
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h8a85ede8;
    ram_cell[       1] = 32'h0;  // 32'hf200f95a;
    ram_cell[       2] = 32'h0;  // 32'h12dab255;
    ram_cell[       3] = 32'h0;  // 32'h542c1f99;
    ram_cell[       4] = 32'h0;  // 32'h24295418;
    ram_cell[       5] = 32'h0;  // 32'h8a0fe7e1;
    ram_cell[       6] = 32'h0;  // 32'hb25e761f;
    ram_cell[       7] = 32'h0;  // 32'hc4d006b4;
    ram_cell[       8] = 32'h0;  // 32'hc1ac13f3;
    ram_cell[       9] = 32'h0;  // 32'h1c618983;
    ram_cell[      10] = 32'h0;  // 32'h9d9e6820;
    ram_cell[      11] = 32'h0;  // 32'h4a7ba8a7;
    ram_cell[      12] = 32'h0;  // 32'h1afbbef1;
    ram_cell[      13] = 32'h0;  // 32'hafd03693;
    ram_cell[      14] = 32'h0;  // 32'h54b1b1bf;
    ram_cell[      15] = 32'h0;  // 32'hb8f4f677;
    ram_cell[      16] = 32'h0;  // 32'h92244e96;
    ram_cell[      17] = 32'h0;  // 32'h396ff671;
    ram_cell[      18] = 32'h0;  // 32'h747a8701;
    ram_cell[      19] = 32'h0;  // 32'hdbab9185;
    ram_cell[      20] = 32'h0;  // 32'h0e4c2306;
    ram_cell[      21] = 32'h0;  // 32'h1c79a259;
    ram_cell[      22] = 32'h0;  // 32'h56c0d1bb;
    ram_cell[      23] = 32'h0;  // 32'ha2853f15;
    ram_cell[      24] = 32'h0;  // 32'h7eda1bb2;
    ram_cell[      25] = 32'h0;  // 32'h47c7616f;
    ram_cell[      26] = 32'h0;  // 32'h8f363449;
    ram_cell[      27] = 32'h0;  // 32'hec2c1852;
    ram_cell[      28] = 32'h0;  // 32'h93d8cf0a;
    ram_cell[      29] = 32'h0;  // 32'h3f7b2df8;
    ram_cell[      30] = 32'h0;  // 32'h1a29d631;
    ram_cell[      31] = 32'h0;  // 32'hea333a90;
    ram_cell[      32] = 32'h0;  // 32'h1f4b8381;
    ram_cell[      33] = 32'h0;  // 32'hd15336cb;
    ram_cell[      34] = 32'h0;  // 32'he02f5180;
    ram_cell[      35] = 32'h0;  // 32'h66acdc8e;
    ram_cell[      36] = 32'h0;  // 32'h1b151614;
    ram_cell[      37] = 32'h0;  // 32'h522c3f9e;
    ram_cell[      38] = 32'h0;  // 32'h8364aab2;
    ram_cell[      39] = 32'h0;  // 32'h3d3b3a27;
    ram_cell[      40] = 32'h0;  // 32'h6d74153f;
    ram_cell[      41] = 32'h0;  // 32'hffe9e025;
    ram_cell[      42] = 32'h0;  // 32'h58d9dbe7;
    ram_cell[      43] = 32'h0;  // 32'h5c80fd59;
    ram_cell[      44] = 32'h0;  // 32'h95226fcb;
    ram_cell[      45] = 32'h0;  // 32'h15943f27;
    ram_cell[      46] = 32'h0;  // 32'h15ecb088;
    ram_cell[      47] = 32'h0;  // 32'hdd0f5116;
    ram_cell[      48] = 32'h0;  // 32'hdc2ed641;
    ram_cell[      49] = 32'h0;  // 32'hb1c68984;
    ram_cell[      50] = 32'h0;  // 32'ha7c126a3;
    ram_cell[      51] = 32'h0;  // 32'h7ecd2f4d;
    ram_cell[      52] = 32'h0;  // 32'h600d2509;
    ram_cell[      53] = 32'h0;  // 32'h1acf7843;
    ram_cell[      54] = 32'h0;  // 32'hf42914da;
    ram_cell[      55] = 32'h0;  // 32'he2ea1d14;
    ram_cell[      56] = 32'h0;  // 32'h75989e8c;
    ram_cell[      57] = 32'h0;  // 32'h8ded9b8a;
    ram_cell[      58] = 32'h0;  // 32'hde45ed70;
    ram_cell[      59] = 32'h0;  // 32'h24ef749e;
    ram_cell[      60] = 32'h0;  // 32'h5fc7f1c3;
    ram_cell[      61] = 32'h0;  // 32'h5c5b1818;
    ram_cell[      62] = 32'h0;  // 32'h50c59809;
    ram_cell[      63] = 32'h0;  // 32'h1f79a586;
    ram_cell[      64] = 32'h0;  // 32'h470eb597;
    ram_cell[      65] = 32'h0;  // 32'ha83de3c9;
    ram_cell[      66] = 32'h0;  // 32'h3f09e736;
    ram_cell[      67] = 32'h0;  // 32'hf6887216;
    ram_cell[      68] = 32'h0;  // 32'h9fceb777;
    ram_cell[      69] = 32'h0;  // 32'h78f1cfc3;
    ram_cell[      70] = 32'h0;  // 32'hdf4dd1d2;
    ram_cell[      71] = 32'h0;  // 32'hb497b362;
    ram_cell[      72] = 32'h0;  // 32'h48d00d9e;
    ram_cell[      73] = 32'h0;  // 32'h137efae6;
    ram_cell[      74] = 32'h0;  // 32'h21c6768d;
    ram_cell[      75] = 32'h0;  // 32'hc09490c0;
    ram_cell[      76] = 32'h0;  // 32'h2e79af96;
    ram_cell[      77] = 32'h0;  // 32'hfb28f4fc;
    ram_cell[      78] = 32'h0;  // 32'h6b1b1266;
    ram_cell[      79] = 32'h0;  // 32'h939ed4dc;
    ram_cell[      80] = 32'h0;  // 32'h2ecefc95;
    ram_cell[      81] = 32'h0;  // 32'h19b5f32f;
    ram_cell[      82] = 32'h0;  // 32'h0fd129fb;
    ram_cell[      83] = 32'h0;  // 32'h855bcf2d;
    ram_cell[      84] = 32'h0;  // 32'h63911ca7;
    ram_cell[      85] = 32'h0;  // 32'hbeba2402;
    ram_cell[      86] = 32'h0;  // 32'hdb4efe4a;
    ram_cell[      87] = 32'h0;  // 32'h8d8efa0e;
    ram_cell[      88] = 32'h0;  // 32'h6faf9d0a;
    ram_cell[      89] = 32'h0;  // 32'h1d7e8482;
    ram_cell[      90] = 32'h0;  // 32'he717498b;
    ram_cell[      91] = 32'h0;  // 32'hf4f96f9b;
    ram_cell[      92] = 32'h0;  // 32'h216adb99;
    ram_cell[      93] = 32'h0;  // 32'h676af661;
    ram_cell[      94] = 32'h0;  // 32'he89e1cde;
    ram_cell[      95] = 32'h0;  // 32'h0aa987ee;
    ram_cell[      96] = 32'h0;  // 32'h0093e782;
    ram_cell[      97] = 32'h0;  // 32'he178087b;
    ram_cell[      98] = 32'h0;  // 32'hc8af43d7;
    ram_cell[      99] = 32'h0;  // 32'h4b5b01ff;
    ram_cell[     100] = 32'h0;  // 32'haf4eb1ce;
    ram_cell[     101] = 32'h0;  // 32'h5ea87b20;
    ram_cell[     102] = 32'h0;  // 32'hc8771020;
    ram_cell[     103] = 32'h0;  // 32'hb3901dfe;
    ram_cell[     104] = 32'h0;  // 32'h96e31f03;
    ram_cell[     105] = 32'h0;  // 32'he4be7eed;
    ram_cell[     106] = 32'h0;  // 32'h9261c09f;
    ram_cell[     107] = 32'h0;  // 32'hef7d562a;
    ram_cell[     108] = 32'h0;  // 32'he2d20a46;
    ram_cell[     109] = 32'h0;  // 32'h69ff9f44;
    ram_cell[     110] = 32'h0;  // 32'h13df006e;
    ram_cell[     111] = 32'h0;  // 32'h4c3f2f42;
    ram_cell[     112] = 32'h0;  // 32'hef7d1fa6;
    ram_cell[     113] = 32'h0;  // 32'hbde9738f;
    ram_cell[     114] = 32'h0;  // 32'h2aad3511;
    ram_cell[     115] = 32'h0;  // 32'h2ae3a94f;
    ram_cell[     116] = 32'h0;  // 32'h12b83ae2;
    ram_cell[     117] = 32'h0;  // 32'h6dd2d770;
    ram_cell[     118] = 32'h0;  // 32'h6aab5c1a;
    ram_cell[     119] = 32'h0;  // 32'h7a65e39d;
    ram_cell[     120] = 32'h0;  // 32'h1f342ef0;
    ram_cell[     121] = 32'h0;  // 32'h57f15797;
    ram_cell[     122] = 32'h0;  // 32'h4022c75c;
    ram_cell[     123] = 32'h0;  // 32'h1e42402c;
    ram_cell[     124] = 32'h0;  // 32'h796a8686;
    ram_cell[     125] = 32'h0;  // 32'h782ff8e3;
    ram_cell[     126] = 32'h0;  // 32'h8be2c8fe;
    ram_cell[     127] = 32'h0;  // 32'h66debddc;
    ram_cell[     128] = 32'h0;  // 32'h0a5ec98b;
    ram_cell[     129] = 32'h0;  // 32'h46dcc4fe;
    ram_cell[     130] = 32'h0;  // 32'h12976ee7;
    ram_cell[     131] = 32'h0;  // 32'hbbf10508;
    ram_cell[     132] = 32'h0;  // 32'h19e8aab3;
    ram_cell[     133] = 32'h0;  // 32'ha6cdd9c2;
    ram_cell[     134] = 32'h0;  // 32'h5be67093;
    ram_cell[     135] = 32'h0;  // 32'h6086c608;
    ram_cell[     136] = 32'h0;  // 32'h54d36bea;
    ram_cell[     137] = 32'h0;  // 32'h002ccf17;
    ram_cell[     138] = 32'h0;  // 32'hd8225e70;
    ram_cell[     139] = 32'h0;  // 32'h95dd6e50;
    ram_cell[     140] = 32'h0;  // 32'h97a99cd8;
    ram_cell[     141] = 32'h0;  // 32'ha8c8ea9d;
    ram_cell[     142] = 32'h0;  // 32'h65b37b2e;
    ram_cell[     143] = 32'h0;  // 32'hcbbade66;
    ram_cell[     144] = 32'h0;  // 32'h50e1464f;
    ram_cell[     145] = 32'h0;  // 32'hef646b15;
    ram_cell[     146] = 32'h0;  // 32'h8e864aaa;
    ram_cell[     147] = 32'h0;  // 32'hdec9f647;
    ram_cell[     148] = 32'h0;  // 32'hd05ddff6;
    ram_cell[     149] = 32'h0;  // 32'h13ec0db3;
    ram_cell[     150] = 32'h0;  // 32'he6c48bbb;
    ram_cell[     151] = 32'h0;  // 32'ha094490f;
    ram_cell[     152] = 32'h0;  // 32'hcae5fcf8;
    ram_cell[     153] = 32'h0;  // 32'hed277ac4;
    ram_cell[     154] = 32'h0;  // 32'h0743565b;
    ram_cell[     155] = 32'h0;  // 32'hf2affadd;
    ram_cell[     156] = 32'h0;  // 32'h82579232;
    ram_cell[     157] = 32'h0;  // 32'h8888e313;
    ram_cell[     158] = 32'h0;  // 32'h824f5ea3;
    ram_cell[     159] = 32'h0;  // 32'h385ac394;
    ram_cell[     160] = 32'h0;  // 32'h4f7872c9;
    ram_cell[     161] = 32'h0;  // 32'hf0fd328c;
    ram_cell[     162] = 32'h0;  // 32'hc99df053;
    ram_cell[     163] = 32'h0;  // 32'he71891e2;
    ram_cell[     164] = 32'h0;  // 32'h233cf720;
    ram_cell[     165] = 32'h0;  // 32'h01768643;
    ram_cell[     166] = 32'h0;  // 32'hef57e30b;
    ram_cell[     167] = 32'h0;  // 32'h0144f8d9;
    ram_cell[     168] = 32'h0;  // 32'h63f9b2c7;
    ram_cell[     169] = 32'h0;  // 32'h98c7b8ae;
    ram_cell[     170] = 32'h0;  // 32'h9cabeef7;
    ram_cell[     171] = 32'h0;  // 32'h18b64631;
    ram_cell[     172] = 32'h0;  // 32'h920dad7c;
    ram_cell[     173] = 32'h0;  // 32'hebabf3b0;
    ram_cell[     174] = 32'h0;  // 32'hc18137fb;
    ram_cell[     175] = 32'h0;  // 32'h4c1f6c04;
    ram_cell[     176] = 32'h0;  // 32'hbb981270;
    ram_cell[     177] = 32'h0;  // 32'he47647a7;
    ram_cell[     178] = 32'h0;  // 32'hd5865d2e;
    ram_cell[     179] = 32'h0;  // 32'h30863016;
    ram_cell[     180] = 32'h0;  // 32'h173da52a;
    ram_cell[     181] = 32'h0;  // 32'h507b5e28;
    ram_cell[     182] = 32'h0;  // 32'h483b199a;
    ram_cell[     183] = 32'h0;  // 32'h46f72a34;
    ram_cell[     184] = 32'h0;  // 32'h84b9775c;
    ram_cell[     185] = 32'h0;  // 32'h4c1a23ab;
    ram_cell[     186] = 32'h0;  // 32'h0b4780bb;
    ram_cell[     187] = 32'h0;  // 32'hd1be9ebe;
    ram_cell[     188] = 32'h0;  // 32'hfc3f79eb;
    ram_cell[     189] = 32'h0;  // 32'h1b4cf376;
    ram_cell[     190] = 32'h0;  // 32'h2dbc7c04;
    ram_cell[     191] = 32'h0;  // 32'h5bad8e49;
    ram_cell[     192] = 32'h0;  // 32'h1dbb1038;
    ram_cell[     193] = 32'h0;  // 32'had0e1e34;
    ram_cell[     194] = 32'h0;  // 32'h825265e5;
    ram_cell[     195] = 32'h0;  // 32'hcebb3638;
    ram_cell[     196] = 32'h0;  // 32'ha4a64f99;
    ram_cell[     197] = 32'h0;  // 32'h6158b03e;
    ram_cell[     198] = 32'h0;  // 32'hc81dc1e2;
    ram_cell[     199] = 32'h0;  // 32'hcb13a146;
    ram_cell[     200] = 32'h0;  // 32'h87c05257;
    ram_cell[     201] = 32'h0;  // 32'h4839d680;
    ram_cell[     202] = 32'h0;  // 32'h3e2f39da;
    ram_cell[     203] = 32'h0;  // 32'h6446260a;
    ram_cell[     204] = 32'h0;  // 32'h174a1864;
    ram_cell[     205] = 32'h0;  // 32'h256aa009;
    ram_cell[     206] = 32'h0;  // 32'h7df06d3b;
    ram_cell[     207] = 32'h0;  // 32'hfe7804a4;
    ram_cell[     208] = 32'h0;  // 32'he779536e;
    ram_cell[     209] = 32'h0;  // 32'hd80ae6a6;
    ram_cell[     210] = 32'h0;  // 32'h5f755ed5;
    ram_cell[     211] = 32'h0;  // 32'h5ece0711;
    ram_cell[     212] = 32'h0;  // 32'h3b22e052;
    ram_cell[     213] = 32'h0;  // 32'haa41d680;
    ram_cell[     214] = 32'h0;  // 32'h7c30d37a;
    ram_cell[     215] = 32'h0;  // 32'h801e80d1;
    ram_cell[     216] = 32'h0;  // 32'h2cf99747;
    ram_cell[     217] = 32'h0;  // 32'he4a86414;
    ram_cell[     218] = 32'h0;  // 32'hba12718a;
    ram_cell[     219] = 32'h0;  // 32'h6a85e929;
    ram_cell[     220] = 32'h0;  // 32'h0f4dca48;
    ram_cell[     221] = 32'h0;  // 32'h1ee766a6;
    ram_cell[     222] = 32'h0;  // 32'h694c2e2e;
    ram_cell[     223] = 32'h0;  // 32'h8a948e44;
    ram_cell[     224] = 32'h0;  // 32'h0bc835a8;
    ram_cell[     225] = 32'h0;  // 32'h63ee42ea;
    ram_cell[     226] = 32'h0;  // 32'h500877dd;
    ram_cell[     227] = 32'h0;  // 32'h9279875f;
    ram_cell[     228] = 32'h0;  // 32'ha00279cb;
    ram_cell[     229] = 32'h0;  // 32'h5ecaf13b;
    ram_cell[     230] = 32'h0;  // 32'hcd1a04c3;
    ram_cell[     231] = 32'h0;  // 32'haeaed285;
    ram_cell[     232] = 32'h0;  // 32'h88d595af;
    ram_cell[     233] = 32'h0;  // 32'h0973f418;
    ram_cell[     234] = 32'h0;  // 32'h036b2141;
    ram_cell[     235] = 32'h0;  // 32'h37fb3f13;
    ram_cell[     236] = 32'h0;  // 32'hff3dd08d;
    ram_cell[     237] = 32'h0;  // 32'h0b37dda2;
    ram_cell[     238] = 32'h0;  // 32'h04549d61;
    ram_cell[     239] = 32'h0;  // 32'h173ce662;
    ram_cell[     240] = 32'h0;  // 32'h2c4c9cba;
    ram_cell[     241] = 32'h0;  // 32'he70aa5f5;
    ram_cell[     242] = 32'h0;  // 32'h2e98fcca;
    ram_cell[     243] = 32'h0;  // 32'hf4d14598;
    ram_cell[     244] = 32'h0;  // 32'h4ee148ae;
    ram_cell[     245] = 32'h0;  // 32'h0abae3ed;
    ram_cell[     246] = 32'h0;  // 32'h298375c3;
    ram_cell[     247] = 32'h0;  // 32'h357bea94;
    ram_cell[     248] = 32'h0;  // 32'haaff261f;
    ram_cell[     249] = 32'h0;  // 32'ha2feab78;
    ram_cell[     250] = 32'h0;  // 32'h4edc0d3a;
    ram_cell[     251] = 32'h0;  // 32'h863fa88d;
    ram_cell[     252] = 32'h0;  // 32'h99c1a071;
    ram_cell[     253] = 32'h0;  // 32'h0fa386ab;
    ram_cell[     254] = 32'h0;  // 32'h480c9db0;
    ram_cell[     255] = 32'h0;  // 32'h8b0040ce;
    ram_cell[     256] = 32'h0;  // 32'h71ffabcc;
    ram_cell[     257] = 32'h0;  // 32'hb5825a5a;
    ram_cell[     258] = 32'h0;  // 32'h223b8b03;
    ram_cell[     259] = 32'h0;  // 32'h077936dd;
    ram_cell[     260] = 32'h0;  // 32'h2631ebfa;
    ram_cell[     261] = 32'h0;  // 32'h37da03a5;
    ram_cell[     262] = 32'h0;  // 32'h351ce60c;
    ram_cell[     263] = 32'h0;  // 32'h555656dc;
    ram_cell[     264] = 32'h0;  // 32'h6c7b8f5c;
    ram_cell[     265] = 32'h0;  // 32'h70ba632a;
    ram_cell[     266] = 32'h0;  // 32'h47360d84;
    ram_cell[     267] = 32'h0;  // 32'hab515be1;
    ram_cell[     268] = 32'h0;  // 32'h6277af10;
    ram_cell[     269] = 32'h0;  // 32'h25a6a6cb;
    ram_cell[     270] = 32'h0;  // 32'h2a4e1071;
    ram_cell[     271] = 32'h0;  // 32'h4a8f191d;
    ram_cell[     272] = 32'h0;  // 32'h40cef21e;
    ram_cell[     273] = 32'h0;  // 32'h2e97407c;
    ram_cell[     274] = 32'h0;  // 32'h4dd16204;
    ram_cell[     275] = 32'h0;  // 32'h8e8e0411;
    ram_cell[     276] = 32'h0;  // 32'h3a17c3cc;
    ram_cell[     277] = 32'h0;  // 32'h168b092c;
    ram_cell[     278] = 32'h0;  // 32'h7b4fc6e2;
    ram_cell[     279] = 32'h0;  // 32'h4a49eb8d;
    ram_cell[     280] = 32'h0;  // 32'hcce9a047;
    ram_cell[     281] = 32'h0;  // 32'h284b0660;
    ram_cell[     282] = 32'h0;  // 32'hfb64dba9;
    ram_cell[     283] = 32'h0;  // 32'hda78414d;
    ram_cell[     284] = 32'h0;  // 32'h9648d115;
    ram_cell[     285] = 32'h0;  // 32'h2d51dddc;
    ram_cell[     286] = 32'h0;  // 32'hec89ba0d;
    ram_cell[     287] = 32'h0;  // 32'h7cc5e489;
    ram_cell[     288] = 32'h0;  // 32'h58de36d4;
    ram_cell[     289] = 32'h0;  // 32'he2db61e5;
    ram_cell[     290] = 32'h0;  // 32'hcf69c611;
    ram_cell[     291] = 32'h0;  // 32'hf7fd0512;
    ram_cell[     292] = 32'h0;  // 32'h2f1ed2bf;
    ram_cell[     293] = 32'h0;  // 32'h2c109663;
    ram_cell[     294] = 32'h0;  // 32'heb2d3316;
    ram_cell[     295] = 32'h0;  // 32'h5f0bd83f;
    ram_cell[     296] = 32'h0;  // 32'hf5e398fd;
    ram_cell[     297] = 32'h0;  // 32'h4f4cb4ab;
    ram_cell[     298] = 32'h0;  // 32'h1ae24208;
    ram_cell[     299] = 32'h0;  // 32'h26fb58b0;
    ram_cell[     300] = 32'h0;  // 32'h6b3aeb4f;
    ram_cell[     301] = 32'h0;  // 32'hc7835e15;
    ram_cell[     302] = 32'h0;  // 32'hd6df5545;
    ram_cell[     303] = 32'h0;  // 32'h1227b2eb;
    ram_cell[     304] = 32'h0;  // 32'hf02a020d;
    ram_cell[     305] = 32'h0;  // 32'hf5f01577;
    ram_cell[     306] = 32'h0;  // 32'h52c18f7c;
    ram_cell[     307] = 32'h0;  // 32'hac96d69b;
    ram_cell[     308] = 32'h0;  // 32'ha1300004;
    ram_cell[     309] = 32'h0;  // 32'h74c4c0f1;
    ram_cell[     310] = 32'h0;  // 32'h126697c2;
    ram_cell[     311] = 32'h0;  // 32'h5a074efe;
    ram_cell[     312] = 32'h0;  // 32'hcc14a0db;
    ram_cell[     313] = 32'h0;  // 32'h3d1e9197;
    ram_cell[     314] = 32'h0;  // 32'h79b7becc;
    ram_cell[     315] = 32'h0;  // 32'hdaf58fdd;
    ram_cell[     316] = 32'h0;  // 32'h7a0c7b48;
    ram_cell[     317] = 32'h0;  // 32'h6c2501c0;
    ram_cell[     318] = 32'h0;  // 32'h08d587ed;
    ram_cell[     319] = 32'h0;  // 32'h84686e6f;
    ram_cell[     320] = 32'h0;  // 32'h4ffdebee;
    ram_cell[     321] = 32'h0;  // 32'ha417e0b5;
    ram_cell[     322] = 32'h0;  // 32'h29516d73;
    ram_cell[     323] = 32'h0;  // 32'h93a0d31e;
    ram_cell[     324] = 32'h0;  // 32'hd36a6fcf;
    ram_cell[     325] = 32'h0;  // 32'h5b9ca3be;
    ram_cell[     326] = 32'h0;  // 32'he22d40d7;
    ram_cell[     327] = 32'h0;  // 32'h4eddedd8;
    ram_cell[     328] = 32'h0;  // 32'h6a9bc3d7;
    ram_cell[     329] = 32'h0;  // 32'hb0165d47;
    ram_cell[     330] = 32'h0;  // 32'ha636b09a;
    ram_cell[     331] = 32'h0;  // 32'hb0dcdb53;
    ram_cell[     332] = 32'h0;  // 32'hb548ec4c;
    ram_cell[     333] = 32'h0;  // 32'h266422f4;
    ram_cell[     334] = 32'h0;  // 32'hbb3d34bf;
    ram_cell[     335] = 32'h0;  // 32'h5c9ffb7f;
    ram_cell[     336] = 32'h0;  // 32'h77f861c0;
    ram_cell[     337] = 32'h0;  // 32'hf20a5129;
    ram_cell[     338] = 32'h0;  // 32'h3f860aec;
    ram_cell[     339] = 32'h0;  // 32'h719e5be0;
    ram_cell[     340] = 32'h0;  // 32'h6189b47b;
    ram_cell[     341] = 32'h0;  // 32'ha24215da;
    ram_cell[     342] = 32'h0;  // 32'h4c6a83fa;
    ram_cell[     343] = 32'h0;  // 32'hae0a73f4;
    ram_cell[     344] = 32'h0;  // 32'h324079ae;
    ram_cell[     345] = 32'h0;  // 32'h35314fad;
    ram_cell[     346] = 32'h0;  // 32'hf9425acd;
    ram_cell[     347] = 32'h0;  // 32'h4aa8f513;
    ram_cell[     348] = 32'h0;  // 32'h4c03dc1a;
    ram_cell[     349] = 32'h0;  // 32'h7f5debb3;
    ram_cell[     350] = 32'h0;  // 32'h636983a8;
    ram_cell[     351] = 32'h0;  // 32'h1a0142d6;
    ram_cell[     352] = 32'h0;  // 32'hd6a43d80;
    ram_cell[     353] = 32'h0;  // 32'h9cc8747e;
    ram_cell[     354] = 32'h0;  // 32'h4e6cc9d5;
    ram_cell[     355] = 32'h0;  // 32'ha890c308;
    ram_cell[     356] = 32'h0;  // 32'he7c6dab5;
    ram_cell[     357] = 32'h0;  // 32'hed1dc55a;
    ram_cell[     358] = 32'h0;  // 32'h8621923f;
    ram_cell[     359] = 32'h0;  // 32'hfb1c57ca;
    ram_cell[     360] = 32'h0;  // 32'h4a61ab14;
    ram_cell[     361] = 32'h0;  // 32'ha99fc6f7;
    ram_cell[     362] = 32'h0;  // 32'h32593047;
    ram_cell[     363] = 32'h0;  // 32'h2e40f806;
    ram_cell[     364] = 32'h0;  // 32'h6a1dec2e;
    ram_cell[     365] = 32'h0;  // 32'hd2830b21;
    ram_cell[     366] = 32'h0;  // 32'hbe45ec91;
    ram_cell[     367] = 32'h0;  // 32'h5b402bac;
    ram_cell[     368] = 32'h0;  // 32'h77fd68a0;
    ram_cell[     369] = 32'h0;  // 32'h9d878f0b;
    ram_cell[     370] = 32'h0;  // 32'hef340082;
    ram_cell[     371] = 32'h0;  // 32'hc977cf7e;
    ram_cell[     372] = 32'h0;  // 32'hd408260b;
    ram_cell[     373] = 32'h0;  // 32'h9c1b7356;
    ram_cell[     374] = 32'h0;  // 32'h20d98d40;
    ram_cell[     375] = 32'h0;  // 32'hb35a08a8;
    ram_cell[     376] = 32'h0;  // 32'hc8bec348;
    ram_cell[     377] = 32'h0;  // 32'h854920f2;
    ram_cell[     378] = 32'h0;  // 32'h23799f72;
    ram_cell[     379] = 32'h0;  // 32'hbea463cd;
    ram_cell[     380] = 32'h0;  // 32'h451cc24a;
    ram_cell[     381] = 32'h0;  // 32'h44d7df74;
    ram_cell[     382] = 32'h0;  // 32'ha8f02768;
    ram_cell[     383] = 32'h0;  // 32'hd36ac33e;
    ram_cell[     384] = 32'h0;  // 32'ha8e87948;
    ram_cell[     385] = 32'h0;  // 32'h383f7c39;
    ram_cell[     386] = 32'h0;  // 32'h6c56a44a;
    ram_cell[     387] = 32'h0;  // 32'h425647bc;
    ram_cell[     388] = 32'h0;  // 32'he9351036;
    ram_cell[     389] = 32'h0;  // 32'hbaa57b3d;
    ram_cell[     390] = 32'h0;  // 32'h502db97b;
    ram_cell[     391] = 32'h0;  // 32'hd10382b1;
    ram_cell[     392] = 32'h0;  // 32'h3a907481;
    ram_cell[     393] = 32'h0;  // 32'h876784f6;
    ram_cell[     394] = 32'h0;  // 32'h2602d29d;
    ram_cell[     395] = 32'h0;  // 32'h4d3a2743;
    ram_cell[     396] = 32'h0;  // 32'h3afd6174;
    ram_cell[     397] = 32'h0;  // 32'h237e7edb;
    ram_cell[     398] = 32'h0;  // 32'h02f57d64;
    ram_cell[     399] = 32'h0;  // 32'h11c30764;
    ram_cell[     400] = 32'h0;  // 32'h30b10a42;
    ram_cell[     401] = 32'h0;  // 32'h4b142dab;
    ram_cell[     402] = 32'h0;  // 32'hebabdd43;
    ram_cell[     403] = 32'h0;  // 32'h591905af;
    ram_cell[     404] = 32'h0;  // 32'h2850c3fe;
    ram_cell[     405] = 32'h0;  // 32'h0f9d72dd;
    ram_cell[     406] = 32'h0;  // 32'hfcbbc781;
    ram_cell[     407] = 32'h0;  // 32'h00d23f97;
    ram_cell[     408] = 32'h0;  // 32'h4a1c6be6;
    ram_cell[     409] = 32'h0;  // 32'h7fbe7743;
    ram_cell[     410] = 32'h0;  // 32'h5572a301;
    ram_cell[     411] = 32'h0;  // 32'h66a321be;
    ram_cell[     412] = 32'h0;  // 32'h4dc957cc;
    ram_cell[     413] = 32'h0;  // 32'h46ae78c5;
    ram_cell[     414] = 32'h0;  // 32'h9ff19a3c;
    ram_cell[     415] = 32'h0;  // 32'h729995de;
    ram_cell[     416] = 32'h0;  // 32'hd5090b7f;
    ram_cell[     417] = 32'h0;  // 32'h61da6b12;
    ram_cell[     418] = 32'h0;  // 32'hdfd5b54e;
    ram_cell[     419] = 32'h0;  // 32'h00cb75bf;
    ram_cell[     420] = 32'h0;  // 32'h2aa8d5d6;
    ram_cell[     421] = 32'h0;  // 32'h889088a3;
    ram_cell[     422] = 32'h0;  // 32'h312650a8;
    ram_cell[     423] = 32'h0;  // 32'hacbc7a9c;
    ram_cell[     424] = 32'h0;  // 32'h3b89988d;
    ram_cell[     425] = 32'h0;  // 32'h722a39bb;
    ram_cell[     426] = 32'h0;  // 32'h9cc2c83c;
    ram_cell[     427] = 32'h0;  // 32'h07efa0c0;
    ram_cell[     428] = 32'h0;  // 32'h4c380b7f;
    ram_cell[     429] = 32'h0;  // 32'h0e75bdb0;
    ram_cell[     430] = 32'h0;  // 32'h5d9d35bd;
    ram_cell[     431] = 32'h0;  // 32'h7d3461de;
    ram_cell[     432] = 32'h0;  // 32'h29f84010;
    ram_cell[     433] = 32'h0;  // 32'h58c2f61c;
    ram_cell[     434] = 32'h0;  // 32'h1e837075;
    ram_cell[     435] = 32'h0;  // 32'hbc2449fd;
    ram_cell[     436] = 32'h0;  // 32'h2aec7cde;
    ram_cell[     437] = 32'h0;  // 32'ha395b02b;
    ram_cell[     438] = 32'h0;  // 32'h5221a9b5;
    ram_cell[     439] = 32'h0;  // 32'h3982aa6c;
    ram_cell[     440] = 32'h0;  // 32'hc95ba4c8;
    ram_cell[     441] = 32'h0;  // 32'h792231e3;
    ram_cell[     442] = 32'h0;  // 32'h7aad02ad;
    ram_cell[     443] = 32'h0;  // 32'hd57b1295;
    ram_cell[     444] = 32'h0;  // 32'h6d515e3d;
    ram_cell[     445] = 32'h0;  // 32'h26d09868;
    ram_cell[     446] = 32'h0;  // 32'he64cec81;
    ram_cell[     447] = 32'h0;  // 32'h63b02bf9;
    ram_cell[     448] = 32'h0;  // 32'h1ee932d8;
    ram_cell[     449] = 32'h0;  // 32'h3e428f29;
    ram_cell[     450] = 32'h0;  // 32'hc6b63697;
    ram_cell[     451] = 32'h0;  // 32'hda2795e4;
    ram_cell[     452] = 32'h0;  // 32'h3d1ae58c;
    ram_cell[     453] = 32'h0;  // 32'hd2bc2839;
    ram_cell[     454] = 32'h0;  // 32'h8e98333b;
    ram_cell[     455] = 32'h0;  // 32'h61c13e58;
    ram_cell[     456] = 32'h0;  // 32'h7061ad1a;
    ram_cell[     457] = 32'h0;  // 32'h246ef588;
    ram_cell[     458] = 32'h0;  // 32'h32e74e25;
    ram_cell[     459] = 32'h0;  // 32'h5593f508;
    ram_cell[     460] = 32'h0;  // 32'h7ab7e0f9;
    ram_cell[     461] = 32'h0;  // 32'hf7bf1f9e;
    ram_cell[     462] = 32'h0;  // 32'h2dbedd5b;
    ram_cell[     463] = 32'h0;  // 32'hdf5fed45;
    ram_cell[     464] = 32'h0;  // 32'hd3e9f879;
    ram_cell[     465] = 32'h0;  // 32'he9aedd21;
    ram_cell[     466] = 32'h0;  // 32'h0289c1d1;
    ram_cell[     467] = 32'h0;  // 32'h3c91e86c;
    ram_cell[     468] = 32'h0;  // 32'h2798ddad;
    ram_cell[     469] = 32'h0;  // 32'hc4836875;
    ram_cell[     470] = 32'h0;  // 32'h6762218d;
    ram_cell[     471] = 32'h0;  // 32'h04723a2f;
    ram_cell[     472] = 32'h0;  // 32'h16d71b4b;
    ram_cell[     473] = 32'h0;  // 32'haa06486f;
    ram_cell[     474] = 32'h0;  // 32'h58daf1b1;
    ram_cell[     475] = 32'h0;  // 32'hd106d65d;
    ram_cell[     476] = 32'h0;  // 32'hbf12bfe7;
    ram_cell[     477] = 32'h0;  // 32'hb0b82b26;
    ram_cell[     478] = 32'h0;  // 32'hbf960efb;
    ram_cell[     479] = 32'h0;  // 32'hb3986003;
    ram_cell[     480] = 32'h0;  // 32'h67bd49b2;
    ram_cell[     481] = 32'h0;  // 32'h6e150284;
    ram_cell[     482] = 32'h0;  // 32'h4b71c5b6;
    ram_cell[     483] = 32'h0;  // 32'h5341c42d;
    ram_cell[     484] = 32'h0;  // 32'hd771e766;
    ram_cell[     485] = 32'h0;  // 32'h5442d5e4;
    ram_cell[     486] = 32'h0;  // 32'h178ffc9d;
    ram_cell[     487] = 32'h0;  // 32'hef5a7a63;
    ram_cell[     488] = 32'h0;  // 32'h68ff78eb;
    ram_cell[     489] = 32'h0;  // 32'hf2ca7453;
    ram_cell[     490] = 32'h0;  // 32'hf120ab20;
    ram_cell[     491] = 32'h0;  // 32'hf3652d84;
    ram_cell[     492] = 32'h0;  // 32'h1c66b2ff;
    ram_cell[     493] = 32'h0;  // 32'h08b74b1c;
    ram_cell[     494] = 32'h0;  // 32'h8ab55933;
    ram_cell[     495] = 32'h0;  // 32'h1ee44b18;
    ram_cell[     496] = 32'h0;  // 32'hb75c0b03;
    ram_cell[     497] = 32'h0;  // 32'h5e4cadf6;
    ram_cell[     498] = 32'h0;  // 32'h71132c00;
    ram_cell[     499] = 32'h0;  // 32'hc754e7af;
    ram_cell[     500] = 32'h0;  // 32'hc48bd5e9;
    ram_cell[     501] = 32'h0;  // 32'h6c4b29c6;
    ram_cell[     502] = 32'h0;  // 32'h823fe642;
    ram_cell[     503] = 32'h0;  // 32'ha20cab6a;
    ram_cell[     504] = 32'h0;  // 32'hfbca592d;
    ram_cell[     505] = 32'h0;  // 32'h81730b32;
    ram_cell[     506] = 32'h0;  // 32'h532ce39f;
    ram_cell[     507] = 32'h0;  // 32'h9d44b012;
    ram_cell[     508] = 32'h0;  // 32'hc0743b1f;
    ram_cell[     509] = 32'h0;  // 32'h554ce126;
    ram_cell[     510] = 32'h0;  // 32'hc97d1788;
    ram_cell[     511] = 32'h0;  // 32'h39359609;
    ram_cell[     512] = 32'h0;  // 32'hb4bdfc3a;
    ram_cell[     513] = 32'h0;  // 32'h3d3d3d82;
    ram_cell[     514] = 32'h0;  // 32'h245e1d0b;
    ram_cell[     515] = 32'h0;  // 32'h9bdbb859;
    ram_cell[     516] = 32'h0;  // 32'hbbeeca4c;
    ram_cell[     517] = 32'h0;  // 32'hf97d09be;
    ram_cell[     518] = 32'h0;  // 32'h504e91d0;
    ram_cell[     519] = 32'h0;  // 32'h7ade7471;
    ram_cell[     520] = 32'h0;  // 32'h461cfcd1;
    ram_cell[     521] = 32'h0;  // 32'h125792b9;
    ram_cell[     522] = 32'h0;  // 32'h6d6cea97;
    ram_cell[     523] = 32'h0;  // 32'h589aab3e;
    ram_cell[     524] = 32'h0;  // 32'hdb59f888;
    ram_cell[     525] = 32'h0;  // 32'h2d3f09ca;
    ram_cell[     526] = 32'h0;  // 32'h667353eb;
    ram_cell[     527] = 32'h0;  // 32'hcdc120fe;
    ram_cell[     528] = 32'h0;  // 32'h1093b22e;
    ram_cell[     529] = 32'h0;  // 32'h88ed91f2;
    ram_cell[     530] = 32'h0;  // 32'hdbe67196;
    ram_cell[     531] = 32'h0;  // 32'h85b0de88;
    ram_cell[     532] = 32'h0;  // 32'h1bbaee4a;
    ram_cell[     533] = 32'h0;  // 32'h498c4cab;
    ram_cell[     534] = 32'h0;  // 32'h9afb5d79;
    ram_cell[     535] = 32'h0;  // 32'h36f9ac4a;
    ram_cell[     536] = 32'h0;  // 32'h0028bd36;
    ram_cell[     537] = 32'h0;  // 32'h2743c1e8;
    ram_cell[     538] = 32'h0;  // 32'h4d926ea3;
    ram_cell[     539] = 32'h0;  // 32'hf9ceb0c5;
    ram_cell[     540] = 32'h0;  // 32'hfdde39f3;
    ram_cell[     541] = 32'h0;  // 32'hfbe56c7c;
    ram_cell[     542] = 32'h0;  // 32'h12fc03b4;
    ram_cell[     543] = 32'h0;  // 32'h9ae9a8b7;
    ram_cell[     544] = 32'h0;  // 32'hf40a496c;
    ram_cell[     545] = 32'h0;  // 32'he6bbc9a2;
    ram_cell[     546] = 32'h0;  // 32'h43c93813;
    ram_cell[     547] = 32'h0;  // 32'h8a4879bb;
    ram_cell[     548] = 32'h0;  // 32'h33c2a3fc;
    ram_cell[     549] = 32'h0;  // 32'hcd475173;
    ram_cell[     550] = 32'h0;  // 32'hf3609092;
    ram_cell[     551] = 32'h0;  // 32'h2223c1a1;
    ram_cell[     552] = 32'h0;  // 32'h142bc881;
    ram_cell[     553] = 32'h0;  // 32'hdc33622f;
    ram_cell[     554] = 32'h0;  // 32'h209d619c;
    ram_cell[     555] = 32'h0;  // 32'hb4e83b05;
    ram_cell[     556] = 32'h0;  // 32'h53fcb762;
    ram_cell[     557] = 32'h0;  // 32'hb4a8d657;
    ram_cell[     558] = 32'h0;  // 32'ha14561f2;
    ram_cell[     559] = 32'h0;  // 32'h13041897;
    ram_cell[     560] = 32'h0;  // 32'h760de09d;
    ram_cell[     561] = 32'h0;  // 32'h8d7b1f2a;
    ram_cell[     562] = 32'h0;  // 32'h98bb632e;
    ram_cell[     563] = 32'h0;  // 32'h30513a34;
    ram_cell[     564] = 32'h0;  // 32'h09291961;
    ram_cell[     565] = 32'h0;  // 32'hefb42897;
    ram_cell[     566] = 32'h0;  // 32'hd868fe3e;
    ram_cell[     567] = 32'h0;  // 32'h40c8a892;
    ram_cell[     568] = 32'h0;  // 32'h9a4fc9cf;
    ram_cell[     569] = 32'h0;  // 32'h354f926f;
    ram_cell[     570] = 32'h0;  // 32'h9e1ee94e;
    ram_cell[     571] = 32'h0;  // 32'hb3d7ab41;
    ram_cell[     572] = 32'h0;  // 32'hd4ee964f;
    ram_cell[     573] = 32'h0;  // 32'ha17d15be;
    ram_cell[     574] = 32'h0;  // 32'hc9405f0f;
    ram_cell[     575] = 32'h0;  // 32'h5c1e68b5;
    ram_cell[     576] = 32'h0;  // 32'h431b917b;
    ram_cell[     577] = 32'h0;  // 32'heedce5e9;
    ram_cell[     578] = 32'h0;  // 32'h8370b675;
    ram_cell[     579] = 32'h0;  // 32'h5233c6e0;
    ram_cell[     580] = 32'h0;  // 32'heddf6a7c;
    ram_cell[     581] = 32'h0;  // 32'hfbbcfcbd;
    ram_cell[     582] = 32'h0;  // 32'hb4985ed6;
    ram_cell[     583] = 32'h0;  // 32'hdd09139d;
    ram_cell[     584] = 32'h0;  // 32'hffb782c5;
    ram_cell[     585] = 32'h0;  // 32'h41f6d920;
    ram_cell[     586] = 32'h0;  // 32'h8c491f1b;
    ram_cell[     587] = 32'h0;  // 32'h976c8a28;
    ram_cell[     588] = 32'h0;  // 32'h2eb4e44c;
    ram_cell[     589] = 32'h0;  // 32'h1f2bed70;
    ram_cell[     590] = 32'h0;  // 32'hb3f32544;
    ram_cell[     591] = 32'h0;  // 32'h05016346;
    ram_cell[     592] = 32'h0;  // 32'h0b1f33e4;
    ram_cell[     593] = 32'h0;  // 32'h8437f54c;
    ram_cell[     594] = 32'h0;  // 32'h99379a8d;
    ram_cell[     595] = 32'h0;  // 32'h876368c4;
    ram_cell[     596] = 32'h0;  // 32'hd5dce853;
    ram_cell[     597] = 32'h0;  // 32'h13664295;
    ram_cell[     598] = 32'h0;  // 32'he36168be;
    ram_cell[     599] = 32'h0;  // 32'hb236f0c3;
    ram_cell[     600] = 32'h0;  // 32'h44f1573b;
    ram_cell[     601] = 32'h0;  // 32'h7c2faa4f;
    ram_cell[     602] = 32'h0;  // 32'h9aabb8c2;
    ram_cell[     603] = 32'h0;  // 32'h9641ca84;
    ram_cell[     604] = 32'h0;  // 32'h4c0a1b68;
    ram_cell[     605] = 32'h0;  // 32'h4059b97f;
    ram_cell[     606] = 32'h0;  // 32'h1bd6bcab;
    ram_cell[     607] = 32'h0;  // 32'h1fff0e16;
    ram_cell[     608] = 32'h0;  // 32'h12c71c35;
    ram_cell[     609] = 32'h0;  // 32'h63078ae7;
    ram_cell[     610] = 32'h0;  // 32'h655282ad;
    ram_cell[     611] = 32'h0;  // 32'h6206beb8;
    ram_cell[     612] = 32'h0;  // 32'h92b0fee8;
    ram_cell[     613] = 32'h0;  // 32'h656fb397;
    ram_cell[     614] = 32'h0;  // 32'h3ec0c30a;
    ram_cell[     615] = 32'h0;  // 32'h8b927eb7;
    ram_cell[     616] = 32'h0;  // 32'h931258d3;
    ram_cell[     617] = 32'h0;  // 32'h0cd349ad;
    ram_cell[     618] = 32'h0;  // 32'h59201642;
    ram_cell[     619] = 32'h0;  // 32'h54d10e40;
    ram_cell[     620] = 32'h0;  // 32'ha1240ea2;
    ram_cell[     621] = 32'h0;  // 32'hd0bec26e;
    ram_cell[     622] = 32'h0;  // 32'h385a26d2;
    ram_cell[     623] = 32'h0;  // 32'h48e08b0a;
    ram_cell[     624] = 32'h0;  // 32'ha2c55590;
    ram_cell[     625] = 32'h0;  // 32'h72bb68ef;
    ram_cell[     626] = 32'h0;  // 32'he7b7e5e1;
    ram_cell[     627] = 32'h0;  // 32'hbcb83b62;
    ram_cell[     628] = 32'h0;  // 32'h61fc93cb;
    ram_cell[     629] = 32'h0;  // 32'h4856e1cf;
    ram_cell[     630] = 32'h0;  // 32'h9d0da943;
    ram_cell[     631] = 32'h0;  // 32'he241365e;
    ram_cell[     632] = 32'h0;  // 32'h8091ac01;
    ram_cell[     633] = 32'h0;  // 32'ha7ef103a;
    ram_cell[     634] = 32'h0;  // 32'ha8143004;
    ram_cell[     635] = 32'h0;  // 32'h1c226849;
    ram_cell[     636] = 32'h0;  // 32'h31c5a9f2;
    ram_cell[     637] = 32'h0;  // 32'h441d28f8;
    ram_cell[     638] = 32'h0;  // 32'hd69afaad;
    ram_cell[     639] = 32'h0;  // 32'h864dcf7b;
    ram_cell[     640] = 32'h0;  // 32'h440cfea3;
    ram_cell[     641] = 32'h0;  // 32'h76cfdd45;
    ram_cell[     642] = 32'h0;  // 32'h65539144;
    ram_cell[     643] = 32'h0;  // 32'hc7ff59bd;
    ram_cell[     644] = 32'h0;  // 32'h2e15a711;
    ram_cell[     645] = 32'h0;  // 32'h03d89dbb;
    ram_cell[     646] = 32'h0;  // 32'he1165cd2;
    ram_cell[     647] = 32'h0;  // 32'h3c16db1d;
    ram_cell[     648] = 32'h0;  // 32'heb7f5236;
    ram_cell[     649] = 32'h0;  // 32'h15063eda;
    ram_cell[     650] = 32'h0;  // 32'h88589c52;
    ram_cell[     651] = 32'h0;  // 32'hba91b210;
    ram_cell[     652] = 32'h0;  // 32'h201b072c;
    ram_cell[     653] = 32'h0;  // 32'h73946f8c;
    ram_cell[     654] = 32'h0;  // 32'h5b2d5019;
    ram_cell[     655] = 32'h0;  // 32'h48f9b728;
    ram_cell[     656] = 32'h0;  // 32'h2a262c6f;
    ram_cell[     657] = 32'h0;  // 32'he6e79f3d;
    ram_cell[     658] = 32'h0;  // 32'h7c55aecf;
    ram_cell[     659] = 32'h0;  // 32'he483716a;
    ram_cell[     660] = 32'h0;  // 32'h6dac190e;
    ram_cell[     661] = 32'h0;  // 32'hbc5aced4;
    ram_cell[     662] = 32'h0;  // 32'hed8458ef;
    ram_cell[     663] = 32'h0;  // 32'h93b8744f;
    ram_cell[     664] = 32'h0;  // 32'h5652d2a6;
    ram_cell[     665] = 32'h0;  // 32'h4806b21e;
    ram_cell[     666] = 32'h0;  // 32'hc07cd9c9;
    ram_cell[     667] = 32'h0;  // 32'h2cb35577;
    ram_cell[     668] = 32'h0;  // 32'h61538cef;
    ram_cell[     669] = 32'h0;  // 32'h2bdb0759;
    ram_cell[     670] = 32'h0;  // 32'hdf66d4da;
    ram_cell[     671] = 32'h0;  // 32'h65b380fd;
    ram_cell[     672] = 32'h0;  // 32'hcc077687;
    ram_cell[     673] = 32'h0;  // 32'hc6bcd012;
    ram_cell[     674] = 32'h0;  // 32'h0184099d;
    ram_cell[     675] = 32'h0;  // 32'h60158d87;
    ram_cell[     676] = 32'h0;  // 32'hb508b8c7;
    ram_cell[     677] = 32'h0;  // 32'h6781226f;
    ram_cell[     678] = 32'h0;  // 32'h77693abc;
    ram_cell[     679] = 32'h0;  // 32'h4bf78cbc;
    ram_cell[     680] = 32'h0;  // 32'h749eb05d;
    ram_cell[     681] = 32'h0;  // 32'h13df2385;
    ram_cell[     682] = 32'h0;  // 32'h3b754d43;
    ram_cell[     683] = 32'h0;  // 32'h63c2166b;
    ram_cell[     684] = 32'h0;  // 32'hcd9bf788;
    ram_cell[     685] = 32'h0;  // 32'hc0b3bf8c;
    ram_cell[     686] = 32'h0;  // 32'h725a5665;
    ram_cell[     687] = 32'h0;  // 32'h14b62795;
    ram_cell[     688] = 32'h0;  // 32'h04a60877;
    ram_cell[     689] = 32'h0;  // 32'h6b935b94;
    ram_cell[     690] = 32'h0;  // 32'hca03ce85;
    ram_cell[     691] = 32'h0;  // 32'hc4e8859c;
    ram_cell[     692] = 32'h0;  // 32'h28f5acd2;
    ram_cell[     693] = 32'h0;  // 32'h8e7f9cfb;
    ram_cell[     694] = 32'h0;  // 32'h335fad8c;
    ram_cell[     695] = 32'h0;  // 32'hfc3af928;
    ram_cell[     696] = 32'h0;  // 32'h882bb38c;
    ram_cell[     697] = 32'h0;  // 32'h05857537;
    ram_cell[     698] = 32'h0;  // 32'h2543b00f;
    ram_cell[     699] = 32'h0;  // 32'he7ec8937;
    ram_cell[     700] = 32'h0;  // 32'he432af5b;
    ram_cell[     701] = 32'h0;  // 32'h626a84ed;
    ram_cell[     702] = 32'h0;  // 32'he93a0016;
    ram_cell[     703] = 32'h0;  // 32'hb11d8337;
    ram_cell[     704] = 32'h0;  // 32'ha3759458;
    ram_cell[     705] = 32'h0;  // 32'h0870be82;
    ram_cell[     706] = 32'h0;  // 32'h3fe623d9;
    ram_cell[     707] = 32'h0;  // 32'hecdd0736;
    ram_cell[     708] = 32'h0;  // 32'h1671a899;
    ram_cell[     709] = 32'h0;  // 32'h85eea8f1;
    ram_cell[     710] = 32'h0;  // 32'h2279d15d;
    ram_cell[     711] = 32'h0;  // 32'h2e3cd907;
    ram_cell[     712] = 32'h0;  // 32'hc895e952;
    ram_cell[     713] = 32'h0;  // 32'h3510b00a;
    ram_cell[     714] = 32'h0;  // 32'hd147f807;
    ram_cell[     715] = 32'h0;  // 32'h17905740;
    ram_cell[     716] = 32'h0;  // 32'hd85981a6;
    ram_cell[     717] = 32'h0;  // 32'h83229e2a;
    ram_cell[     718] = 32'h0;  // 32'hb41b6b57;
    ram_cell[     719] = 32'h0;  // 32'h337e804b;
    ram_cell[     720] = 32'h0;  // 32'h55b96848;
    ram_cell[     721] = 32'h0;  // 32'hdcdf9b05;
    ram_cell[     722] = 32'h0;  // 32'h83f02f73;
    ram_cell[     723] = 32'h0;  // 32'h68be2847;
    ram_cell[     724] = 32'h0;  // 32'he8fff38e;
    ram_cell[     725] = 32'h0;  // 32'hedc940b4;
    ram_cell[     726] = 32'h0;  // 32'hb7e24249;
    ram_cell[     727] = 32'h0;  // 32'h342f1359;
    ram_cell[     728] = 32'h0;  // 32'hbff490d5;
    ram_cell[     729] = 32'h0;  // 32'ha33b2fe5;
    ram_cell[     730] = 32'h0;  // 32'h581888a0;
    ram_cell[     731] = 32'h0;  // 32'he364a1d3;
    ram_cell[     732] = 32'h0;  // 32'hb5ec1481;
    ram_cell[     733] = 32'h0;  // 32'hf2050513;
    ram_cell[     734] = 32'h0;  // 32'ha514f865;
    ram_cell[     735] = 32'h0;  // 32'hce86efc6;
    ram_cell[     736] = 32'h0;  // 32'hd4624901;
    ram_cell[     737] = 32'h0;  // 32'hf83c8be2;
    ram_cell[     738] = 32'h0;  // 32'h00ee5d69;
    ram_cell[     739] = 32'h0;  // 32'hb28753af;
    ram_cell[     740] = 32'h0;  // 32'h7f9bcfac;
    ram_cell[     741] = 32'h0;  // 32'h690035bd;
    ram_cell[     742] = 32'h0;  // 32'h0622c05f;
    ram_cell[     743] = 32'h0;  // 32'hf29487cb;
    ram_cell[     744] = 32'h0;  // 32'h0aa96f82;
    ram_cell[     745] = 32'h0;  // 32'hf3b63760;
    ram_cell[     746] = 32'h0;  // 32'h3a34af25;
    ram_cell[     747] = 32'h0;  // 32'hc5b05d90;
    ram_cell[     748] = 32'h0;  // 32'h291ce427;
    ram_cell[     749] = 32'h0;  // 32'had9b8877;
    ram_cell[     750] = 32'h0;  // 32'h90668763;
    ram_cell[     751] = 32'h0;  // 32'hec696399;
    ram_cell[     752] = 32'h0;  // 32'h5249aa11;
    ram_cell[     753] = 32'h0;  // 32'h8e2d97e0;
    ram_cell[     754] = 32'h0;  // 32'h4136be47;
    ram_cell[     755] = 32'h0;  // 32'h8d2c8896;
    ram_cell[     756] = 32'h0;  // 32'h0cbe47cb;
    ram_cell[     757] = 32'h0;  // 32'h4fbed163;
    ram_cell[     758] = 32'h0;  // 32'h99f8788c;
    ram_cell[     759] = 32'h0;  // 32'h0cf1e2c4;
    ram_cell[     760] = 32'h0;  // 32'hc91adcb2;
    ram_cell[     761] = 32'h0;  // 32'h97bb38a9;
    ram_cell[     762] = 32'h0;  // 32'h1581cd6d;
    ram_cell[     763] = 32'h0;  // 32'hfb591d42;
    ram_cell[     764] = 32'h0;  // 32'h55ed3feb;
    ram_cell[     765] = 32'h0;  // 32'h94f18064;
    ram_cell[     766] = 32'h0;  // 32'h3d312a9f;
    ram_cell[     767] = 32'h0;  // 32'h844094b5;
    ram_cell[     768] = 32'h0;  // 32'h553ed1dd;
    ram_cell[     769] = 32'h0;  // 32'hd2197734;
    ram_cell[     770] = 32'h0;  // 32'h815dbabf;
    ram_cell[     771] = 32'h0;  // 32'hfe2537a2;
    ram_cell[     772] = 32'h0;  // 32'h75222e9b;
    ram_cell[     773] = 32'h0;  // 32'h9820a496;
    ram_cell[     774] = 32'h0;  // 32'h0ee5a81a;
    ram_cell[     775] = 32'h0;  // 32'h53a4851c;
    ram_cell[     776] = 32'h0;  // 32'h659d4bd2;
    ram_cell[     777] = 32'h0;  // 32'h513f865a;
    ram_cell[     778] = 32'h0;  // 32'h23c661c5;
    ram_cell[     779] = 32'h0;  // 32'he1af8d97;
    ram_cell[     780] = 32'h0;  // 32'hf42e45c5;
    ram_cell[     781] = 32'h0;  // 32'hdceb9045;
    ram_cell[     782] = 32'h0;  // 32'ha2f0cd8f;
    ram_cell[     783] = 32'h0;  // 32'hf77131c3;
    ram_cell[     784] = 32'h0;  // 32'h0d5a2260;
    ram_cell[     785] = 32'h0;  // 32'hc579e35b;
    ram_cell[     786] = 32'h0;  // 32'h3e3d801a;
    ram_cell[     787] = 32'h0;  // 32'h147216c5;
    ram_cell[     788] = 32'h0;  // 32'h93f77868;
    ram_cell[     789] = 32'h0;  // 32'ha52e1041;
    ram_cell[     790] = 32'h0;  // 32'h4da878ed;
    ram_cell[     791] = 32'h0;  // 32'h9126dcb5;
    ram_cell[     792] = 32'h0;  // 32'h3a697653;
    ram_cell[     793] = 32'h0;  // 32'h6991df96;
    ram_cell[     794] = 32'h0;  // 32'h0e8c0557;
    ram_cell[     795] = 32'h0;  // 32'h64b95c45;
    ram_cell[     796] = 32'h0;  // 32'hfbf7e1ac;
    ram_cell[     797] = 32'h0;  // 32'h9283ae6a;
    ram_cell[     798] = 32'h0;  // 32'h38fa03d6;
    ram_cell[     799] = 32'h0;  // 32'hc4b009b0;
    ram_cell[     800] = 32'h0;  // 32'he29c470a;
    ram_cell[     801] = 32'h0;  // 32'h14fdd57f;
    ram_cell[     802] = 32'h0;  // 32'hd0c21f19;
    ram_cell[     803] = 32'h0;  // 32'hd298cc06;
    ram_cell[     804] = 32'h0;  // 32'hd4553262;
    ram_cell[     805] = 32'h0;  // 32'h82bab81f;
    ram_cell[     806] = 32'h0;  // 32'hdcd3f55c;
    ram_cell[     807] = 32'h0;  // 32'h088e9cb3;
    ram_cell[     808] = 32'h0;  // 32'h115e75c4;
    ram_cell[     809] = 32'h0;  // 32'h25d73312;
    ram_cell[     810] = 32'h0;  // 32'h8a52380d;
    ram_cell[     811] = 32'h0;  // 32'h16387b1e;
    ram_cell[     812] = 32'h0;  // 32'h25a1a934;
    ram_cell[     813] = 32'h0;  // 32'h62ac3b34;
    ram_cell[     814] = 32'h0;  // 32'h0198aed5;
    ram_cell[     815] = 32'h0;  // 32'h0cd345e8;
    ram_cell[     816] = 32'h0;  // 32'hb2fbfff9;
    ram_cell[     817] = 32'h0;  // 32'h7855ee16;
    ram_cell[     818] = 32'h0;  // 32'hca1ef591;
    ram_cell[     819] = 32'h0;  // 32'h2027734d;
    ram_cell[     820] = 32'h0;  // 32'h364b7383;
    ram_cell[     821] = 32'h0;  // 32'he147bdec;
    ram_cell[     822] = 32'h0;  // 32'ha51220cc;
    ram_cell[     823] = 32'h0;  // 32'h2817b15f;
    ram_cell[     824] = 32'h0;  // 32'hcb661be7;
    ram_cell[     825] = 32'h0;  // 32'h7224ddfe;
    ram_cell[     826] = 32'h0;  // 32'h3a129fbf;
    ram_cell[     827] = 32'h0;  // 32'hd9d558e8;
    ram_cell[     828] = 32'h0;  // 32'h485bc579;
    ram_cell[     829] = 32'h0;  // 32'hf79f4db8;
    ram_cell[     830] = 32'h0;  // 32'ha0cfebdc;
    ram_cell[     831] = 32'h0;  // 32'hb127957d;
    ram_cell[     832] = 32'h0;  // 32'hf4959413;
    ram_cell[     833] = 32'h0;  // 32'hab8b38c4;
    ram_cell[     834] = 32'h0;  // 32'h7bd21d04;
    ram_cell[     835] = 32'h0;  // 32'h1585a9e8;
    ram_cell[     836] = 32'h0;  // 32'hcd4ba194;
    ram_cell[     837] = 32'h0;  // 32'heeab9c80;
    ram_cell[     838] = 32'h0;  // 32'h35343dff;
    ram_cell[     839] = 32'h0;  // 32'h4aa8ae80;
    ram_cell[     840] = 32'h0;  // 32'h1fa59870;
    ram_cell[     841] = 32'h0;  // 32'hb9566dc5;
    ram_cell[     842] = 32'h0;  // 32'hd97bcfca;
    ram_cell[     843] = 32'h0;  // 32'h5163215d;
    ram_cell[     844] = 32'h0;  // 32'h35b8205f;
    ram_cell[     845] = 32'h0;  // 32'h032a0e27;
    ram_cell[     846] = 32'h0;  // 32'ha9a8c4e0;
    ram_cell[     847] = 32'h0;  // 32'h636a90b7;
    ram_cell[     848] = 32'h0;  // 32'haf85b068;
    ram_cell[     849] = 32'h0;  // 32'h98b48904;
    ram_cell[     850] = 32'h0;  // 32'he8df67e3;
    ram_cell[     851] = 32'h0;  // 32'hc92fcfd4;
    ram_cell[     852] = 32'h0;  // 32'hea672fcd;
    ram_cell[     853] = 32'h0;  // 32'hbaa19f3f;
    ram_cell[     854] = 32'h0;  // 32'hd8a25d32;
    ram_cell[     855] = 32'h0;  // 32'h3057d1cc;
    ram_cell[     856] = 32'h0;  // 32'hf271ad3d;
    ram_cell[     857] = 32'h0;  // 32'h890ac7cc;
    ram_cell[     858] = 32'h0;  // 32'hc861fb4a;
    ram_cell[     859] = 32'h0;  // 32'hbcd8e381;
    ram_cell[     860] = 32'h0;  // 32'h621584c8;
    ram_cell[     861] = 32'h0;  // 32'h6d35b5f2;
    ram_cell[     862] = 32'h0;  // 32'h01266247;
    ram_cell[     863] = 32'h0;  // 32'ha7ed91a3;
    ram_cell[     864] = 32'h0;  // 32'ha53976e6;
    ram_cell[     865] = 32'h0;  // 32'h830eacce;
    ram_cell[     866] = 32'h0;  // 32'h16eafccd;
    ram_cell[     867] = 32'h0;  // 32'hb7b48ceb;
    ram_cell[     868] = 32'h0;  // 32'heeecea55;
    ram_cell[     869] = 32'h0;  // 32'h6db8a6eb;
    ram_cell[     870] = 32'h0;  // 32'h8986e54c;
    ram_cell[     871] = 32'h0;  // 32'hdfd64ae5;
    ram_cell[     872] = 32'h0;  // 32'h3d1ef428;
    ram_cell[     873] = 32'h0;  // 32'hb3f6c204;
    ram_cell[     874] = 32'h0;  // 32'hf50fba94;
    ram_cell[     875] = 32'h0;  // 32'h6319efea;
    ram_cell[     876] = 32'h0;  // 32'h72e34646;
    ram_cell[     877] = 32'h0;  // 32'habd6ac4f;
    ram_cell[     878] = 32'h0;  // 32'h69ecacf9;
    ram_cell[     879] = 32'h0;  // 32'h8e9851fc;
    ram_cell[     880] = 32'h0;  // 32'h5db2bc11;
    ram_cell[     881] = 32'h0;  // 32'h433216b2;
    ram_cell[     882] = 32'h0;  // 32'h8fda39ab;
    ram_cell[     883] = 32'h0;  // 32'h83ce1366;
    ram_cell[     884] = 32'h0;  // 32'hfab76c7f;
    ram_cell[     885] = 32'h0;  // 32'h90f3738b;
    ram_cell[     886] = 32'h0;  // 32'h58d2e5d8;
    ram_cell[     887] = 32'h0;  // 32'ha9d2f9e2;
    ram_cell[     888] = 32'h0;  // 32'hb5d4b5e4;
    ram_cell[     889] = 32'h0;  // 32'hd8d58507;
    ram_cell[     890] = 32'h0;  // 32'hb0fab1f2;
    ram_cell[     891] = 32'h0;  // 32'h8f07d5c2;
    ram_cell[     892] = 32'h0;  // 32'h2dcbf480;
    ram_cell[     893] = 32'h0;  // 32'h9b8344e5;
    ram_cell[     894] = 32'h0;  // 32'h5678282b;
    ram_cell[     895] = 32'h0;  // 32'h7d600dc9;
    ram_cell[     896] = 32'h0;  // 32'hc5a2d79d;
    ram_cell[     897] = 32'h0;  // 32'h6a89f9ff;
    ram_cell[     898] = 32'h0;  // 32'hcd6f14cb;
    ram_cell[     899] = 32'h0;  // 32'h6c5bdab8;
    ram_cell[     900] = 32'h0;  // 32'he86fa1c7;
    ram_cell[     901] = 32'h0;  // 32'h7da07d8e;
    ram_cell[     902] = 32'h0;  // 32'h3c7d0da5;
    ram_cell[     903] = 32'h0;  // 32'h1cb7bf52;
    ram_cell[     904] = 32'h0;  // 32'hd708db1d;
    ram_cell[     905] = 32'h0;  // 32'hbb4cdd0b;
    ram_cell[     906] = 32'h0;  // 32'hb3123b0e;
    ram_cell[     907] = 32'h0;  // 32'hbb8de5d0;
    ram_cell[     908] = 32'h0;  // 32'h6fc337fd;
    ram_cell[     909] = 32'h0;  // 32'ha7f0bec4;
    ram_cell[     910] = 32'h0;  // 32'h9dd4259a;
    ram_cell[     911] = 32'h0;  // 32'haece1e30;
    ram_cell[     912] = 32'h0;  // 32'ha0d75638;
    ram_cell[     913] = 32'h0;  // 32'he2549db3;
    ram_cell[     914] = 32'h0;  // 32'h7f4b0406;
    ram_cell[     915] = 32'h0;  // 32'h7e75d732;
    ram_cell[     916] = 32'h0;  // 32'h93c2b607;
    ram_cell[     917] = 32'h0;  // 32'h9ae90142;
    ram_cell[     918] = 32'h0;  // 32'hc70d94ad;
    ram_cell[     919] = 32'h0;  // 32'hfeb97c15;
    ram_cell[     920] = 32'h0;  // 32'hfffbf4f1;
    ram_cell[     921] = 32'h0;  // 32'h4937fa3c;
    ram_cell[     922] = 32'h0;  // 32'h230f0d44;
    ram_cell[     923] = 32'h0;  // 32'h221dbdd7;
    ram_cell[     924] = 32'h0;  // 32'h717b744e;
    ram_cell[     925] = 32'h0;  // 32'heb1f476a;
    ram_cell[     926] = 32'h0;  // 32'hd6a162f0;
    ram_cell[     927] = 32'h0;  // 32'hd3b52438;
    ram_cell[     928] = 32'h0;  // 32'hcafcc562;
    ram_cell[     929] = 32'h0;  // 32'h46e8ccb2;
    ram_cell[     930] = 32'h0;  // 32'h3ff54461;
    ram_cell[     931] = 32'h0;  // 32'hd6fba0ce;
    ram_cell[     932] = 32'h0;  // 32'h7299d0e9;
    ram_cell[     933] = 32'h0;  // 32'h69fb5fa4;
    ram_cell[     934] = 32'h0;  // 32'ha74e4518;
    ram_cell[     935] = 32'h0;  // 32'h5b403edd;
    ram_cell[     936] = 32'h0;  // 32'h2fd2ed0e;
    ram_cell[     937] = 32'h0;  // 32'h98916255;
    ram_cell[     938] = 32'h0;  // 32'h17d4e081;
    ram_cell[     939] = 32'h0;  // 32'h2a3b56fe;
    ram_cell[     940] = 32'h0;  // 32'hee32d707;
    ram_cell[     941] = 32'h0;  // 32'h28aac570;
    ram_cell[     942] = 32'h0;  // 32'h0242096b;
    ram_cell[     943] = 32'h0;  // 32'h0558dec8;
    ram_cell[     944] = 32'h0;  // 32'h24e868fc;
    ram_cell[     945] = 32'h0;  // 32'h6ccf8094;
    ram_cell[     946] = 32'h0;  // 32'hfb9b377c;
    ram_cell[     947] = 32'h0;  // 32'hc10cbff2;
    ram_cell[     948] = 32'h0;  // 32'h5942c01f;
    ram_cell[     949] = 32'h0;  // 32'h3c8fcefa;
    ram_cell[     950] = 32'h0;  // 32'h6f23602d;
    ram_cell[     951] = 32'h0;  // 32'h039fee0b;
    ram_cell[     952] = 32'h0;  // 32'hd29b6dd3;
    ram_cell[     953] = 32'h0;  // 32'h33db9950;
    ram_cell[     954] = 32'h0;  // 32'h75cf6b1d;
    ram_cell[     955] = 32'h0;  // 32'h690b1fd1;
    ram_cell[     956] = 32'h0;  // 32'hd6ea7547;
    ram_cell[     957] = 32'h0;  // 32'hda752168;
    ram_cell[     958] = 32'h0;  // 32'h38a96553;
    ram_cell[     959] = 32'h0;  // 32'h18580eb5;
    ram_cell[     960] = 32'h0;  // 32'h6757f17a;
    ram_cell[     961] = 32'h0;  // 32'hb71e9472;
    ram_cell[     962] = 32'h0;  // 32'hf26dc669;
    ram_cell[     963] = 32'h0;  // 32'h8586c349;
    ram_cell[     964] = 32'h0;  // 32'h39792f0b;
    ram_cell[     965] = 32'h0;  // 32'h0a9f1a1c;
    ram_cell[     966] = 32'h0;  // 32'hda8d4d35;
    ram_cell[     967] = 32'h0;  // 32'h80255b74;
    ram_cell[     968] = 32'h0;  // 32'hc1acc2ea;
    ram_cell[     969] = 32'h0;  // 32'hbf523e20;
    ram_cell[     970] = 32'h0;  // 32'h29798fcd;
    ram_cell[     971] = 32'h0;  // 32'h150bad01;
    ram_cell[     972] = 32'h0;  // 32'hf8663f30;
    ram_cell[     973] = 32'h0;  // 32'h5e7ddfbd;
    ram_cell[     974] = 32'h0;  // 32'hd35ce0bf;
    ram_cell[     975] = 32'h0;  // 32'h8d5b9d6f;
    ram_cell[     976] = 32'h0;  // 32'h627cbb58;
    ram_cell[     977] = 32'h0;  // 32'hf4a7bc74;
    ram_cell[     978] = 32'h0;  // 32'h020f234e;
    ram_cell[     979] = 32'h0;  // 32'hd4d9afa2;
    ram_cell[     980] = 32'h0;  // 32'hf507fefe;
    ram_cell[     981] = 32'h0;  // 32'h024650c4;
    ram_cell[     982] = 32'h0;  // 32'hd1d23c0c;
    ram_cell[     983] = 32'h0;  // 32'hce099e08;
    ram_cell[     984] = 32'h0;  // 32'h0c3b43fa;
    ram_cell[     985] = 32'h0;  // 32'hd340df0c;
    ram_cell[     986] = 32'h0;  // 32'hb7a3cec1;
    ram_cell[     987] = 32'h0;  // 32'h34a086db;
    ram_cell[     988] = 32'h0;  // 32'h7e157fad;
    ram_cell[     989] = 32'h0;  // 32'h3680c542;
    ram_cell[     990] = 32'h0;  // 32'h19f3c878;
    ram_cell[     991] = 32'h0;  // 32'h78f18681;
    ram_cell[     992] = 32'h0;  // 32'he98b9859;
    ram_cell[     993] = 32'h0;  // 32'h6b6088cf;
    ram_cell[     994] = 32'h0;  // 32'ha258a0d5;
    ram_cell[     995] = 32'h0;  // 32'he9b44659;
    ram_cell[     996] = 32'h0;  // 32'h406fbaa7;
    ram_cell[     997] = 32'h0;  // 32'hec74dfbd;
    ram_cell[     998] = 32'h0;  // 32'had4d135d;
    ram_cell[     999] = 32'h0;  // 32'h17b4dce0;
    ram_cell[    1000] = 32'h0;  // 32'h02b5252c;
    ram_cell[    1001] = 32'h0;  // 32'hd96e885c;
    ram_cell[    1002] = 32'h0;  // 32'h1995c928;
    ram_cell[    1003] = 32'h0;  // 32'h4ced7c99;
    ram_cell[    1004] = 32'h0;  // 32'h9a9d6ce9;
    ram_cell[    1005] = 32'h0;  // 32'h56664355;
    ram_cell[    1006] = 32'h0;  // 32'hbfd8b9b2;
    ram_cell[    1007] = 32'h0;  // 32'h53602ad4;
    ram_cell[    1008] = 32'h0;  // 32'hcab43933;
    ram_cell[    1009] = 32'h0;  // 32'hce7cda89;
    ram_cell[    1010] = 32'h0;  // 32'hea9ca55c;
    ram_cell[    1011] = 32'h0;  // 32'h8ebe07f8;
    ram_cell[    1012] = 32'h0;  // 32'ha842bf3d;
    ram_cell[    1013] = 32'h0;  // 32'hd4a50a10;
    ram_cell[    1014] = 32'h0;  // 32'h72912e2c;
    ram_cell[    1015] = 32'h0;  // 32'he2b6a67c;
    ram_cell[    1016] = 32'h0;  // 32'hf815a8f5;
    ram_cell[    1017] = 32'h0;  // 32'h2fdf62d0;
    ram_cell[    1018] = 32'h0;  // 32'h2586ccc2;
    ram_cell[    1019] = 32'h0;  // 32'hfe11036c;
    ram_cell[    1020] = 32'h0;  // 32'h175d798a;
    ram_cell[    1021] = 32'h0;  // 32'hedc99f11;
    ram_cell[    1022] = 32'h0;  // 32'h55d55b17;
    ram_cell[    1023] = 32'h0;  // 32'hc84a05f0;
    // src matrix A
    ram_cell[    1024] = 32'h3c1ce27a;
    ram_cell[    1025] = 32'hc16c2315;
    ram_cell[    1026] = 32'h010512e5;
    ram_cell[    1027] = 32'h5153fe35;
    ram_cell[    1028] = 32'hd3299bb4;
    ram_cell[    1029] = 32'hc46c8baf;
    ram_cell[    1030] = 32'hf3ad1690;
    ram_cell[    1031] = 32'h19c7342f;
    ram_cell[    1032] = 32'hf3d01cfe;
    ram_cell[    1033] = 32'hefa138ca;
    ram_cell[    1034] = 32'h2a52745f;
    ram_cell[    1035] = 32'h675d92c6;
    ram_cell[    1036] = 32'h967342d7;
    ram_cell[    1037] = 32'h9d6fdb43;
    ram_cell[    1038] = 32'hd29630f0;
    ram_cell[    1039] = 32'h11326693;
    ram_cell[    1040] = 32'hb82486f1;
    ram_cell[    1041] = 32'h79e6f940;
    ram_cell[    1042] = 32'h22634391;
    ram_cell[    1043] = 32'h490481e3;
    ram_cell[    1044] = 32'hbd4faf1d;
    ram_cell[    1045] = 32'h1ab69812;
    ram_cell[    1046] = 32'h911801cb;
    ram_cell[    1047] = 32'h41c63f24;
    ram_cell[    1048] = 32'h9bc806dd;
    ram_cell[    1049] = 32'hf0554829;
    ram_cell[    1050] = 32'h816b6c7b;
    ram_cell[    1051] = 32'h58d2a01c;
    ram_cell[    1052] = 32'h7bfde9d9;
    ram_cell[    1053] = 32'haed066c9;
    ram_cell[    1054] = 32'hdc9f945f;
    ram_cell[    1055] = 32'h6165177c;
    ram_cell[    1056] = 32'h6f79c1fa;
    ram_cell[    1057] = 32'h744b2a0f;
    ram_cell[    1058] = 32'h229a055a;
    ram_cell[    1059] = 32'h3bf67cc0;
    ram_cell[    1060] = 32'hd4e315c2;
    ram_cell[    1061] = 32'had7c5f84;
    ram_cell[    1062] = 32'h07a5932a;
    ram_cell[    1063] = 32'h2e34a6f3;
    ram_cell[    1064] = 32'hc3584403;
    ram_cell[    1065] = 32'h52af0c2b;
    ram_cell[    1066] = 32'h01418069;
    ram_cell[    1067] = 32'h06326b3f;
    ram_cell[    1068] = 32'hbdb4348a;
    ram_cell[    1069] = 32'h70553be7;
    ram_cell[    1070] = 32'hb50b7494;
    ram_cell[    1071] = 32'h77e42961;
    ram_cell[    1072] = 32'hd34cf638;
    ram_cell[    1073] = 32'h88a054ca;
    ram_cell[    1074] = 32'h1e2e95e6;
    ram_cell[    1075] = 32'heef1a825;
    ram_cell[    1076] = 32'h3f84255c;
    ram_cell[    1077] = 32'h403e7539;
    ram_cell[    1078] = 32'h4c773097;
    ram_cell[    1079] = 32'ha99d9291;
    ram_cell[    1080] = 32'h7fd0ffb9;
    ram_cell[    1081] = 32'h73cb59c0;
    ram_cell[    1082] = 32'h5d6e756a;
    ram_cell[    1083] = 32'hf45a9504;
    ram_cell[    1084] = 32'h015c1113;
    ram_cell[    1085] = 32'h0570610a;
    ram_cell[    1086] = 32'h0ec576b9;
    ram_cell[    1087] = 32'h83b1db2f;
    ram_cell[    1088] = 32'ha8e77732;
    ram_cell[    1089] = 32'h8eb8f7e5;
    ram_cell[    1090] = 32'hcf0bdbba;
    ram_cell[    1091] = 32'h6027532f;
    ram_cell[    1092] = 32'h0007ee23;
    ram_cell[    1093] = 32'h1b1f3908;
    ram_cell[    1094] = 32'h0eceec87;
    ram_cell[    1095] = 32'h674c5f39;
    ram_cell[    1096] = 32'h2bd39773;
    ram_cell[    1097] = 32'h0942bc0d;
    ram_cell[    1098] = 32'h0e0b2228;
    ram_cell[    1099] = 32'h618751e3;
    ram_cell[    1100] = 32'h6ce97d51;
    ram_cell[    1101] = 32'hda6aa42a;
    ram_cell[    1102] = 32'h95c59082;
    ram_cell[    1103] = 32'hcf593dea;
    ram_cell[    1104] = 32'h0481ae90;
    ram_cell[    1105] = 32'h4898d693;
    ram_cell[    1106] = 32'h79f593f8;
    ram_cell[    1107] = 32'hd69bf96c;
    ram_cell[    1108] = 32'hf61b815a;
    ram_cell[    1109] = 32'h75fafb6a;
    ram_cell[    1110] = 32'h00e1b1e7;
    ram_cell[    1111] = 32'h85e43da5;
    ram_cell[    1112] = 32'h006d6700;
    ram_cell[    1113] = 32'hc55aedf9;
    ram_cell[    1114] = 32'h438b57b0;
    ram_cell[    1115] = 32'hf92cefd1;
    ram_cell[    1116] = 32'h5b9ae8b0;
    ram_cell[    1117] = 32'hf0564d1a;
    ram_cell[    1118] = 32'hc87ecb88;
    ram_cell[    1119] = 32'hc767b390;
    ram_cell[    1120] = 32'haae0d53e;
    ram_cell[    1121] = 32'hd29905a4;
    ram_cell[    1122] = 32'h112617ba;
    ram_cell[    1123] = 32'hdbff510b;
    ram_cell[    1124] = 32'hcd1969af;
    ram_cell[    1125] = 32'h7ec89f0d;
    ram_cell[    1126] = 32'h60625e7d;
    ram_cell[    1127] = 32'h16e7c7eb;
    ram_cell[    1128] = 32'hc3c9139b;
    ram_cell[    1129] = 32'h99eb9006;
    ram_cell[    1130] = 32'he52ecf6d;
    ram_cell[    1131] = 32'h88d6ed47;
    ram_cell[    1132] = 32'h8095cfe2;
    ram_cell[    1133] = 32'h7211bbb4;
    ram_cell[    1134] = 32'h6bff3ed7;
    ram_cell[    1135] = 32'he452a0a7;
    ram_cell[    1136] = 32'hbaa01b27;
    ram_cell[    1137] = 32'haee166b9;
    ram_cell[    1138] = 32'h0ccd756f;
    ram_cell[    1139] = 32'h864b3186;
    ram_cell[    1140] = 32'h2d60ed18;
    ram_cell[    1141] = 32'h996abc73;
    ram_cell[    1142] = 32'h310abab2;
    ram_cell[    1143] = 32'hb32a55c0;
    ram_cell[    1144] = 32'h9ab93bdf;
    ram_cell[    1145] = 32'h195be18e;
    ram_cell[    1146] = 32'h3265266a;
    ram_cell[    1147] = 32'h5687917c;
    ram_cell[    1148] = 32'heea483f0;
    ram_cell[    1149] = 32'ha9b736b4;
    ram_cell[    1150] = 32'h063850ed;
    ram_cell[    1151] = 32'hb2817ebe;
    ram_cell[    1152] = 32'ha1f937f4;
    ram_cell[    1153] = 32'he4d03c78;
    ram_cell[    1154] = 32'h8d9a175e;
    ram_cell[    1155] = 32'haedbd0be;
    ram_cell[    1156] = 32'h8d0e48ee;
    ram_cell[    1157] = 32'h3967640a;
    ram_cell[    1158] = 32'h18560cfd;
    ram_cell[    1159] = 32'h9636f4b7;
    ram_cell[    1160] = 32'hff9e3ffe;
    ram_cell[    1161] = 32'h1ba4d317;
    ram_cell[    1162] = 32'h5721f0aa;
    ram_cell[    1163] = 32'h9fbc1647;
    ram_cell[    1164] = 32'h5021519d;
    ram_cell[    1165] = 32'h972eb2de;
    ram_cell[    1166] = 32'hf689a928;
    ram_cell[    1167] = 32'h494f1c28;
    ram_cell[    1168] = 32'hf246365b;
    ram_cell[    1169] = 32'h908cb105;
    ram_cell[    1170] = 32'h6b4aeccc;
    ram_cell[    1171] = 32'h44d0890b;
    ram_cell[    1172] = 32'hf1e2761f;
    ram_cell[    1173] = 32'hbe14fbcc;
    ram_cell[    1174] = 32'h97c62599;
    ram_cell[    1175] = 32'hbd87700f;
    ram_cell[    1176] = 32'h9d54a559;
    ram_cell[    1177] = 32'h46f2b4a0;
    ram_cell[    1178] = 32'hb5d6e358;
    ram_cell[    1179] = 32'h8c3c5965;
    ram_cell[    1180] = 32'ha862bd03;
    ram_cell[    1181] = 32'hd58a1958;
    ram_cell[    1182] = 32'h23775bfd;
    ram_cell[    1183] = 32'h4206daeb;
    ram_cell[    1184] = 32'h68b2f6dc;
    ram_cell[    1185] = 32'h0b35eeea;
    ram_cell[    1186] = 32'hf3cc76f3;
    ram_cell[    1187] = 32'h59318f1e;
    ram_cell[    1188] = 32'hdf5292b1;
    ram_cell[    1189] = 32'ha642648e;
    ram_cell[    1190] = 32'h02ea30dc;
    ram_cell[    1191] = 32'h0b7d2e33;
    ram_cell[    1192] = 32'h862f72ca;
    ram_cell[    1193] = 32'hc49020c4;
    ram_cell[    1194] = 32'h6a6550b0;
    ram_cell[    1195] = 32'hb43ea9ff;
    ram_cell[    1196] = 32'h8198b117;
    ram_cell[    1197] = 32'hce9dd383;
    ram_cell[    1198] = 32'h3d89b7e0;
    ram_cell[    1199] = 32'haf49c7b1;
    ram_cell[    1200] = 32'h5467dcfe;
    ram_cell[    1201] = 32'hdfe156cb;
    ram_cell[    1202] = 32'he13126c1;
    ram_cell[    1203] = 32'h25c7f001;
    ram_cell[    1204] = 32'h8e0418ad;
    ram_cell[    1205] = 32'hc5692372;
    ram_cell[    1206] = 32'h0a2b7eb2;
    ram_cell[    1207] = 32'h4bbc0261;
    ram_cell[    1208] = 32'h9d1e480e;
    ram_cell[    1209] = 32'he755896b;
    ram_cell[    1210] = 32'ha3ccdb7e;
    ram_cell[    1211] = 32'h0372f149;
    ram_cell[    1212] = 32'he5dfbcfd;
    ram_cell[    1213] = 32'h19c2b472;
    ram_cell[    1214] = 32'h9f6b8491;
    ram_cell[    1215] = 32'h7a17f1ec;
    ram_cell[    1216] = 32'hdb0e5020;
    ram_cell[    1217] = 32'hf14fb157;
    ram_cell[    1218] = 32'hd1b54321;
    ram_cell[    1219] = 32'h892f608d;
    ram_cell[    1220] = 32'h56d7d335;
    ram_cell[    1221] = 32'hbcb30281;
    ram_cell[    1222] = 32'h83f09819;
    ram_cell[    1223] = 32'hc1915a0d;
    ram_cell[    1224] = 32'h846a47d6;
    ram_cell[    1225] = 32'hd5555e73;
    ram_cell[    1226] = 32'haf7fc2b1;
    ram_cell[    1227] = 32'h582e6d42;
    ram_cell[    1228] = 32'h1bb72851;
    ram_cell[    1229] = 32'hb1426ada;
    ram_cell[    1230] = 32'h7c478191;
    ram_cell[    1231] = 32'he40e9497;
    ram_cell[    1232] = 32'heb033c17;
    ram_cell[    1233] = 32'hb0f954b5;
    ram_cell[    1234] = 32'h61413d5a;
    ram_cell[    1235] = 32'h0ef6b989;
    ram_cell[    1236] = 32'h0a5db9ea;
    ram_cell[    1237] = 32'ha665f5b2;
    ram_cell[    1238] = 32'h63cca392;
    ram_cell[    1239] = 32'h94a3f7e0;
    ram_cell[    1240] = 32'hce1a41fd;
    ram_cell[    1241] = 32'hd65c254e;
    ram_cell[    1242] = 32'hbc4a5bbd;
    ram_cell[    1243] = 32'h0e0fd07d;
    ram_cell[    1244] = 32'h0b629207;
    ram_cell[    1245] = 32'hdaf7b884;
    ram_cell[    1246] = 32'h09784ab0;
    ram_cell[    1247] = 32'h136f4aca;
    ram_cell[    1248] = 32'h3adfb06b;
    ram_cell[    1249] = 32'h0bce999f;
    ram_cell[    1250] = 32'h15148fe5;
    ram_cell[    1251] = 32'h6fa1fbc3;
    ram_cell[    1252] = 32'h605e5934;
    ram_cell[    1253] = 32'hde061908;
    ram_cell[    1254] = 32'he3b73c1b;
    ram_cell[    1255] = 32'ha7b6273c;
    ram_cell[    1256] = 32'hefe2d3e7;
    ram_cell[    1257] = 32'h360a989d;
    ram_cell[    1258] = 32'h94353e71;
    ram_cell[    1259] = 32'h1de1993f;
    ram_cell[    1260] = 32'h801d9d91;
    ram_cell[    1261] = 32'hb696f1b0;
    ram_cell[    1262] = 32'h5b3c7b36;
    ram_cell[    1263] = 32'h51498d5b;
    ram_cell[    1264] = 32'hc02eceae;
    ram_cell[    1265] = 32'hd7514cae;
    ram_cell[    1266] = 32'h5d726ba8;
    ram_cell[    1267] = 32'h60abd90c;
    ram_cell[    1268] = 32'h136d8e51;
    ram_cell[    1269] = 32'ha42d1e55;
    ram_cell[    1270] = 32'hc8e87564;
    ram_cell[    1271] = 32'h0a27b4ab;
    ram_cell[    1272] = 32'hb832c299;
    ram_cell[    1273] = 32'h8b42e1ed;
    ram_cell[    1274] = 32'hed5add2d;
    ram_cell[    1275] = 32'h7e48f341;
    ram_cell[    1276] = 32'hc8bccc95;
    ram_cell[    1277] = 32'h437dd432;
    ram_cell[    1278] = 32'h92b5cdfa;
    ram_cell[    1279] = 32'h79e77023;
    ram_cell[    1280] = 32'h5e6a212c;
    ram_cell[    1281] = 32'h06976990;
    ram_cell[    1282] = 32'h51e65627;
    ram_cell[    1283] = 32'h896a9f9f;
    ram_cell[    1284] = 32'he51f4da5;
    ram_cell[    1285] = 32'he0f48e62;
    ram_cell[    1286] = 32'h973f7f40;
    ram_cell[    1287] = 32'h81059168;
    ram_cell[    1288] = 32'ha1d39da4;
    ram_cell[    1289] = 32'hc4ec7576;
    ram_cell[    1290] = 32'hf7ca072b;
    ram_cell[    1291] = 32'h70789b7c;
    ram_cell[    1292] = 32'h3bf63ecc;
    ram_cell[    1293] = 32'h574de49a;
    ram_cell[    1294] = 32'h5d60227d;
    ram_cell[    1295] = 32'h4ddf6c17;
    ram_cell[    1296] = 32'h185a93f2;
    ram_cell[    1297] = 32'h5c9184f8;
    ram_cell[    1298] = 32'hacb5b075;
    ram_cell[    1299] = 32'h1909b70f;
    ram_cell[    1300] = 32'h8574c6d0;
    ram_cell[    1301] = 32'h5fe8093b;
    ram_cell[    1302] = 32'hbde69267;
    ram_cell[    1303] = 32'h8957df00;
    ram_cell[    1304] = 32'hb9d28283;
    ram_cell[    1305] = 32'h4ed82b16;
    ram_cell[    1306] = 32'he831ff39;
    ram_cell[    1307] = 32'hea5f0220;
    ram_cell[    1308] = 32'haa245f99;
    ram_cell[    1309] = 32'he22dd40e;
    ram_cell[    1310] = 32'h23756a4e;
    ram_cell[    1311] = 32'h19d82a31;
    ram_cell[    1312] = 32'hb7ad992b;
    ram_cell[    1313] = 32'hefb2b5ba;
    ram_cell[    1314] = 32'haa98bbdf;
    ram_cell[    1315] = 32'h917b9e37;
    ram_cell[    1316] = 32'h153a95c8;
    ram_cell[    1317] = 32'h3df327f0;
    ram_cell[    1318] = 32'hbb1931b9;
    ram_cell[    1319] = 32'h9336913a;
    ram_cell[    1320] = 32'h809dc97b;
    ram_cell[    1321] = 32'h658dd266;
    ram_cell[    1322] = 32'h2fe67dc8;
    ram_cell[    1323] = 32'h81cd2111;
    ram_cell[    1324] = 32'h8bf9dd25;
    ram_cell[    1325] = 32'hd1c1366b;
    ram_cell[    1326] = 32'h09243a2d;
    ram_cell[    1327] = 32'hb2993d8e;
    ram_cell[    1328] = 32'h05b4d60d;
    ram_cell[    1329] = 32'hb1cf3afb;
    ram_cell[    1330] = 32'hcdfe67ae;
    ram_cell[    1331] = 32'h04fedf70;
    ram_cell[    1332] = 32'he9650308;
    ram_cell[    1333] = 32'heca716e2;
    ram_cell[    1334] = 32'h38ea5376;
    ram_cell[    1335] = 32'h2f367c9d;
    ram_cell[    1336] = 32'hefdf96c8;
    ram_cell[    1337] = 32'hb144d4a6;
    ram_cell[    1338] = 32'habcf8dda;
    ram_cell[    1339] = 32'h859c0ebd;
    ram_cell[    1340] = 32'hcdcd4e1e;
    ram_cell[    1341] = 32'h34597ca8;
    ram_cell[    1342] = 32'h7d197bfb;
    ram_cell[    1343] = 32'ha8a549d5;
    ram_cell[    1344] = 32'h1548a57d;
    ram_cell[    1345] = 32'hef2923bd;
    ram_cell[    1346] = 32'h7ddd7f50;
    ram_cell[    1347] = 32'hd134dca4;
    ram_cell[    1348] = 32'hdea0115e;
    ram_cell[    1349] = 32'hdc7fc1cd;
    ram_cell[    1350] = 32'hb97353d3;
    ram_cell[    1351] = 32'h570f76eb;
    ram_cell[    1352] = 32'he5b2ef14;
    ram_cell[    1353] = 32'h71ba9156;
    ram_cell[    1354] = 32'hc6f0e0c9;
    ram_cell[    1355] = 32'hfb79a646;
    ram_cell[    1356] = 32'h1d2582fc;
    ram_cell[    1357] = 32'h09598344;
    ram_cell[    1358] = 32'h370c790f;
    ram_cell[    1359] = 32'hb9e12602;
    ram_cell[    1360] = 32'hce5cdebd;
    ram_cell[    1361] = 32'hd678dfc2;
    ram_cell[    1362] = 32'h00b07709;
    ram_cell[    1363] = 32'hdfa3c762;
    ram_cell[    1364] = 32'hffda0f00;
    ram_cell[    1365] = 32'h4650947a;
    ram_cell[    1366] = 32'h11dae664;
    ram_cell[    1367] = 32'h499aed73;
    ram_cell[    1368] = 32'hc82fa59d;
    ram_cell[    1369] = 32'h906548e1;
    ram_cell[    1370] = 32'h9107bf98;
    ram_cell[    1371] = 32'ha9aac440;
    ram_cell[    1372] = 32'heb5ca284;
    ram_cell[    1373] = 32'h36d32637;
    ram_cell[    1374] = 32'hc661fc02;
    ram_cell[    1375] = 32'hedda45ba;
    ram_cell[    1376] = 32'hf63e7ae6;
    ram_cell[    1377] = 32'h7cf70dcf;
    ram_cell[    1378] = 32'h3cbc053a;
    ram_cell[    1379] = 32'h8183057a;
    ram_cell[    1380] = 32'h58f1af69;
    ram_cell[    1381] = 32'h6ae259f4;
    ram_cell[    1382] = 32'h55a73350;
    ram_cell[    1383] = 32'h48c6c93f;
    ram_cell[    1384] = 32'hb1b7f409;
    ram_cell[    1385] = 32'h15d12cb2;
    ram_cell[    1386] = 32'hcc923b35;
    ram_cell[    1387] = 32'h5f8fd90e;
    ram_cell[    1388] = 32'hfb20fcd7;
    ram_cell[    1389] = 32'h9b9b3a61;
    ram_cell[    1390] = 32'hd832dc02;
    ram_cell[    1391] = 32'h05f576bc;
    ram_cell[    1392] = 32'h8f6959ac;
    ram_cell[    1393] = 32'h8597e135;
    ram_cell[    1394] = 32'h7d8f0e28;
    ram_cell[    1395] = 32'h2a71b054;
    ram_cell[    1396] = 32'ha779f9ec;
    ram_cell[    1397] = 32'he784f6f3;
    ram_cell[    1398] = 32'h613a9a27;
    ram_cell[    1399] = 32'h1be61269;
    ram_cell[    1400] = 32'h46399617;
    ram_cell[    1401] = 32'hbb4cd0dd;
    ram_cell[    1402] = 32'h1d3de62f;
    ram_cell[    1403] = 32'h2056e150;
    ram_cell[    1404] = 32'h4e334ae2;
    ram_cell[    1405] = 32'h7c67349b;
    ram_cell[    1406] = 32'h8a1b130e;
    ram_cell[    1407] = 32'hcdca181e;
    ram_cell[    1408] = 32'h6c5cc639;
    ram_cell[    1409] = 32'hf26c8324;
    ram_cell[    1410] = 32'h25c3b451;
    ram_cell[    1411] = 32'h2bd388e0;
    ram_cell[    1412] = 32'hf30f050c;
    ram_cell[    1413] = 32'h95ac5771;
    ram_cell[    1414] = 32'ha5b92cc0;
    ram_cell[    1415] = 32'h3443c51d;
    ram_cell[    1416] = 32'h94fbfe76;
    ram_cell[    1417] = 32'hbc339750;
    ram_cell[    1418] = 32'hf496a0d6;
    ram_cell[    1419] = 32'hacf2c570;
    ram_cell[    1420] = 32'hb4429245;
    ram_cell[    1421] = 32'h8dbb0526;
    ram_cell[    1422] = 32'ha647d40a;
    ram_cell[    1423] = 32'h02dbf9fd;
    ram_cell[    1424] = 32'h1572408f;
    ram_cell[    1425] = 32'hfb3a654d;
    ram_cell[    1426] = 32'hc539e414;
    ram_cell[    1427] = 32'hde6c365c;
    ram_cell[    1428] = 32'hc8fe505b;
    ram_cell[    1429] = 32'h9ebeb4e7;
    ram_cell[    1430] = 32'h3ead5ce9;
    ram_cell[    1431] = 32'h440ff9ed;
    ram_cell[    1432] = 32'ha2a3658b;
    ram_cell[    1433] = 32'hd6a1887f;
    ram_cell[    1434] = 32'h637dedc7;
    ram_cell[    1435] = 32'h0cf991e6;
    ram_cell[    1436] = 32'hb24f5047;
    ram_cell[    1437] = 32'h9ca7df1c;
    ram_cell[    1438] = 32'hb531ef84;
    ram_cell[    1439] = 32'h12c9cd8b;
    ram_cell[    1440] = 32'h1c4b42b9;
    ram_cell[    1441] = 32'hd6fab503;
    ram_cell[    1442] = 32'h4a43c459;
    ram_cell[    1443] = 32'h0953241a;
    ram_cell[    1444] = 32'hb01ed7d9;
    ram_cell[    1445] = 32'h3322abf0;
    ram_cell[    1446] = 32'hae61281e;
    ram_cell[    1447] = 32'h1f606580;
    ram_cell[    1448] = 32'h3b85bb26;
    ram_cell[    1449] = 32'h7638a7b0;
    ram_cell[    1450] = 32'hfc5b731e;
    ram_cell[    1451] = 32'hced5ad45;
    ram_cell[    1452] = 32'h67d84d1a;
    ram_cell[    1453] = 32'h13dbe658;
    ram_cell[    1454] = 32'h467e7049;
    ram_cell[    1455] = 32'h79d18c6a;
    ram_cell[    1456] = 32'h94912ab6;
    ram_cell[    1457] = 32'hc82fbaaf;
    ram_cell[    1458] = 32'h2682aa75;
    ram_cell[    1459] = 32'hf3f8493e;
    ram_cell[    1460] = 32'h22ed7bdd;
    ram_cell[    1461] = 32'h28cbdf1c;
    ram_cell[    1462] = 32'h862ce8c3;
    ram_cell[    1463] = 32'hef972d3d;
    ram_cell[    1464] = 32'hb16b6733;
    ram_cell[    1465] = 32'h0244a519;
    ram_cell[    1466] = 32'h11ec4904;
    ram_cell[    1467] = 32'h0a3486a3;
    ram_cell[    1468] = 32'h941a697f;
    ram_cell[    1469] = 32'h15414846;
    ram_cell[    1470] = 32'hd94fabcc;
    ram_cell[    1471] = 32'h0b985628;
    ram_cell[    1472] = 32'h81912810;
    ram_cell[    1473] = 32'h8be6f42f;
    ram_cell[    1474] = 32'h8cd6e47a;
    ram_cell[    1475] = 32'h8e462c20;
    ram_cell[    1476] = 32'ha8ac5ae7;
    ram_cell[    1477] = 32'he3388262;
    ram_cell[    1478] = 32'hf14f0ce0;
    ram_cell[    1479] = 32'hef9e8800;
    ram_cell[    1480] = 32'hcc9fc31f;
    ram_cell[    1481] = 32'h55ce3969;
    ram_cell[    1482] = 32'h273e5b35;
    ram_cell[    1483] = 32'h46fcea8f;
    ram_cell[    1484] = 32'h6131bd80;
    ram_cell[    1485] = 32'h3d9d8086;
    ram_cell[    1486] = 32'h98d4213f;
    ram_cell[    1487] = 32'h1a43a4a9;
    ram_cell[    1488] = 32'h85435a69;
    ram_cell[    1489] = 32'h50a801ef;
    ram_cell[    1490] = 32'h696076bb;
    ram_cell[    1491] = 32'hcd608111;
    ram_cell[    1492] = 32'h040d7dbf;
    ram_cell[    1493] = 32'he6d5f0df;
    ram_cell[    1494] = 32'h84f4eae6;
    ram_cell[    1495] = 32'h712901c1;
    ram_cell[    1496] = 32'h8e8be67b;
    ram_cell[    1497] = 32'he5e6fcaa;
    ram_cell[    1498] = 32'hb7bc58b4;
    ram_cell[    1499] = 32'h7458deb0;
    ram_cell[    1500] = 32'hb85b6d49;
    ram_cell[    1501] = 32'h2472ced4;
    ram_cell[    1502] = 32'h973c063b;
    ram_cell[    1503] = 32'h8732b1b7;
    ram_cell[    1504] = 32'ha9fb8821;
    ram_cell[    1505] = 32'h2cef5cb0;
    ram_cell[    1506] = 32'he4b53047;
    ram_cell[    1507] = 32'h829440bc;
    ram_cell[    1508] = 32'h0a9b3aa8;
    ram_cell[    1509] = 32'h2177d535;
    ram_cell[    1510] = 32'hf7454f8b;
    ram_cell[    1511] = 32'hd45ba30f;
    ram_cell[    1512] = 32'hbd0deee7;
    ram_cell[    1513] = 32'h6e42bd0c;
    ram_cell[    1514] = 32'h8433706e;
    ram_cell[    1515] = 32'h96ca92e9;
    ram_cell[    1516] = 32'hb172b156;
    ram_cell[    1517] = 32'h90e75162;
    ram_cell[    1518] = 32'h7426e8ea;
    ram_cell[    1519] = 32'h3233be64;
    ram_cell[    1520] = 32'h869fa3cd;
    ram_cell[    1521] = 32'h6c5b9bc4;
    ram_cell[    1522] = 32'h6e701e78;
    ram_cell[    1523] = 32'hdb4d95fb;
    ram_cell[    1524] = 32'h46ffb7bd;
    ram_cell[    1525] = 32'hb613af2a;
    ram_cell[    1526] = 32'h6c6a2a4a;
    ram_cell[    1527] = 32'h9185b278;
    ram_cell[    1528] = 32'h6f84846d;
    ram_cell[    1529] = 32'h7aed5ab0;
    ram_cell[    1530] = 32'hfb061840;
    ram_cell[    1531] = 32'he575fc67;
    ram_cell[    1532] = 32'h3386e7d3;
    ram_cell[    1533] = 32'h0b6e175a;
    ram_cell[    1534] = 32'h2f65f4f2;
    ram_cell[    1535] = 32'ha9c52c03;
    ram_cell[    1536] = 32'h88378741;
    ram_cell[    1537] = 32'h8bd73478;
    ram_cell[    1538] = 32'hc12ed77f;
    ram_cell[    1539] = 32'hd3a35f7e;
    ram_cell[    1540] = 32'hf29bb41e;
    ram_cell[    1541] = 32'h2e3f4024;
    ram_cell[    1542] = 32'h971027e3;
    ram_cell[    1543] = 32'h872d2130;
    ram_cell[    1544] = 32'hff31cf02;
    ram_cell[    1545] = 32'h5bbe2830;
    ram_cell[    1546] = 32'h64056af5;
    ram_cell[    1547] = 32'h41d6e76a;
    ram_cell[    1548] = 32'h7ce4ab65;
    ram_cell[    1549] = 32'hadb7ad58;
    ram_cell[    1550] = 32'he0c52f3c;
    ram_cell[    1551] = 32'h3b0366ca;
    ram_cell[    1552] = 32'h8a6f1336;
    ram_cell[    1553] = 32'h4593e082;
    ram_cell[    1554] = 32'h3a1c11c1;
    ram_cell[    1555] = 32'hc7ad2d77;
    ram_cell[    1556] = 32'h828ddb78;
    ram_cell[    1557] = 32'h134dcb30;
    ram_cell[    1558] = 32'h23927520;
    ram_cell[    1559] = 32'hdea3dcd3;
    ram_cell[    1560] = 32'h3e2a0897;
    ram_cell[    1561] = 32'h1aaed18a;
    ram_cell[    1562] = 32'hc5322cb2;
    ram_cell[    1563] = 32'h79878ad6;
    ram_cell[    1564] = 32'h5ff36545;
    ram_cell[    1565] = 32'h6a8eeed7;
    ram_cell[    1566] = 32'h89edb72e;
    ram_cell[    1567] = 32'h26e054da;
    ram_cell[    1568] = 32'ha7f1ea14;
    ram_cell[    1569] = 32'h151e9750;
    ram_cell[    1570] = 32'h8399bd6e;
    ram_cell[    1571] = 32'hbb990a17;
    ram_cell[    1572] = 32'h6a6a46e0;
    ram_cell[    1573] = 32'hb6391c01;
    ram_cell[    1574] = 32'he9f3a358;
    ram_cell[    1575] = 32'h2bbe53b0;
    ram_cell[    1576] = 32'h47d3c004;
    ram_cell[    1577] = 32'h55154ca0;
    ram_cell[    1578] = 32'h43489220;
    ram_cell[    1579] = 32'hd8ecfcc6;
    ram_cell[    1580] = 32'h36d8c0cc;
    ram_cell[    1581] = 32'h3cb6c8ba;
    ram_cell[    1582] = 32'h20820552;
    ram_cell[    1583] = 32'he3f4b6b3;
    ram_cell[    1584] = 32'hbb459194;
    ram_cell[    1585] = 32'h1fed5385;
    ram_cell[    1586] = 32'hbbaaecb6;
    ram_cell[    1587] = 32'h36cba288;
    ram_cell[    1588] = 32'h540cae23;
    ram_cell[    1589] = 32'h1774dbc9;
    ram_cell[    1590] = 32'hb9288dd6;
    ram_cell[    1591] = 32'hb5349c73;
    ram_cell[    1592] = 32'h251dd750;
    ram_cell[    1593] = 32'h9f827543;
    ram_cell[    1594] = 32'h244f9bc3;
    ram_cell[    1595] = 32'h57d8846c;
    ram_cell[    1596] = 32'hfe016d94;
    ram_cell[    1597] = 32'h85de026b;
    ram_cell[    1598] = 32'h006e1ab9;
    ram_cell[    1599] = 32'h68cc1580;
    ram_cell[    1600] = 32'hc950df8e;
    ram_cell[    1601] = 32'h0e2edb95;
    ram_cell[    1602] = 32'h4e247b18;
    ram_cell[    1603] = 32'h7a9f1868;
    ram_cell[    1604] = 32'h4b68084a;
    ram_cell[    1605] = 32'hb89cbc29;
    ram_cell[    1606] = 32'h07b57dda;
    ram_cell[    1607] = 32'h69516654;
    ram_cell[    1608] = 32'h59055ff3;
    ram_cell[    1609] = 32'ha557c804;
    ram_cell[    1610] = 32'hae379f25;
    ram_cell[    1611] = 32'hb7c2ce82;
    ram_cell[    1612] = 32'hd1103d19;
    ram_cell[    1613] = 32'h18d1f88d;
    ram_cell[    1614] = 32'h0990fcf6;
    ram_cell[    1615] = 32'hff34ca98;
    ram_cell[    1616] = 32'hfaf75caf;
    ram_cell[    1617] = 32'h7ac419f4;
    ram_cell[    1618] = 32'h51e99f75;
    ram_cell[    1619] = 32'ha01d2ce8;
    ram_cell[    1620] = 32'h4ee6784c;
    ram_cell[    1621] = 32'h074134e9;
    ram_cell[    1622] = 32'haa1149d5;
    ram_cell[    1623] = 32'h7f9822ad;
    ram_cell[    1624] = 32'h14f91630;
    ram_cell[    1625] = 32'h34b303ec;
    ram_cell[    1626] = 32'hba9ab250;
    ram_cell[    1627] = 32'he993b2b3;
    ram_cell[    1628] = 32'h157a5881;
    ram_cell[    1629] = 32'h5a342b8e;
    ram_cell[    1630] = 32'h282bbe40;
    ram_cell[    1631] = 32'hf87db4c4;
    ram_cell[    1632] = 32'h4835c23c;
    ram_cell[    1633] = 32'hbb814c86;
    ram_cell[    1634] = 32'h195428fa;
    ram_cell[    1635] = 32'h0c92666a;
    ram_cell[    1636] = 32'h916f5c27;
    ram_cell[    1637] = 32'h43f2892e;
    ram_cell[    1638] = 32'h1c9d610c;
    ram_cell[    1639] = 32'h12ca7eaf;
    ram_cell[    1640] = 32'h6488ecf9;
    ram_cell[    1641] = 32'h77fac7c2;
    ram_cell[    1642] = 32'h62e015fe;
    ram_cell[    1643] = 32'h1c75ed55;
    ram_cell[    1644] = 32'hbbd12ffb;
    ram_cell[    1645] = 32'h61701507;
    ram_cell[    1646] = 32'h39db61a8;
    ram_cell[    1647] = 32'h38df94a1;
    ram_cell[    1648] = 32'h3e0e2049;
    ram_cell[    1649] = 32'h16ce2b9e;
    ram_cell[    1650] = 32'hd4d1d919;
    ram_cell[    1651] = 32'hbfdf4969;
    ram_cell[    1652] = 32'h70de3e4c;
    ram_cell[    1653] = 32'h6f68e690;
    ram_cell[    1654] = 32'h77051229;
    ram_cell[    1655] = 32'hd1037138;
    ram_cell[    1656] = 32'hca20927a;
    ram_cell[    1657] = 32'hfbbda139;
    ram_cell[    1658] = 32'he2424f44;
    ram_cell[    1659] = 32'h4de79fa1;
    ram_cell[    1660] = 32'hb0d85091;
    ram_cell[    1661] = 32'h67839a7d;
    ram_cell[    1662] = 32'h39cdd6e3;
    ram_cell[    1663] = 32'hfd52b0f4;
    ram_cell[    1664] = 32'hf02c2c26;
    ram_cell[    1665] = 32'h1c2a24ba;
    ram_cell[    1666] = 32'hcd117794;
    ram_cell[    1667] = 32'hacc1ac03;
    ram_cell[    1668] = 32'had0c73b8;
    ram_cell[    1669] = 32'hfba4ad13;
    ram_cell[    1670] = 32'h525fcbfe;
    ram_cell[    1671] = 32'h23eacd07;
    ram_cell[    1672] = 32'hd0e7fd1a;
    ram_cell[    1673] = 32'h6a4d49a7;
    ram_cell[    1674] = 32'hc443753f;
    ram_cell[    1675] = 32'h7e2bdfea;
    ram_cell[    1676] = 32'hd694a847;
    ram_cell[    1677] = 32'h0d33d7ca;
    ram_cell[    1678] = 32'h1158fc64;
    ram_cell[    1679] = 32'h68b56778;
    ram_cell[    1680] = 32'h2e67653c;
    ram_cell[    1681] = 32'hc7b5dbcf;
    ram_cell[    1682] = 32'h6f91474b;
    ram_cell[    1683] = 32'hb02f9168;
    ram_cell[    1684] = 32'hc29240aa;
    ram_cell[    1685] = 32'hf3c18db1;
    ram_cell[    1686] = 32'hfba3321c;
    ram_cell[    1687] = 32'h16c18a5e;
    ram_cell[    1688] = 32'hc7caae94;
    ram_cell[    1689] = 32'hb0c5cf71;
    ram_cell[    1690] = 32'heba0e970;
    ram_cell[    1691] = 32'h020be33b;
    ram_cell[    1692] = 32'h2c480a1c;
    ram_cell[    1693] = 32'h57eefee6;
    ram_cell[    1694] = 32'h95340474;
    ram_cell[    1695] = 32'hc7a9a4d7;
    ram_cell[    1696] = 32'h7a779dcf;
    ram_cell[    1697] = 32'h37add476;
    ram_cell[    1698] = 32'hd2f6b288;
    ram_cell[    1699] = 32'h15f09e95;
    ram_cell[    1700] = 32'hd359f637;
    ram_cell[    1701] = 32'h785cad6f;
    ram_cell[    1702] = 32'h7ffa2da0;
    ram_cell[    1703] = 32'h5b4b33c0;
    ram_cell[    1704] = 32'h59aba5e0;
    ram_cell[    1705] = 32'h10bcc6d1;
    ram_cell[    1706] = 32'h5deaabe5;
    ram_cell[    1707] = 32'he488ec53;
    ram_cell[    1708] = 32'h6a00dfc7;
    ram_cell[    1709] = 32'hb1d3d4b3;
    ram_cell[    1710] = 32'heff92f45;
    ram_cell[    1711] = 32'h2d814729;
    ram_cell[    1712] = 32'h143445b3;
    ram_cell[    1713] = 32'hf98315e7;
    ram_cell[    1714] = 32'h1868707b;
    ram_cell[    1715] = 32'h809a5a85;
    ram_cell[    1716] = 32'h171e32b2;
    ram_cell[    1717] = 32'h774f01b5;
    ram_cell[    1718] = 32'h4f641b8d;
    ram_cell[    1719] = 32'hb274a330;
    ram_cell[    1720] = 32'h77fd5449;
    ram_cell[    1721] = 32'h83a165b3;
    ram_cell[    1722] = 32'h42c99858;
    ram_cell[    1723] = 32'h9da0bb3c;
    ram_cell[    1724] = 32'h35c97652;
    ram_cell[    1725] = 32'h2cd8e3be;
    ram_cell[    1726] = 32'h4160d7cb;
    ram_cell[    1727] = 32'hf7340d44;
    ram_cell[    1728] = 32'h320a4c9c;
    ram_cell[    1729] = 32'h0fd1e24c;
    ram_cell[    1730] = 32'h26ae1226;
    ram_cell[    1731] = 32'hc7b828b8;
    ram_cell[    1732] = 32'h16eeb5bb;
    ram_cell[    1733] = 32'h91fe1107;
    ram_cell[    1734] = 32'hf91991ac;
    ram_cell[    1735] = 32'he4b29e91;
    ram_cell[    1736] = 32'hbb02e0c9;
    ram_cell[    1737] = 32'ha029ecc6;
    ram_cell[    1738] = 32'h3a60c4c0;
    ram_cell[    1739] = 32'h2cfe668c;
    ram_cell[    1740] = 32'h35978d27;
    ram_cell[    1741] = 32'hfe88ff53;
    ram_cell[    1742] = 32'hf057bd4b;
    ram_cell[    1743] = 32'h1178772e;
    ram_cell[    1744] = 32'he48fe743;
    ram_cell[    1745] = 32'h40d10b9b;
    ram_cell[    1746] = 32'h4c336547;
    ram_cell[    1747] = 32'h68638a2d;
    ram_cell[    1748] = 32'hbb303ed9;
    ram_cell[    1749] = 32'h7d8e6ae3;
    ram_cell[    1750] = 32'h364383a4;
    ram_cell[    1751] = 32'hf3a22358;
    ram_cell[    1752] = 32'h14c8a4f1;
    ram_cell[    1753] = 32'hd7dec5b4;
    ram_cell[    1754] = 32'h8522fe53;
    ram_cell[    1755] = 32'hd1e8a187;
    ram_cell[    1756] = 32'hb8c0e78e;
    ram_cell[    1757] = 32'ha5fb35e1;
    ram_cell[    1758] = 32'h00bb1e60;
    ram_cell[    1759] = 32'h89250767;
    ram_cell[    1760] = 32'hce554e0a;
    ram_cell[    1761] = 32'h4f87b4ad;
    ram_cell[    1762] = 32'h531af8a8;
    ram_cell[    1763] = 32'hef1d4235;
    ram_cell[    1764] = 32'h9c59ada1;
    ram_cell[    1765] = 32'hc5562238;
    ram_cell[    1766] = 32'hbd543cf2;
    ram_cell[    1767] = 32'hebce2984;
    ram_cell[    1768] = 32'h222c924c;
    ram_cell[    1769] = 32'h5f0179dc;
    ram_cell[    1770] = 32'he43f6ef1;
    ram_cell[    1771] = 32'h6b9689de;
    ram_cell[    1772] = 32'hbc8162bc;
    ram_cell[    1773] = 32'h2ba81299;
    ram_cell[    1774] = 32'h8f0a15fd;
    ram_cell[    1775] = 32'h668de4f5;
    ram_cell[    1776] = 32'h6237e97b;
    ram_cell[    1777] = 32'h114950a1;
    ram_cell[    1778] = 32'hfebe6aef;
    ram_cell[    1779] = 32'h78cfcdb2;
    ram_cell[    1780] = 32'h3a8d443c;
    ram_cell[    1781] = 32'h678ca9b9;
    ram_cell[    1782] = 32'h961ebe19;
    ram_cell[    1783] = 32'hc7887b5d;
    ram_cell[    1784] = 32'h82f9d4e3;
    ram_cell[    1785] = 32'h808a9f01;
    ram_cell[    1786] = 32'h32202179;
    ram_cell[    1787] = 32'h7b611261;
    ram_cell[    1788] = 32'h83896d89;
    ram_cell[    1789] = 32'hb868cfe4;
    ram_cell[    1790] = 32'h8c555a8a;
    ram_cell[    1791] = 32'hfef3070a;
    ram_cell[    1792] = 32'h89e6f77f;
    ram_cell[    1793] = 32'h55d09131;
    ram_cell[    1794] = 32'h8eb92c1c;
    ram_cell[    1795] = 32'h18032e67;
    ram_cell[    1796] = 32'h1d8922b3;
    ram_cell[    1797] = 32'h8f696f9d;
    ram_cell[    1798] = 32'h2ed19f7c;
    ram_cell[    1799] = 32'h3683273e;
    ram_cell[    1800] = 32'h6b4b0868;
    ram_cell[    1801] = 32'h14871e66;
    ram_cell[    1802] = 32'h50ec3b06;
    ram_cell[    1803] = 32'h02786e88;
    ram_cell[    1804] = 32'h8831fb8e;
    ram_cell[    1805] = 32'hd9fbda0e;
    ram_cell[    1806] = 32'h2fc4ca11;
    ram_cell[    1807] = 32'h2e2ce60d;
    ram_cell[    1808] = 32'h4cfa60f9;
    ram_cell[    1809] = 32'h8891a1e9;
    ram_cell[    1810] = 32'h84d96d93;
    ram_cell[    1811] = 32'had3d2341;
    ram_cell[    1812] = 32'hd8e32218;
    ram_cell[    1813] = 32'h871f4592;
    ram_cell[    1814] = 32'h0d0dce21;
    ram_cell[    1815] = 32'h524c6c69;
    ram_cell[    1816] = 32'h2eab2aa2;
    ram_cell[    1817] = 32'h6ea9af04;
    ram_cell[    1818] = 32'h0acea33b;
    ram_cell[    1819] = 32'he87b67d4;
    ram_cell[    1820] = 32'h1630581e;
    ram_cell[    1821] = 32'h39529e60;
    ram_cell[    1822] = 32'h413ea388;
    ram_cell[    1823] = 32'h3432af9a;
    ram_cell[    1824] = 32'h95fb4c77;
    ram_cell[    1825] = 32'h0402bf19;
    ram_cell[    1826] = 32'h914fba78;
    ram_cell[    1827] = 32'h890e818c;
    ram_cell[    1828] = 32'h8b52971a;
    ram_cell[    1829] = 32'h73e1bc18;
    ram_cell[    1830] = 32'h209d39de;
    ram_cell[    1831] = 32'h4e754546;
    ram_cell[    1832] = 32'h44d46129;
    ram_cell[    1833] = 32'h046087f4;
    ram_cell[    1834] = 32'hcf77e353;
    ram_cell[    1835] = 32'hfb1bbbcf;
    ram_cell[    1836] = 32'hdac48450;
    ram_cell[    1837] = 32'hf60946fe;
    ram_cell[    1838] = 32'hd37cc34a;
    ram_cell[    1839] = 32'hdd63b0e1;
    ram_cell[    1840] = 32'hca00082a;
    ram_cell[    1841] = 32'h0fb291ff;
    ram_cell[    1842] = 32'hda066ab6;
    ram_cell[    1843] = 32'h855fdc6f;
    ram_cell[    1844] = 32'h69bd5349;
    ram_cell[    1845] = 32'h04164ebd;
    ram_cell[    1846] = 32'h00943f77;
    ram_cell[    1847] = 32'h7c689887;
    ram_cell[    1848] = 32'h608790a7;
    ram_cell[    1849] = 32'hb4045fbb;
    ram_cell[    1850] = 32'h5a243267;
    ram_cell[    1851] = 32'hfbb8efe5;
    ram_cell[    1852] = 32'h30c5b3ca;
    ram_cell[    1853] = 32'hb2b27a1f;
    ram_cell[    1854] = 32'hd5449118;
    ram_cell[    1855] = 32'hb9b40203;
    ram_cell[    1856] = 32'h92845351;
    ram_cell[    1857] = 32'he023161a;
    ram_cell[    1858] = 32'h4584a169;
    ram_cell[    1859] = 32'h90ae426c;
    ram_cell[    1860] = 32'he96269c7;
    ram_cell[    1861] = 32'he1aa25c2;
    ram_cell[    1862] = 32'h8024adbc;
    ram_cell[    1863] = 32'h9ce86518;
    ram_cell[    1864] = 32'h331bfef2;
    ram_cell[    1865] = 32'h6b329ffc;
    ram_cell[    1866] = 32'h39c7133e;
    ram_cell[    1867] = 32'h62c63481;
    ram_cell[    1868] = 32'h64137ab6;
    ram_cell[    1869] = 32'hd90f5c2d;
    ram_cell[    1870] = 32'hc12a7b09;
    ram_cell[    1871] = 32'h130aecfc;
    ram_cell[    1872] = 32'h7e1bf162;
    ram_cell[    1873] = 32'hf0924e92;
    ram_cell[    1874] = 32'hf78448ca;
    ram_cell[    1875] = 32'hd370b82b;
    ram_cell[    1876] = 32'hb5249f8e;
    ram_cell[    1877] = 32'h6440d045;
    ram_cell[    1878] = 32'h7302fe35;
    ram_cell[    1879] = 32'h8cb2f4ff;
    ram_cell[    1880] = 32'hc900aa86;
    ram_cell[    1881] = 32'hac001769;
    ram_cell[    1882] = 32'h10ed187f;
    ram_cell[    1883] = 32'h889b5b53;
    ram_cell[    1884] = 32'he97627eb;
    ram_cell[    1885] = 32'he9fee1e2;
    ram_cell[    1886] = 32'h84c25a97;
    ram_cell[    1887] = 32'hecac618f;
    ram_cell[    1888] = 32'h69927744;
    ram_cell[    1889] = 32'hf82a5b38;
    ram_cell[    1890] = 32'hdec56e75;
    ram_cell[    1891] = 32'hbbf439f6;
    ram_cell[    1892] = 32'h6db5bf93;
    ram_cell[    1893] = 32'h959e83fd;
    ram_cell[    1894] = 32'h7f2ed3dd;
    ram_cell[    1895] = 32'h51cacb4c;
    ram_cell[    1896] = 32'h1fc2debe;
    ram_cell[    1897] = 32'h098a9f3b;
    ram_cell[    1898] = 32'h1231d8be;
    ram_cell[    1899] = 32'h36d250f6;
    ram_cell[    1900] = 32'h4b47110d;
    ram_cell[    1901] = 32'h63771a93;
    ram_cell[    1902] = 32'ha5b796e9;
    ram_cell[    1903] = 32'hd5dd5be1;
    ram_cell[    1904] = 32'h37fa1ba9;
    ram_cell[    1905] = 32'h5a5dff97;
    ram_cell[    1906] = 32'h676debe4;
    ram_cell[    1907] = 32'hfa16839f;
    ram_cell[    1908] = 32'h00302a89;
    ram_cell[    1909] = 32'h18d71b0d;
    ram_cell[    1910] = 32'h5d33b58f;
    ram_cell[    1911] = 32'h253b299f;
    ram_cell[    1912] = 32'h6c398666;
    ram_cell[    1913] = 32'h5ea3de01;
    ram_cell[    1914] = 32'hca409629;
    ram_cell[    1915] = 32'h97529825;
    ram_cell[    1916] = 32'h255a38da;
    ram_cell[    1917] = 32'h46d65de9;
    ram_cell[    1918] = 32'h03cab196;
    ram_cell[    1919] = 32'h1c398266;
    ram_cell[    1920] = 32'h54a6028b;
    ram_cell[    1921] = 32'h49d2055c;
    ram_cell[    1922] = 32'hc2264e5f;
    ram_cell[    1923] = 32'hfc4aa1cc;
    ram_cell[    1924] = 32'h6d117587;
    ram_cell[    1925] = 32'h65afe10a;
    ram_cell[    1926] = 32'hc19aab39;
    ram_cell[    1927] = 32'h4013a320;
    ram_cell[    1928] = 32'h3c9e14d5;
    ram_cell[    1929] = 32'h5d2ea40c;
    ram_cell[    1930] = 32'h980d8eb2;
    ram_cell[    1931] = 32'he8b84410;
    ram_cell[    1932] = 32'he99aaab6;
    ram_cell[    1933] = 32'h03d9c637;
    ram_cell[    1934] = 32'hc3eefd37;
    ram_cell[    1935] = 32'h11572dc4;
    ram_cell[    1936] = 32'h7e34ff4b;
    ram_cell[    1937] = 32'hc6aa4f45;
    ram_cell[    1938] = 32'hfae50b16;
    ram_cell[    1939] = 32'he5cdd72c;
    ram_cell[    1940] = 32'h222aade6;
    ram_cell[    1941] = 32'h01337294;
    ram_cell[    1942] = 32'h3e38aa83;
    ram_cell[    1943] = 32'hd3414a3c;
    ram_cell[    1944] = 32'h134d0af7;
    ram_cell[    1945] = 32'hc77bbfe3;
    ram_cell[    1946] = 32'he4297c11;
    ram_cell[    1947] = 32'h96139b57;
    ram_cell[    1948] = 32'habcf2b43;
    ram_cell[    1949] = 32'hc46525fc;
    ram_cell[    1950] = 32'hb7f8b90f;
    ram_cell[    1951] = 32'hf4e53e9d;
    ram_cell[    1952] = 32'h6a18f05b;
    ram_cell[    1953] = 32'h2a3cd79c;
    ram_cell[    1954] = 32'hf00570e8;
    ram_cell[    1955] = 32'h34d5d98e;
    ram_cell[    1956] = 32'hcf5dd808;
    ram_cell[    1957] = 32'h409ef09c;
    ram_cell[    1958] = 32'h42ed76b4;
    ram_cell[    1959] = 32'h54e368c0;
    ram_cell[    1960] = 32'hb5dd3119;
    ram_cell[    1961] = 32'h1b156fdc;
    ram_cell[    1962] = 32'he2b70d1a;
    ram_cell[    1963] = 32'h251d67c3;
    ram_cell[    1964] = 32'ha3f5e273;
    ram_cell[    1965] = 32'h80194626;
    ram_cell[    1966] = 32'h900dab60;
    ram_cell[    1967] = 32'hf193384e;
    ram_cell[    1968] = 32'h717c53cc;
    ram_cell[    1969] = 32'hf4259415;
    ram_cell[    1970] = 32'h13e2863c;
    ram_cell[    1971] = 32'h18398769;
    ram_cell[    1972] = 32'h9c8c17df;
    ram_cell[    1973] = 32'h324195aa;
    ram_cell[    1974] = 32'h4d104f5e;
    ram_cell[    1975] = 32'h86152d62;
    ram_cell[    1976] = 32'hefc0b7e0;
    ram_cell[    1977] = 32'hdcb4ecf2;
    ram_cell[    1978] = 32'ha97aab23;
    ram_cell[    1979] = 32'ha174ccae;
    ram_cell[    1980] = 32'hfdcfe7ad;
    ram_cell[    1981] = 32'h134e1564;
    ram_cell[    1982] = 32'h5128807b;
    ram_cell[    1983] = 32'h4cebcb0b;
    ram_cell[    1984] = 32'hf470dd59;
    ram_cell[    1985] = 32'hf459aa3e;
    ram_cell[    1986] = 32'h4e49ab34;
    ram_cell[    1987] = 32'h12c89a4c;
    ram_cell[    1988] = 32'h8ebd9c01;
    ram_cell[    1989] = 32'hf29cb187;
    ram_cell[    1990] = 32'hc227a70f;
    ram_cell[    1991] = 32'h3187623b;
    ram_cell[    1992] = 32'ha9ffb306;
    ram_cell[    1993] = 32'h2407f159;
    ram_cell[    1994] = 32'heed8f2b0;
    ram_cell[    1995] = 32'hd75c28de;
    ram_cell[    1996] = 32'hfa288cfc;
    ram_cell[    1997] = 32'he1a827b3;
    ram_cell[    1998] = 32'h0a183391;
    ram_cell[    1999] = 32'hdf45e9ec;
    ram_cell[    2000] = 32'hef037396;
    ram_cell[    2001] = 32'hfebef5e8;
    ram_cell[    2002] = 32'h45d23f07;
    ram_cell[    2003] = 32'h439a253c;
    ram_cell[    2004] = 32'h45e8ebb0;
    ram_cell[    2005] = 32'ha5e1e1c5;
    ram_cell[    2006] = 32'h0ca9cfa8;
    ram_cell[    2007] = 32'h1b99333f;
    ram_cell[    2008] = 32'hd35fc38e;
    ram_cell[    2009] = 32'ha6938464;
    ram_cell[    2010] = 32'h28c388e5;
    ram_cell[    2011] = 32'h03f1bae3;
    ram_cell[    2012] = 32'h47ad78f6;
    ram_cell[    2013] = 32'hcac32c90;
    ram_cell[    2014] = 32'hd0ff0c8c;
    ram_cell[    2015] = 32'h5e7cfdb4;
    ram_cell[    2016] = 32'he05bd074;
    ram_cell[    2017] = 32'hb71d03cc;
    ram_cell[    2018] = 32'hdc02271c;
    ram_cell[    2019] = 32'h134983d8;
    ram_cell[    2020] = 32'hb82138bd;
    ram_cell[    2021] = 32'h6cecf187;
    ram_cell[    2022] = 32'hacf4abbc;
    ram_cell[    2023] = 32'hd46b56c3;
    ram_cell[    2024] = 32'he5972381;
    ram_cell[    2025] = 32'h92a7e264;
    ram_cell[    2026] = 32'h65351453;
    ram_cell[    2027] = 32'hd04ee3a6;
    ram_cell[    2028] = 32'h6d026dae;
    ram_cell[    2029] = 32'h4aebee82;
    ram_cell[    2030] = 32'hb1477ed8;
    ram_cell[    2031] = 32'h5cc65573;
    ram_cell[    2032] = 32'h50d2cb5b;
    ram_cell[    2033] = 32'h7592d4a8;
    ram_cell[    2034] = 32'h17d6d0fb;
    ram_cell[    2035] = 32'h268d3756;
    ram_cell[    2036] = 32'h56a89024;
    ram_cell[    2037] = 32'h0de4018c;
    ram_cell[    2038] = 32'h2ea4e24f;
    ram_cell[    2039] = 32'hd766311f;
    ram_cell[    2040] = 32'hb1daa1a4;
    ram_cell[    2041] = 32'h168b9d43;
    ram_cell[    2042] = 32'h20704f69;
    ram_cell[    2043] = 32'hf22295ed;
    ram_cell[    2044] = 32'ha8cbbac6;
    ram_cell[    2045] = 32'h8deafc74;
    ram_cell[    2046] = 32'h37862fd0;
    ram_cell[    2047] = 32'h4b795190;
    // src matrix B
    ram_cell[    2048] = 32'h3e607f2c;
    ram_cell[    2049] = 32'h441f3fdb;
    ram_cell[    2050] = 32'hd4e79616;
    ram_cell[    2051] = 32'hfae49ce8;
    ram_cell[    2052] = 32'hc8ecc566;
    ram_cell[    2053] = 32'h5e2dbd52;
    ram_cell[    2054] = 32'h889e461a;
    ram_cell[    2055] = 32'h188379ed;
    ram_cell[    2056] = 32'hc85f0e38;
    ram_cell[    2057] = 32'hf31643ab;
    ram_cell[    2058] = 32'hde0ccf28;
    ram_cell[    2059] = 32'hcdd3c9ce;
    ram_cell[    2060] = 32'h0238c2dd;
    ram_cell[    2061] = 32'hb27a4807;
    ram_cell[    2062] = 32'h618f6cf5;
    ram_cell[    2063] = 32'h7308dad9;
    ram_cell[    2064] = 32'hd51b0b96;
    ram_cell[    2065] = 32'h83a8c218;
    ram_cell[    2066] = 32'hdda7a003;
    ram_cell[    2067] = 32'hc3680e59;
    ram_cell[    2068] = 32'h565c580b;
    ram_cell[    2069] = 32'he5741856;
    ram_cell[    2070] = 32'h5d3f4665;
    ram_cell[    2071] = 32'h8240d900;
    ram_cell[    2072] = 32'hb172c5c2;
    ram_cell[    2073] = 32'hb19ec839;
    ram_cell[    2074] = 32'h7a254e79;
    ram_cell[    2075] = 32'h7884274d;
    ram_cell[    2076] = 32'h51eeec53;
    ram_cell[    2077] = 32'h84c8314a;
    ram_cell[    2078] = 32'h4db05973;
    ram_cell[    2079] = 32'h65c09b98;
    ram_cell[    2080] = 32'h4f51e69a;
    ram_cell[    2081] = 32'h3ac3935f;
    ram_cell[    2082] = 32'h9ed9f701;
    ram_cell[    2083] = 32'h3f4f951c;
    ram_cell[    2084] = 32'hdd2e47f2;
    ram_cell[    2085] = 32'hb5619c5a;
    ram_cell[    2086] = 32'h26cd56a2;
    ram_cell[    2087] = 32'h1ceeadda;
    ram_cell[    2088] = 32'h9a19f8ae;
    ram_cell[    2089] = 32'hc95e18c2;
    ram_cell[    2090] = 32'h004c5b8a;
    ram_cell[    2091] = 32'h1a631e97;
    ram_cell[    2092] = 32'he2e572ec;
    ram_cell[    2093] = 32'he4680132;
    ram_cell[    2094] = 32'h7610817e;
    ram_cell[    2095] = 32'h61629652;
    ram_cell[    2096] = 32'h63038208;
    ram_cell[    2097] = 32'h617fc5c0;
    ram_cell[    2098] = 32'hc32aa43a;
    ram_cell[    2099] = 32'h1de267af;
    ram_cell[    2100] = 32'he818eb4f;
    ram_cell[    2101] = 32'h2e9404ca;
    ram_cell[    2102] = 32'h1bc674ef;
    ram_cell[    2103] = 32'hc67cbe54;
    ram_cell[    2104] = 32'h7e3453c5;
    ram_cell[    2105] = 32'hc0060d4e;
    ram_cell[    2106] = 32'h19ed3ae6;
    ram_cell[    2107] = 32'heb6298f3;
    ram_cell[    2108] = 32'h8cd40381;
    ram_cell[    2109] = 32'ha02af960;
    ram_cell[    2110] = 32'hc51b6869;
    ram_cell[    2111] = 32'h420967a0;
    ram_cell[    2112] = 32'h3a5327d3;
    ram_cell[    2113] = 32'h895b8b75;
    ram_cell[    2114] = 32'hb3060625;
    ram_cell[    2115] = 32'h2fcd8b25;
    ram_cell[    2116] = 32'he8ffd594;
    ram_cell[    2117] = 32'he7eb1f99;
    ram_cell[    2118] = 32'hf3725c34;
    ram_cell[    2119] = 32'h12c397c9;
    ram_cell[    2120] = 32'h49c4480c;
    ram_cell[    2121] = 32'h5ca67b29;
    ram_cell[    2122] = 32'h27db9ed6;
    ram_cell[    2123] = 32'hb5f19466;
    ram_cell[    2124] = 32'h9b98f282;
    ram_cell[    2125] = 32'h49233913;
    ram_cell[    2126] = 32'hee968b9d;
    ram_cell[    2127] = 32'h768d9f75;
    ram_cell[    2128] = 32'hdf083609;
    ram_cell[    2129] = 32'h9cabe629;
    ram_cell[    2130] = 32'head7d48f;
    ram_cell[    2131] = 32'hb6911ecc;
    ram_cell[    2132] = 32'h5e02266f;
    ram_cell[    2133] = 32'h62ce36c8;
    ram_cell[    2134] = 32'h0efbeeb6;
    ram_cell[    2135] = 32'h13589c01;
    ram_cell[    2136] = 32'h3eb338d6;
    ram_cell[    2137] = 32'hc644285e;
    ram_cell[    2138] = 32'h483c5b56;
    ram_cell[    2139] = 32'h124c6c6c;
    ram_cell[    2140] = 32'hde8b96f4;
    ram_cell[    2141] = 32'h78cdb88a;
    ram_cell[    2142] = 32'hb763cbf1;
    ram_cell[    2143] = 32'h573b8022;
    ram_cell[    2144] = 32'h04fe7740;
    ram_cell[    2145] = 32'h90e10eb5;
    ram_cell[    2146] = 32'h603d7e54;
    ram_cell[    2147] = 32'he0b16eb6;
    ram_cell[    2148] = 32'hb62ec517;
    ram_cell[    2149] = 32'hdc46de7e;
    ram_cell[    2150] = 32'h028519c7;
    ram_cell[    2151] = 32'hf1055af6;
    ram_cell[    2152] = 32'ha88ea4dc;
    ram_cell[    2153] = 32'h13ed4467;
    ram_cell[    2154] = 32'h4e296100;
    ram_cell[    2155] = 32'h865b213c;
    ram_cell[    2156] = 32'h46bacf30;
    ram_cell[    2157] = 32'h3eca9cdf;
    ram_cell[    2158] = 32'h82890883;
    ram_cell[    2159] = 32'hb2ee1b8c;
    ram_cell[    2160] = 32'ha12efea1;
    ram_cell[    2161] = 32'ha81351d6;
    ram_cell[    2162] = 32'hc3d3495c;
    ram_cell[    2163] = 32'h65fce1e6;
    ram_cell[    2164] = 32'hbc98de28;
    ram_cell[    2165] = 32'he46c9863;
    ram_cell[    2166] = 32'ha72d50f4;
    ram_cell[    2167] = 32'h74c5e167;
    ram_cell[    2168] = 32'h9c11d423;
    ram_cell[    2169] = 32'h61bb23ce;
    ram_cell[    2170] = 32'h1e136de3;
    ram_cell[    2171] = 32'h8e0ef3f6;
    ram_cell[    2172] = 32'hbfac6853;
    ram_cell[    2173] = 32'habcfa564;
    ram_cell[    2174] = 32'hdfa9a02f;
    ram_cell[    2175] = 32'hb0cde1a4;
    ram_cell[    2176] = 32'h870b044d;
    ram_cell[    2177] = 32'h33510212;
    ram_cell[    2178] = 32'h094ad04b;
    ram_cell[    2179] = 32'h456aeef6;
    ram_cell[    2180] = 32'hf1d75804;
    ram_cell[    2181] = 32'h1664300b;
    ram_cell[    2182] = 32'hd7221ff5;
    ram_cell[    2183] = 32'h1c007412;
    ram_cell[    2184] = 32'h40eab029;
    ram_cell[    2185] = 32'h53ca38cf;
    ram_cell[    2186] = 32'h7d6ca16c;
    ram_cell[    2187] = 32'h11bc0d95;
    ram_cell[    2188] = 32'h81bb52b0;
    ram_cell[    2189] = 32'h06a4c9a4;
    ram_cell[    2190] = 32'h3cd716a8;
    ram_cell[    2191] = 32'hebc22ac2;
    ram_cell[    2192] = 32'h45733e53;
    ram_cell[    2193] = 32'hdfbf44e1;
    ram_cell[    2194] = 32'he57c2ca5;
    ram_cell[    2195] = 32'h3c616ce1;
    ram_cell[    2196] = 32'hfa05a4de;
    ram_cell[    2197] = 32'hd191c72b;
    ram_cell[    2198] = 32'h288b920a;
    ram_cell[    2199] = 32'h1dbfdfb7;
    ram_cell[    2200] = 32'h27bc25ad;
    ram_cell[    2201] = 32'h53e52180;
    ram_cell[    2202] = 32'h4f35cb72;
    ram_cell[    2203] = 32'hef8d411c;
    ram_cell[    2204] = 32'h3c0addf0;
    ram_cell[    2205] = 32'h11f561fa;
    ram_cell[    2206] = 32'hd5a466ba;
    ram_cell[    2207] = 32'hd44bcc61;
    ram_cell[    2208] = 32'h6834b490;
    ram_cell[    2209] = 32'h24fa9d42;
    ram_cell[    2210] = 32'h545faf41;
    ram_cell[    2211] = 32'ha423e81d;
    ram_cell[    2212] = 32'h6b7a23f5;
    ram_cell[    2213] = 32'h2230a2bd;
    ram_cell[    2214] = 32'hcf3e800b;
    ram_cell[    2215] = 32'h3b34b3e9;
    ram_cell[    2216] = 32'hf377568f;
    ram_cell[    2217] = 32'h6f4fa03e;
    ram_cell[    2218] = 32'h342b6427;
    ram_cell[    2219] = 32'h30a6b0f3;
    ram_cell[    2220] = 32'hd231456f;
    ram_cell[    2221] = 32'hca51fa54;
    ram_cell[    2222] = 32'h7a47301d;
    ram_cell[    2223] = 32'h90ae2ba8;
    ram_cell[    2224] = 32'he92fc243;
    ram_cell[    2225] = 32'h8051cbae;
    ram_cell[    2226] = 32'h3d441d90;
    ram_cell[    2227] = 32'h539be8b1;
    ram_cell[    2228] = 32'h56274482;
    ram_cell[    2229] = 32'hccb77cd0;
    ram_cell[    2230] = 32'h3bedf4be;
    ram_cell[    2231] = 32'hbd7fd58d;
    ram_cell[    2232] = 32'hf530a0fa;
    ram_cell[    2233] = 32'hd1f21170;
    ram_cell[    2234] = 32'h5eb961ab;
    ram_cell[    2235] = 32'hcf22b5d0;
    ram_cell[    2236] = 32'h030496c7;
    ram_cell[    2237] = 32'h061acdb5;
    ram_cell[    2238] = 32'h389bcc92;
    ram_cell[    2239] = 32'h816b6f8d;
    ram_cell[    2240] = 32'h2f18e6be;
    ram_cell[    2241] = 32'h17f79a9c;
    ram_cell[    2242] = 32'hdc89a934;
    ram_cell[    2243] = 32'h19f022c8;
    ram_cell[    2244] = 32'hf0914ab4;
    ram_cell[    2245] = 32'h63f839c7;
    ram_cell[    2246] = 32'hd4d7fadd;
    ram_cell[    2247] = 32'hb0989f17;
    ram_cell[    2248] = 32'h9e14a69f;
    ram_cell[    2249] = 32'h1f49707f;
    ram_cell[    2250] = 32'h1e9ecb4d;
    ram_cell[    2251] = 32'hea2bf5ed;
    ram_cell[    2252] = 32'hae12cfab;
    ram_cell[    2253] = 32'h94040195;
    ram_cell[    2254] = 32'h8b5d1e8f;
    ram_cell[    2255] = 32'he59ce105;
    ram_cell[    2256] = 32'h5a23b510;
    ram_cell[    2257] = 32'hbc77d43f;
    ram_cell[    2258] = 32'hf4adf04b;
    ram_cell[    2259] = 32'h2f06bc0e;
    ram_cell[    2260] = 32'had782d2d;
    ram_cell[    2261] = 32'h8e47f1e4;
    ram_cell[    2262] = 32'hda7bb9d3;
    ram_cell[    2263] = 32'h1524597f;
    ram_cell[    2264] = 32'h2c72828b;
    ram_cell[    2265] = 32'he9fb5d72;
    ram_cell[    2266] = 32'h081a4e74;
    ram_cell[    2267] = 32'h90b181cd;
    ram_cell[    2268] = 32'hbcd9e051;
    ram_cell[    2269] = 32'h37fcf2c5;
    ram_cell[    2270] = 32'he2fa3c59;
    ram_cell[    2271] = 32'he2294f25;
    ram_cell[    2272] = 32'hf4f0369f;
    ram_cell[    2273] = 32'hbf46ffa6;
    ram_cell[    2274] = 32'ha991977e;
    ram_cell[    2275] = 32'h25917491;
    ram_cell[    2276] = 32'h3a225109;
    ram_cell[    2277] = 32'h9bd062b3;
    ram_cell[    2278] = 32'hf2eb84e1;
    ram_cell[    2279] = 32'h81b1bf5b;
    ram_cell[    2280] = 32'h562d1bec;
    ram_cell[    2281] = 32'h30fa79ca;
    ram_cell[    2282] = 32'hb1ef9bdc;
    ram_cell[    2283] = 32'hd499cc46;
    ram_cell[    2284] = 32'hb0cef92a;
    ram_cell[    2285] = 32'h6124fb4d;
    ram_cell[    2286] = 32'h72501c45;
    ram_cell[    2287] = 32'h21ea2a4d;
    ram_cell[    2288] = 32'h8d424f40;
    ram_cell[    2289] = 32'h8e9ba4c9;
    ram_cell[    2290] = 32'h39f5f795;
    ram_cell[    2291] = 32'hb4931a43;
    ram_cell[    2292] = 32'h1d7d2811;
    ram_cell[    2293] = 32'h97bf2a8c;
    ram_cell[    2294] = 32'h747e12d9;
    ram_cell[    2295] = 32'hadd6f426;
    ram_cell[    2296] = 32'h4427baec;
    ram_cell[    2297] = 32'hc1ee0298;
    ram_cell[    2298] = 32'h2c8d3244;
    ram_cell[    2299] = 32'h4d5465eb;
    ram_cell[    2300] = 32'h19d70bb4;
    ram_cell[    2301] = 32'hd0b2f87c;
    ram_cell[    2302] = 32'h3b51ff7c;
    ram_cell[    2303] = 32'h4d5a4f29;
    ram_cell[    2304] = 32'hf01eeb1b;
    ram_cell[    2305] = 32'h8b88f2cf;
    ram_cell[    2306] = 32'h209be0ca;
    ram_cell[    2307] = 32'h063d0eed;
    ram_cell[    2308] = 32'h5038dca8;
    ram_cell[    2309] = 32'hc3c7d79a;
    ram_cell[    2310] = 32'ha5eacf4b;
    ram_cell[    2311] = 32'hb2873be6;
    ram_cell[    2312] = 32'ha24bec1e;
    ram_cell[    2313] = 32'hcd4d1e9b;
    ram_cell[    2314] = 32'h3b73fdde;
    ram_cell[    2315] = 32'h91d2e299;
    ram_cell[    2316] = 32'h1e533977;
    ram_cell[    2317] = 32'h2fa50385;
    ram_cell[    2318] = 32'hede57b82;
    ram_cell[    2319] = 32'hc1cd9404;
    ram_cell[    2320] = 32'h07ca397d;
    ram_cell[    2321] = 32'h13897bc1;
    ram_cell[    2322] = 32'he22b3ca2;
    ram_cell[    2323] = 32'h2d944f0b;
    ram_cell[    2324] = 32'h181f5e7e;
    ram_cell[    2325] = 32'h6a3fe013;
    ram_cell[    2326] = 32'h035b414d;
    ram_cell[    2327] = 32'h4ab511c8;
    ram_cell[    2328] = 32'h3527ad77;
    ram_cell[    2329] = 32'h906b4499;
    ram_cell[    2330] = 32'he8354728;
    ram_cell[    2331] = 32'h403d87f9;
    ram_cell[    2332] = 32'h54f78539;
    ram_cell[    2333] = 32'h4ea55ffd;
    ram_cell[    2334] = 32'h5ba7ef1b;
    ram_cell[    2335] = 32'h8e425102;
    ram_cell[    2336] = 32'ha481c717;
    ram_cell[    2337] = 32'h087e0dd2;
    ram_cell[    2338] = 32'hb1a82e17;
    ram_cell[    2339] = 32'h6afbee3a;
    ram_cell[    2340] = 32'hffcb0690;
    ram_cell[    2341] = 32'hf86f2938;
    ram_cell[    2342] = 32'hf498c490;
    ram_cell[    2343] = 32'h08d143c7;
    ram_cell[    2344] = 32'hdd973b79;
    ram_cell[    2345] = 32'h7905d29a;
    ram_cell[    2346] = 32'h449ad6ad;
    ram_cell[    2347] = 32'hc9f455a7;
    ram_cell[    2348] = 32'h1e8b2dbe;
    ram_cell[    2349] = 32'h3595f647;
    ram_cell[    2350] = 32'ha90b2d6c;
    ram_cell[    2351] = 32'h6b994875;
    ram_cell[    2352] = 32'he0eac077;
    ram_cell[    2353] = 32'he16199b8;
    ram_cell[    2354] = 32'h66ca4d9a;
    ram_cell[    2355] = 32'hb204eb89;
    ram_cell[    2356] = 32'h92dece5c;
    ram_cell[    2357] = 32'h3d7ad9ec;
    ram_cell[    2358] = 32'h3556866c;
    ram_cell[    2359] = 32'h95c72022;
    ram_cell[    2360] = 32'hb5cec863;
    ram_cell[    2361] = 32'h6a384cac;
    ram_cell[    2362] = 32'h9708bd55;
    ram_cell[    2363] = 32'h0a5e2ce0;
    ram_cell[    2364] = 32'h4d70f7ef;
    ram_cell[    2365] = 32'h3b14ad13;
    ram_cell[    2366] = 32'h0c11b305;
    ram_cell[    2367] = 32'h1f5b66ea;
    ram_cell[    2368] = 32'h9854aebe;
    ram_cell[    2369] = 32'h92023e0a;
    ram_cell[    2370] = 32'h22cce97d;
    ram_cell[    2371] = 32'h186ba720;
    ram_cell[    2372] = 32'h8d189448;
    ram_cell[    2373] = 32'h8bc4a146;
    ram_cell[    2374] = 32'haff5b9c5;
    ram_cell[    2375] = 32'hed4ab101;
    ram_cell[    2376] = 32'hfbe22fbf;
    ram_cell[    2377] = 32'h2fc97639;
    ram_cell[    2378] = 32'h89b14755;
    ram_cell[    2379] = 32'h28a58705;
    ram_cell[    2380] = 32'h56c55720;
    ram_cell[    2381] = 32'h171399c1;
    ram_cell[    2382] = 32'h88bad59e;
    ram_cell[    2383] = 32'h7a039e34;
    ram_cell[    2384] = 32'h273893d4;
    ram_cell[    2385] = 32'h9f4d7694;
    ram_cell[    2386] = 32'h9b70d5e1;
    ram_cell[    2387] = 32'he36a6478;
    ram_cell[    2388] = 32'hff2ac936;
    ram_cell[    2389] = 32'h8e023fda;
    ram_cell[    2390] = 32'h1a656143;
    ram_cell[    2391] = 32'h81140fee;
    ram_cell[    2392] = 32'h550aa7b5;
    ram_cell[    2393] = 32'h2d540e51;
    ram_cell[    2394] = 32'h95088d88;
    ram_cell[    2395] = 32'hed60e7f4;
    ram_cell[    2396] = 32'hed13fe6c;
    ram_cell[    2397] = 32'ha611e744;
    ram_cell[    2398] = 32'h8278cd23;
    ram_cell[    2399] = 32'hfda784f6;
    ram_cell[    2400] = 32'h6dfa32e7;
    ram_cell[    2401] = 32'hc1896dbc;
    ram_cell[    2402] = 32'h2612775e;
    ram_cell[    2403] = 32'h9ed57b37;
    ram_cell[    2404] = 32'hd17db52f;
    ram_cell[    2405] = 32'h04c75615;
    ram_cell[    2406] = 32'h1c4c936a;
    ram_cell[    2407] = 32'hfed22c69;
    ram_cell[    2408] = 32'hb7f47d37;
    ram_cell[    2409] = 32'ha71c376f;
    ram_cell[    2410] = 32'h3053b095;
    ram_cell[    2411] = 32'hc7844ff3;
    ram_cell[    2412] = 32'h8fc33e85;
    ram_cell[    2413] = 32'h8689c86b;
    ram_cell[    2414] = 32'h7eac5e33;
    ram_cell[    2415] = 32'h5665c7c9;
    ram_cell[    2416] = 32'h99ad433a;
    ram_cell[    2417] = 32'h0465f549;
    ram_cell[    2418] = 32'hc6d81778;
    ram_cell[    2419] = 32'ha11e8139;
    ram_cell[    2420] = 32'h8a303a5a;
    ram_cell[    2421] = 32'hf435027d;
    ram_cell[    2422] = 32'h5a84d418;
    ram_cell[    2423] = 32'h3be40eb3;
    ram_cell[    2424] = 32'hbcf8046a;
    ram_cell[    2425] = 32'h8f10cfc8;
    ram_cell[    2426] = 32'h8d9ec474;
    ram_cell[    2427] = 32'h54156a7d;
    ram_cell[    2428] = 32'h71e50047;
    ram_cell[    2429] = 32'he1be0094;
    ram_cell[    2430] = 32'h2cf8fd99;
    ram_cell[    2431] = 32'h8c54342c;
    ram_cell[    2432] = 32'h743c022e;
    ram_cell[    2433] = 32'h64be50ea;
    ram_cell[    2434] = 32'h365ffb5a;
    ram_cell[    2435] = 32'h815d7be4;
    ram_cell[    2436] = 32'h10727613;
    ram_cell[    2437] = 32'h471edd16;
    ram_cell[    2438] = 32'hfa12f29d;
    ram_cell[    2439] = 32'h6233b2c7;
    ram_cell[    2440] = 32'h92c9514f;
    ram_cell[    2441] = 32'ha619b2ab;
    ram_cell[    2442] = 32'h52314155;
    ram_cell[    2443] = 32'h3779cd08;
    ram_cell[    2444] = 32'h71fb8a17;
    ram_cell[    2445] = 32'hefcdbb7a;
    ram_cell[    2446] = 32'h9dc64f83;
    ram_cell[    2447] = 32'h96a30126;
    ram_cell[    2448] = 32'h999cbd13;
    ram_cell[    2449] = 32'h0b0fb46c;
    ram_cell[    2450] = 32'hd827fd37;
    ram_cell[    2451] = 32'hc898632c;
    ram_cell[    2452] = 32'h6923a5e6;
    ram_cell[    2453] = 32'hfa9f1130;
    ram_cell[    2454] = 32'h9138fb51;
    ram_cell[    2455] = 32'h7ba7053a;
    ram_cell[    2456] = 32'hdb0a9bc6;
    ram_cell[    2457] = 32'h1624b575;
    ram_cell[    2458] = 32'h6e7c0aa8;
    ram_cell[    2459] = 32'h0818899d;
    ram_cell[    2460] = 32'hf81db3d0;
    ram_cell[    2461] = 32'h4863c54a;
    ram_cell[    2462] = 32'h0ef7bd9b;
    ram_cell[    2463] = 32'h9dba889d;
    ram_cell[    2464] = 32'h077f9cf5;
    ram_cell[    2465] = 32'h98438732;
    ram_cell[    2466] = 32'h8a645b49;
    ram_cell[    2467] = 32'h961a6448;
    ram_cell[    2468] = 32'h5165f280;
    ram_cell[    2469] = 32'hfbee8c02;
    ram_cell[    2470] = 32'h2c9e0718;
    ram_cell[    2471] = 32'h8bc7b404;
    ram_cell[    2472] = 32'he6b4b12a;
    ram_cell[    2473] = 32'h1e14879b;
    ram_cell[    2474] = 32'h2b08962e;
    ram_cell[    2475] = 32'h6e16c289;
    ram_cell[    2476] = 32'h7f99c7c0;
    ram_cell[    2477] = 32'hd489520a;
    ram_cell[    2478] = 32'he89ca85f;
    ram_cell[    2479] = 32'hc98312fc;
    ram_cell[    2480] = 32'h895da33f;
    ram_cell[    2481] = 32'h4954493e;
    ram_cell[    2482] = 32'h6fb54b44;
    ram_cell[    2483] = 32'h337ac9bd;
    ram_cell[    2484] = 32'hd9f787ac;
    ram_cell[    2485] = 32'h8e9de5d8;
    ram_cell[    2486] = 32'hcbef6f0e;
    ram_cell[    2487] = 32'ha734e298;
    ram_cell[    2488] = 32'hb7498699;
    ram_cell[    2489] = 32'h9a995036;
    ram_cell[    2490] = 32'h15c71cc7;
    ram_cell[    2491] = 32'h011ab683;
    ram_cell[    2492] = 32'h73067526;
    ram_cell[    2493] = 32'haa8cf341;
    ram_cell[    2494] = 32'h951ee053;
    ram_cell[    2495] = 32'ha78f9756;
    ram_cell[    2496] = 32'h53f3a132;
    ram_cell[    2497] = 32'h65c5a58b;
    ram_cell[    2498] = 32'h730fb56e;
    ram_cell[    2499] = 32'h56ac50a1;
    ram_cell[    2500] = 32'hc8d48cca;
    ram_cell[    2501] = 32'h48d91995;
    ram_cell[    2502] = 32'h60d9df8b;
    ram_cell[    2503] = 32'h58ec73f7;
    ram_cell[    2504] = 32'h9da18701;
    ram_cell[    2505] = 32'hd04b709f;
    ram_cell[    2506] = 32'hd93f857d;
    ram_cell[    2507] = 32'hbe070ef8;
    ram_cell[    2508] = 32'h3958c661;
    ram_cell[    2509] = 32'ha7109939;
    ram_cell[    2510] = 32'h4b7c89f6;
    ram_cell[    2511] = 32'h195d517a;
    ram_cell[    2512] = 32'h8ec7f0ce;
    ram_cell[    2513] = 32'h70baec5a;
    ram_cell[    2514] = 32'h98216ce5;
    ram_cell[    2515] = 32'h720e046c;
    ram_cell[    2516] = 32'hf121a64a;
    ram_cell[    2517] = 32'hb26f2676;
    ram_cell[    2518] = 32'h9ceae1e2;
    ram_cell[    2519] = 32'ha800c8f1;
    ram_cell[    2520] = 32'he3c25484;
    ram_cell[    2521] = 32'hc7511d71;
    ram_cell[    2522] = 32'h4947c6fd;
    ram_cell[    2523] = 32'h68547571;
    ram_cell[    2524] = 32'hfb4a6b55;
    ram_cell[    2525] = 32'he3050d2c;
    ram_cell[    2526] = 32'h110f7f1a;
    ram_cell[    2527] = 32'h46a2864c;
    ram_cell[    2528] = 32'hef25a847;
    ram_cell[    2529] = 32'h580bcc83;
    ram_cell[    2530] = 32'hd4e7855d;
    ram_cell[    2531] = 32'h26fd6af4;
    ram_cell[    2532] = 32'h5af86487;
    ram_cell[    2533] = 32'h35472d94;
    ram_cell[    2534] = 32'h5e98d3c3;
    ram_cell[    2535] = 32'h18f152e8;
    ram_cell[    2536] = 32'h265cacbc;
    ram_cell[    2537] = 32'h4bd1d0d5;
    ram_cell[    2538] = 32'h00ccb4f8;
    ram_cell[    2539] = 32'hef0b8d45;
    ram_cell[    2540] = 32'ha8b1e031;
    ram_cell[    2541] = 32'hafb089ef;
    ram_cell[    2542] = 32'hceb3223d;
    ram_cell[    2543] = 32'hf3f9f74d;
    ram_cell[    2544] = 32'h4a3ed0f9;
    ram_cell[    2545] = 32'h290e32d6;
    ram_cell[    2546] = 32'h571d099d;
    ram_cell[    2547] = 32'hb1ccc113;
    ram_cell[    2548] = 32'h8017e1d4;
    ram_cell[    2549] = 32'hc1cf89ff;
    ram_cell[    2550] = 32'hbeffea81;
    ram_cell[    2551] = 32'h353cf7f2;
    ram_cell[    2552] = 32'hb51a8131;
    ram_cell[    2553] = 32'h7c899527;
    ram_cell[    2554] = 32'haadce387;
    ram_cell[    2555] = 32'h97ac46a3;
    ram_cell[    2556] = 32'h32f501b3;
    ram_cell[    2557] = 32'hc789a9fd;
    ram_cell[    2558] = 32'hc2d40995;
    ram_cell[    2559] = 32'h0bd4eac7;
    ram_cell[    2560] = 32'hba998a3d;
    ram_cell[    2561] = 32'hd4657cbd;
    ram_cell[    2562] = 32'h2747ee5b;
    ram_cell[    2563] = 32'h003969f5;
    ram_cell[    2564] = 32'h93eaa496;
    ram_cell[    2565] = 32'h3304304e;
    ram_cell[    2566] = 32'h8369651c;
    ram_cell[    2567] = 32'hd18e3259;
    ram_cell[    2568] = 32'h47f32dac;
    ram_cell[    2569] = 32'h205a0cbd;
    ram_cell[    2570] = 32'h58313d87;
    ram_cell[    2571] = 32'h7ef27e65;
    ram_cell[    2572] = 32'h48ab4abc;
    ram_cell[    2573] = 32'h71d05253;
    ram_cell[    2574] = 32'h1cad349a;
    ram_cell[    2575] = 32'h36a67370;
    ram_cell[    2576] = 32'hb3b7c236;
    ram_cell[    2577] = 32'h478ba010;
    ram_cell[    2578] = 32'hc7b463a8;
    ram_cell[    2579] = 32'hd8d39662;
    ram_cell[    2580] = 32'hb34f1d60;
    ram_cell[    2581] = 32'h47299a72;
    ram_cell[    2582] = 32'h57e6ffe2;
    ram_cell[    2583] = 32'h77caca48;
    ram_cell[    2584] = 32'h97a2e7e7;
    ram_cell[    2585] = 32'hcc496da8;
    ram_cell[    2586] = 32'hbde6ac88;
    ram_cell[    2587] = 32'h7ec793bd;
    ram_cell[    2588] = 32'h39088df4;
    ram_cell[    2589] = 32'h9a72f664;
    ram_cell[    2590] = 32'h4f6b3bcb;
    ram_cell[    2591] = 32'h45a8d260;
    ram_cell[    2592] = 32'hddf54171;
    ram_cell[    2593] = 32'hcbf55d46;
    ram_cell[    2594] = 32'h7c78d7e3;
    ram_cell[    2595] = 32'ha47cb47d;
    ram_cell[    2596] = 32'ha9849d94;
    ram_cell[    2597] = 32'h1a40f690;
    ram_cell[    2598] = 32'h37157c69;
    ram_cell[    2599] = 32'h0c94f27d;
    ram_cell[    2600] = 32'hdff31f7c;
    ram_cell[    2601] = 32'h964939a8;
    ram_cell[    2602] = 32'hbad53f48;
    ram_cell[    2603] = 32'h9b097d82;
    ram_cell[    2604] = 32'h039a5b6a;
    ram_cell[    2605] = 32'hd5b45432;
    ram_cell[    2606] = 32'h0958f1ba;
    ram_cell[    2607] = 32'ha9eb0eec;
    ram_cell[    2608] = 32'h7c16296e;
    ram_cell[    2609] = 32'h9744cff5;
    ram_cell[    2610] = 32'h34a93bce;
    ram_cell[    2611] = 32'hb8efabf4;
    ram_cell[    2612] = 32'hc4b29234;
    ram_cell[    2613] = 32'h559a2ab7;
    ram_cell[    2614] = 32'h6ddd1e90;
    ram_cell[    2615] = 32'hf7c6d009;
    ram_cell[    2616] = 32'h8c1915a6;
    ram_cell[    2617] = 32'h0b8e2236;
    ram_cell[    2618] = 32'h6be2c265;
    ram_cell[    2619] = 32'h7ed28480;
    ram_cell[    2620] = 32'he0b54d00;
    ram_cell[    2621] = 32'h7bccbba1;
    ram_cell[    2622] = 32'h4bc68b64;
    ram_cell[    2623] = 32'h7af46e02;
    ram_cell[    2624] = 32'hf16151b5;
    ram_cell[    2625] = 32'hbe335b1a;
    ram_cell[    2626] = 32'h344e2bcf;
    ram_cell[    2627] = 32'h311ccd02;
    ram_cell[    2628] = 32'h37b9817f;
    ram_cell[    2629] = 32'hc27d5d5d;
    ram_cell[    2630] = 32'hfd9b4001;
    ram_cell[    2631] = 32'h578fd045;
    ram_cell[    2632] = 32'h3996b363;
    ram_cell[    2633] = 32'h9567cc90;
    ram_cell[    2634] = 32'h2c06f27c;
    ram_cell[    2635] = 32'hf4f321e6;
    ram_cell[    2636] = 32'h15598208;
    ram_cell[    2637] = 32'ha9b46454;
    ram_cell[    2638] = 32'h6dd21d8d;
    ram_cell[    2639] = 32'had790f07;
    ram_cell[    2640] = 32'h51a86bbf;
    ram_cell[    2641] = 32'h97c07844;
    ram_cell[    2642] = 32'h3903e263;
    ram_cell[    2643] = 32'ha1b178d7;
    ram_cell[    2644] = 32'h9c3ba1b0;
    ram_cell[    2645] = 32'h601cbd32;
    ram_cell[    2646] = 32'hd9f790e3;
    ram_cell[    2647] = 32'h60f7e5dc;
    ram_cell[    2648] = 32'h0cdb3e1a;
    ram_cell[    2649] = 32'h20668d9d;
    ram_cell[    2650] = 32'hf275f1a2;
    ram_cell[    2651] = 32'h7f6ddf5a;
    ram_cell[    2652] = 32'h5d37d650;
    ram_cell[    2653] = 32'hafa9a821;
    ram_cell[    2654] = 32'hedb93da5;
    ram_cell[    2655] = 32'h47cecbd3;
    ram_cell[    2656] = 32'h86e106b3;
    ram_cell[    2657] = 32'h800edad5;
    ram_cell[    2658] = 32'hb15e9a0f;
    ram_cell[    2659] = 32'h5a760c49;
    ram_cell[    2660] = 32'h99d470f2;
    ram_cell[    2661] = 32'h9bf944dc;
    ram_cell[    2662] = 32'hda21b0df;
    ram_cell[    2663] = 32'h8dea0879;
    ram_cell[    2664] = 32'hb948ea0c;
    ram_cell[    2665] = 32'hfd6c32c1;
    ram_cell[    2666] = 32'hfe899eb6;
    ram_cell[    2667] = 32'h50a3204e;
    ram_cell[    2668] = 32'h552e21f3;
    ram_cell[    2669] = 32'h215315f9;
    ram_cell[    2670] = 32'hf23ad3f3;
    ram_cell[    2671] = 32'h4cd326f1;
    ram_cell[    2672] = 32'ha37833d7;
    ram_cell[    2673] = 32'h92dabc0c;
    ram_cell[    2674] = 32'h266a6daa;
    ram_cell[    2675] = 32'h61a85933;
    ram_cell[    2676] = 32'hcfc2b539;
    ram_cell[    2677] = 32'hfc090adb;
    ram_cell[    2678] = 32'h59add5cf;
    ram_cell[    2679] = 32'h1f81b3a1;
    ram_cell[    2680] = 32'hd2ccb4f1;
    ram_cell[    2681] = 32'hcadb4758;
    ram_cell[    2682] = 32'hb82377b3;
    ram_cell[    2683] = 32'he60ff2ff;
    ram_cell[    2684] = 32'h2a8eefec;
    ram_cell[    2685] = 32'h8beefde4;
    ram_cell[    2686] = 32'h0e44b0f4;
    ram_cell[    2687] = 32'h495710b3;
    ram_cell[    2688] = 32'h2d30869d;
    ram_cell[    2689] = 32'hfdb0eae5;
    ram_cell[    2690] = 32'hd1f455f3;
    ram_cell[    2691] = 32'h81e45e98;
    ram_cell[    2692] = 32'h65673929;
    ram_cell[    2693] = 32'hd1d58588;
    ram_cell[    2694] = 32'h62b0b60f;
    ram_cell[    2695] = 32'hff29cb89;
    ram_cell[    2696] = 32'h27c65c5d;
    ram_cell[    2697] = 32'hdc1d627e;
    ram_cell[    2698] = 32'h63d65b43;
    ram_cell[    2699] = 32'h041089e8;
    ram_cell[    2700] = 32'h353e69e6;
    ram_cell[    2701] = 32'h20a8cd1c;
    ram_cell[    2702] = 32'hd73db99f;
    ram_cell[    2703] = 32'hb74e2aa9;
    ram_cell[    2704] = 32'h8753a756;
    ram_cell[    2705] = 32'hdf6449a2;
    ram_cell[    2706] = 32'h54955c0b;
    ram_cell[    2707] = 32'hc6ca4e3e;
    ram_cell[    2708] = 32'h370e3740;
    ram_cell[    2709] = 32'h8fa62b74;
    ram_cell[    2710] = 32'h7353061d;
    ram_cell[    2711] = 32'h2c16299d;
    ram_cell[    2712] = 32'h7b7e7a0e;
    ram_cell[    2713] = 32'h446cdd3d;
    ram_cell[    2714] = 32'h3bc0d7af;
    ram_cell[    2715] = 32'h0eb759f7;
    ram_cell[    2716] = 32'h24066c2c;
    ram_cell[    2717] = 32'h99b609e6;
    ram_cell[    2718] = 32'hd0cd5980;
    ram_cell[    2719] = 32'h34898f68;
    ram_cell[    2720] = 32'h0aab158c;
    ram_cell[    2721] = 32'h4e1d2b48;
    ram_cell[    2722] = 32'h6ec2283c;
    ram_cell[    2723] = 32'h53d07d86;
    ram_cell[    2724] = 32'h9547f034;
    ram_cell[    2725] = 32'h68082c84;
    ram_cell[    2726] = 32'hd8093e40;
    ram_cell[    2727] = 32'h947a6826;
    ram_cell[    2728] = 32'h78c015ed;
    ram_cell[    2729] = 32'h2e22fce4;
    ram_cell[    2730] = 32'h5dda5d09;
    ram_cell[    2731] = 32'h80ac313a;
    ram_cell[    2732] = 32'h3e66d6c3;
    ram_cell[    2733] = 32'h06d746ba;
    ram_cell[    2734] = 32'h4742952a;
    ram_cell[    2735] = 32'h089f6e7f;
    ram_cell[    2736] = 32'he1ff2c41;
    ram_cell[    2737] = 32'h2da12519;
    ram_cell[    2738] = 32'h77438a21;
    ram_cell[    2739] = 32'h1ed3b96a;
    ram_cell[    2740] = 32'h8151bb5b;
    ram_cell[    2741] = 32'he260886d;
    ram_cell[    2742] = 32'h0294ab65;
    ram_cell[    2743] = 32'h1266cf69;
    ram_cell[    2744] = 32'h1c1c434b;
    ram_cell[    2745] = 32'h6d2662c4;
    ram_cell[    2746] = 32'hcddec0bb;
    ram_cell[    2747] = 32'hedd584c6;
    ram_cell[    2748] = 32'h1ab77ba0;
    ram_cell[    2749] = 32'hfc773aa0;
    ram_cell[    2750] = 32'hc31efd1b;
    ram_cell[    2751] = 32'h3be1ac24;
    ram_cell[    2752] = 32'h248684da;
    ram_cell[    2753] = 32'h86bcffef;
    ram_cell[    2754] = 32'h239e3fcb;
    ram_cell[    2755] = 32'h77edf314;
    ram_cell[    2756] = 32'h72e97dc9;
    ram_cell[    2757] = 32'h715bc15f;
    ram_cell[    2758] = 32'h90fdc0b5;
    ram_cell[    2759] = 32'h3ad1840b;
    ram_cell[    2760] = 32'hb7c76f1d;
    ram_cell[    2761] = 32'h405cad15;
    ram_cell[    2762] = 32'h9020f9a7;
    ram_cell[    2763] = 32'had4e58e6;
    ram_cell[    2764] = 32'hb7a143b1;
    ram_cell[    2765] = 32'h6d79f432;
    ram_cell[    2766] = 32'hf9a4011b;
    ram_cell[    2767] = 32'h71a36074;
    ram_cell[    2768] = 32'h5638128b;
    ram_cell[    2769] = 32'h7724e7ce;
    ram_cell[    2770] = 32'h993ea7ab;
    ram_cell[    2771] = 32'h40d11f8f;
    ram_cell[    2772] = 32'h86329f97;
    ram_cell[    2773] = 32'h963318de;
    ram_cell[    2774] = 32'h3cc2e992;
    ram_cell[    2775] = 32'h269c1ea9;
    ram_cell[    2776] = 32'h1236ce7c;
    ram_cell[    2777] = 32'h9fd1efa2;
    ram_cell[    2778] = 32'h0f26f09f;
    ram_cell[    2779] = 32'hba4dffac;
    ram_cell[    2780] = 32'h4c09ce61;
    ram_cell[    2781] = 32'h5db4f009;
    ram_cell[    2782] = 32'h4a416789;
    ram_cell[    2783] = 32'h4b6af9f8;
    ram_cell[    2784] = 32'hbd6f4ce9;
    ram_cell[    2785] = 32'h7bf985d0;
    ram_cell[    2786] = 32'hea638fa1;
    ram_cell[    2787] = 32'hd694e376;
    ram_cell[    2788] = 32'h057f31c2;
    ram_cell[    2789] = 32'h055b6405;
    ram_cell[    2790] = 32'hdeabe3fe;
    ram_cell[    2791] = 32'h9e5ce6ed;
    ram_cell[    2792] = 32'hd6348cfc;
    ram_cell[    2793] = 32'he7353b7d;
    ram_cell[    2794] = 32'h777286ff;
    ram_cell[    2795] = 32'hc1077a37;
    ram_cell[    2796] = 32'hc401d69f;
    ram_cell[    2797] = 32'h6b1da257;
    ram_cell[    2798] = 32'h26f1683d;
    ram_cell[    2799] = 32'h58e9bd9a;
    ram_cell[    2800] = 32'h7e8fda4d;
    ram_cell[    2801] = 32'h8d3495a8;
    ram_cell[    2802] = 32'hb1e71968;
    ram_cell[    2803] = 32'h744e05e0;
    ram_cell[    2804] = 32'hb4de29ea;
    ram_cell[    2805] = 32'hd0fdb392;
    ram_cell[    2806] = 32'h73bcf000;
    ram_cell[    2807] = 32'hf8f6c943;
    ram_cell[    2808] = 32'ha88f29b9;
    ram_cell[    2809] = 32'h6a7919e6;
    ram_cell[    2810] = 32'hfdf91aad;
    ram_cell[    2811] = 32'hbbc283a0;
    ram_cell[    2812] = 32'hbf5d326d;
    ram_cell[    2813] = 32'h58c8972f;
    ram_cell[    2814] = 32'hf1d0aac0;
    ram_cell[    2815] = 32'h92c7f9bc;
    ram_cell[    2816] = 32'ha7159462;
    ram_cell[    2817] = 32'h49596c62;
    ram_cell[    2818] = 32'hc28ecf81;
    ram_cell[    2819] = 32'h95d9915b;
    ram_cell[    2820] = 32'h896d765c;
    ram_cell[    2821] = 32'h0d0c88d3;
    ram_cell[    2822] = 32'h5ee99526;
    ram_cell[    2823] = 32'he70db012;
    ram_cell[    2824] = 32'ha2b45306;
    ram_cell[    2825] = 32'h70b08fd0;
    ram_cell[    2826] = 32'hf42de233;
    ram_cell[    2827] = 32'h57dbaeb0;
    ram_cell[    2828] = 32'h9e157dfa;
    ram_cell[    2829] = 32'h813ddb0f;
    ram_cell[    2830] = 32'hc176d454;
    ram_cell[    2831] = 32'h3bf9c29b;
    ram_cell[    2832] = 32'h2b210fac;
    ram_cell[    2833] = 32'h1ee2585a;
    ram_cell[    2834] = 32'ha374626f;
    ram_cell[    2835] = 32'h53e8dd37;
    ram_cell[    2836] = 32'h5a5dbe63;
    ram_cell[    2837] = 32'h0d5bb844;
    ram_cell[    2838] = 32'h7beb5917;
    ram_cell[    2839] = 32'h92820803;
    ram_cell[    2840] = 32'h5cc350e8;
    ram_cell[    2841] = 32'h9b0380c3;
    ram_cell[    2842] = 32'hb593e38a;
    ram_cell[    2843] = 32'h140c1605;
    ram_cell[    2844] = 32'hab38e624;
    ram_cell[    2845] = 32'ha1936878;
    ram_cell[    2846] = 32'hec19ee56;
    ram_cell[    2847] = 32'h8682a085;
    ram_cell[    2848] = 32'he67e81b4;
    ram_cell[    2849] = 32'h2c5259b9;
    ram_cell[    2850] = 32'h882b8ca6;
    ram_cell[    2851] = 32'hfe407e15;
    ram_cell[    2852] = 32'h6106182e;
    ram_cell[    2853] = 32'h7a806cdc;
    ram_cell[    2854] = 32'h7529dde0;
    ram_cell[    2855] = 32'h72c6d45b;
    ram_cell[    2856] = 32'h774adf28;
    ram_cell[    2857] = 32'hf79c4c1d;
    ram_cell[    2858] = 32'hfa2046e0;
    ram_cell[    2859] = 32'h5edf2a95;
    ram_cell[    2860] = 32'h9a1e6c26;
    ram_cell[    2861] = 32'hc9ea0a18;
    ram_cell[    2862] = 32'h19b62c6a;
    ram_cell[    2863] = 32'h5a465628;
    ram_cell[    2864] = 32'h3b790c65;
    ram_cell[    2865] = 32'h9274fd28;
    ram_cell[    2866] = 32'hbcb99933;
    ram_cell[    2867] = 32'hb3bd7c20;
    ram_cell[    2868] = 32'he5e3b365;
    ram_cell[    2869] = 32'h7715a117;
    ram_cell[    2870] = 32'h05954de6;
    ram_cell[    2871] = 32'hff9cf64c;
    ram_cell[    2872] = 32'ha71696f3;
    ram_cell[    2873] = 32'h987e2249;
    ram_cell[    2874] = 32'hdbd06896;
    ram_cell[    2875] = 32'h510bab7c;
    ram_cell[    2876] = 32'hbdace668;
    ram_cell[    2877] = 32'h3fb7ccff;
    ram_cell[    2878] = 32'hd7cfad9b;
    ram_cell[    2879] = 32'h33a48f91;
    ram_cell[    2880] = 32'hd162dc9c;
    ram_cell[    2881] = 32'h9988bfa8;
    ram_cell[    2882] = 32'hed294a61;
    ram_cell[    2883] = 32'hed0cd32f;
    ram_cell[    2884] = 32'hc6f0b852;
    ram_cell[    2885] = 32'h58f76ca8;
    ram_cell[    2886] = 32'h84cc7347;
    ram_cell[    2887] = 32'hc997c439;
    ram_cell[    2888] = 32'h9675d023;
    ram_cell[    2889] = 32'hce3c1897;
    ram_cell[    2890] = 32'ha6e0677c;
    ram_cell[    2891] = 32'h171cc19b;
    ram_cell[    2892] = 32'h18dd5b5c;
    ram_cell[    2893] = 32'heb06e91c;
    ram_cell[    2894] = 32'h2823eb03;
    ram_cell[    2895] = 32'h0e7e3e3b;
    ram_cell[    2896] = 32'h8fe652d2;
    ram_cell[    2897] = 32'hdf9633f1;
    ram_cell[    2898] = 32'hc634bfb2;
    ram_cell[    2899] = 32'h5be98573;
    ram_cell[    2900] = 32'h8ca195fa;
    ram_cell[    2901] = 32'h1fef8e36;
    ram_cell[    2902] = 32'h799f54ee;
    ram_cell[    2903] = 32'hbd54e21f;
    ram_cell[    2904] = 32'hee3e64c6;
    ram_cell[    2905] = 32'h89a84782;
    ram_cell[    2906] = 32'h6fcd1eec;
    ram_cell[    2907] = 32'head276e7;
    ram_cell[    2908] = 32'h2a49d098;
    ram_cell[    2909] = 32'h102cbe36;
    ram_cell[    2910] = 32'hdddff63f;
    ram_cell[    2911] = 32'h7214da83;
    ram_cell[    2912] = 32'h5e244648;
    ram_cell[    2913] = 32'h8ddfbb50;
    ram_cell[    2914] = 32'h796586c0;
    ram_cell[    2915] = 32'h21c62c81;
    ram_cell[    2916] = 32'he0411784;
    ram_cell[    2917] = 32'h763ec029;
    ram_cell[    2918] = 32'h54fbfbe0;
    ram_cell[    2919] = 32'h7a94ef37;
    ram_cell[    2920] = 32'h4d146428;
    ram_cell[    2921] = 32'h4153c7b7;
    ram_cell[    2922] = 32'hf98273f3;
    ram_cell[    2923] = 32'h25ee056c;
    ram_cell[    2924] = 32'hd41d63d2;
    ram_cell[    2925] = 32'h174c81f3;
    ram_cell[    2926] = 32'h89d28201;
    ram_cell[    2927] = 32'he88385ba;
    ram_cell[    2928] = 32'h740303c5;
    ram_cell[    2929] = 32'hf3c07b7b;
    ram_cell[    2930] = 32'hc8c34cd3;
    ram_cell[    2931] = 32'he6d1a1bc;
    ram_cell[    2932] = 32'ha129aaa4;
    ram_cell[    2933] = 32'h40b7eef0;
    ram_cell[    2934] = 32'hfd8a6c53;
    ram_cell[    2935] = 32'h03529701;
    ram_cell[    2936] = 32'h983644f2;
    ram_cell[    2937] = 32'h889e34d5;
    ram_cell[    2938] = 32'hbf2da934;
    ram_cell[    2939] = 32'h52e56811;
    ram_cell[    2940] = 32'hcde1ba4d;
    ram_cell[    2941] = 32'h1c957e0a;
    ram_cell[    2942] = 32'h5ce0415d;
    ram_cell[    2943] = 32'h552d9ba3;
    ram_cell[    2944] = 32'he49a87a8;
    ram_cell[    2945] = 32'hec7329c3;
    ram_cell[    2946] = 32'h4de9aead;
    ram_cell[    2947] = 32'hf12f33e4;
    ram_cell[    2948] = 32'hbc081cb2;
    ram_cell[    2949] = 32'h608dda6a;
    ram_cell[    2950] = 32'h310df8ca;
    ram_cell[    2951] = 32'h5d035347;
    ram_cell[    2952] = 32'h62e9dabf;
    ram_cell[    2953] = 32'h35e62988;
    ram_cell[    2954] = 32'h4bf29923;
    ram_cell[    2955] = 32'ha736f693;
    ram_cell[    2956] = 32'hdb3ee158;
    ram_cell[    2957] = 32'hcb8641e5;
    ram_cell[    2958] = 32'h47454d67;
    ram_cell[    2959] = 32'hc007fd76;
    ram_cell[    2960] = 32'h701602fb;
    ram_cell[    2961] = 32'h85d9b4a5;
    ram_cell[    2962] = 32'h29c5c2d7;
    ram_cell[    2963] = 32'hdc56ff00;
    ram_cell[    2964] = 32'h73a9dfb2;
    ram_cell[    2965] = 32'hd44b8129;
    ram_cell[    2966] = 32'h863cca4f;
    ram_cell[    2967] = 32'h64c601fa;
    ram_cell[    2968] = 32'h4149f8fe;
    ram_cell[    2969] = 32'hbaaf063e;
    ram_cell[    2970] = 32'h6545f059;
    ram_cell[    2971] = 32'ha37fb93c;
    ram_cell[    2972] = 32'hda137508;
    ram_cell[    2973] = 32'h389f2195;
    ram_cell[    2974] = 32'h2385544f;
    ram_cell[    2975] = 32'h85b8d30a;
    ram_cell[    2976] = 32'h78129776;
    ram_cell[    2977] = 32'ha37d5254;
    ram_cell[    2978] = 32'hc4a0738c;
    ram_cell[    2979] = 32'h1d0d637c;
    ram_cell[    2980] = 32'hfab378fc;
    ram_cell[    2981] = 32'he7084563;
    ram_cell[    2982] = 32'hc8ec9ead;
    ram_cell[    2983] = 32'h4c2e9a46;
    ram_cell[    2984] = 32'h65a7fd4c;
    ram_cell[    2985] = 32'hcedbf0f6;
    ram_cell[    2986] = 32'h504aa0dd;
    ram_cell[    2987] = 32'he2b0ee00;
    ram_cell[    2988] = 32'h783c1fd9;
    ram_cell[    2989] = 32'h0a1ded26;
    ram_cell[    2990] = 32'hf9774003;
    ram_cell[    2991] = 32'h864faa46;
    ram_cell[    2992] = 32'h616dcb24;
    ram_cell[    2993] = 32'hf4baecaf;
    ram_cell[    2994] = 32'hf626a78e;
    ram_cell[    2995] = 32'hc1d768a4;
    ram_cell[    2996] = 32'h8628ac0f;
    ram_cell[    2997] = 32'h3a123ac5;
    ram_cell[    2998] = 32'h61957f4d;
    ram_cell[    2999] = 32'h41e3333d;
    ram_cell[    3000] = 32'hd90b234c;
    ram_cell[    3001] = 32'hb63a20e5;
    ram_cell[    3002] = 32'h200bd7e7;
    ram_cell[    3003] = 32'hb2511406;
    ram_cell[    3004] = 32'hc75b334a;
    ram_cell[    3005] = 32'he96ddcea;
    ram_cell[    3006] = 32'hf10dcf3f;
    ram_cell[    3007] = 32'hededbc12;
    ram_cell[    3008] = 32'h3482fc8a;
    ram_cell[    3009] = 32'hb9556f20;
    ram_cell[    3010] = 32'h93ac3483;
    ram_cell[    3011] = 32'h13790689;
    ram_cell[    3012] = 32'hfd75fdf0;
    ram_cell[    3013] = 32'h73aa292c;
    ram_cell[    3014] = 32'h5568c5a5;
    ram_cell[    3015] = 32'h510fe497;
    ram_cell[    3016] = 32'h792e8dc1;
    ram_cell[    3017] = 32'h4c7ab3de;
    ram_cell[    3018] = 32'hd1dc4bd5;
    ram_cell[    3019] = 32'h17a40748;
    ram_cell[    3020] = 32'h763614b5;
    ram_cell[    3021] = 32'h1c196a96;
    ram_cell[    3022] = 32'h8901665f;
    ram_cell[    3023] = 32'hc4a90585;
    ram_cell[    3024] = 32'h9cf954d1;
    ram_cell[    3025] = 32'h9e1e9b44;
    ram_cell[    3026] = 32'h3baeb198;
    ram_cell[    3027] = 32'he8552f29;
    ram_cell[    3028] = 32'h8e303d7c;
    ram_cell[    3029] = 32'h70c87cd1;
    ram_cell[    3030] = 32'h648857d0;
    ram_cell[    3031] = 32'h3eb2fa26;
    ram_cell[    3032] = 32'heece0a46;
    ram_cell[    3033] = 32'hc86f5c83;
    ram_cell[    3034] = 32'h225caac4;
    ram_cell[    3035] = 32'hfab115b4;
    ram_cell[    3036] = 32'h0b2bad39;
    ram_cell[    3037] = 32'hfb22e41d;
    ram_cell[    3038] = 32'h7b493e93;
    ram_cell[    3039] = 32'h399dd841;
    ram_cell[    3040] = 32'he1794f55;
    ram_cell[    3041] = 32'h0d027771;
    ram_cell[    3042] = 32'hc18ca9a1;
    ram_cell[    3043] = 32'ha892d68e;
    ram_cell[    3044] = 32'ha3739b9a;
    ram_cell[    3045] = 32'h58f9c1d3;
    ram_cell[    3046] = 32'h09d57183;
    ram_cell[    3047] = 32'h747c5aaa;
    ram_cell[    3048] = 32'h1bbf38ae;
    ram_cell[    3049] = 32'h5595e7b5;
    ram_cell[    3050] = 32'h0f654fd6;
    ram_cell[    3051] = 32'h84e52dee;
    ram_cell[    3052] = 32'h9270e09d;
    ram_cell[    3053] = 32'hb0d68b4d;
    ram_cell[    3054] = 32'h195316f1;
    ram_cell[    3055] = 32'h2394bf0c;
    ram_cell[    3056] = 32'h8bda2e31;
    ram_cell[    3057] = 32'h1d9d9b5b;
    ram_cell[    3058] = 32'hce616b62;
    ram_cell[    3059] = 32'hfbce2330;
    ram_cell[    3060] = 32'h433b110d;
    ram_cell[    3061] = 32'h51a9d1ec;
    ram_cell[    3062] = 32'h95247fdb;
    ram_cell[    3063] = 32'h829d2e96;
    ram_cell[    3064] = 32'h12b8793d;
    ram_cell[    3065] = 32'hc832ed49;
    ram_cell[    3066] = 32'hbe7bcf7e;
    ram_cell[    3067] = 32'h52017e9a;
    ram_cell[    3068] = 32'h3edac005;
    ram_cell[    3069] = 32'h7747536e;
    ram_cell[    3070] = 32'hee2c35a2;
    ram_cell[    3071] = 32'h464bb547;
end

endmodule



module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h9a446be4;
    ram_cell[       1] = 32'h0;  // 32'h6c211748;
    ram_cell[       2] = 32'h0;  // 32'h56a91f67;
    ram_cell[       3] = 32'h0;  // 32'h2547b0f7;
    ram_cell[       4] = 32'h0;  // 32'h275853fa;
    ram_cell[       5] = 32'h0;  // 32'hf36b55f6;
    ram_cell[       6] = 32'h0;  // 32'h8100eb96;
    ram_cell[       7] = 32'h0;  // 32'h8b3b3d11;
    ram_cell[       8] = 32'h0;  // 32'h4879d4db;
    ram_cell[       9] = 32'h0;  // 32'hfd826dd9;
    ram_cell[      10] = 32'h0;  // 32'hca26ef65;
    ram_cell[      11] = 32'h0;  // 32'h865127c0;
    ram_cell[      12] = 32'h0;  // 32'h6b591b79;
    ram_cell[      13] = 32'h0;  // 32'h6653eef2;
    ram_cell[      14] = 32'h0;  // 32'he9a8beab;
    ram_cell[      15] = 32'h0;  // 32'h5c965bf0;
    ram_cell[      16] = 32'h0;  // 32'h8d93995b;
    ram_cell[      17] = 32'h0;  // 32'hfb2c6b4e;
    ram_cell[      18] = 32'h0;  // 32'h047d8981;
    ram_cell[      19] = 32'h0;  // 32'h8056c228;
    ram_cell[      20] = 32'h0;  // 32'hf13b3b6d;
    ram_cell[      21] = 32'h0;  // 32'h4886a1f8;
    ram_cell[      22] = 32'h0;  // 32'hd03d9e12;
    ram_cell[      23] = 32'h0;  // 32'h26298c3c;
    ram_cell[      24] = 32'h0;  // 32'h1685fd3b;
    ram_cell[      25] = 32'h0;  // 32'h0eb44305;
    ram_cell[      26] = 32'h0;  // 32'hcd73e7b8;
    ram_cell[      27] = 32'h0;  // 32'haf6d8532;
    ram_cell[      28] = 32'h0;  // 32'h8dbc8986;
    ram_cell[      29] = 32'h0;  // 32'ha68e70e8;
    ram_cell[      30] = 32'h0;  // 32'h03b03dcd;
    ram_cell[      31] = 32'h0;  // 32'hf34d86c3;
    ram_cell[      32] = 32'h0;  // 32'h0079ab9c;
    ram_cell[      33] = 32'h0;  // 32'h2addcacb;
    ram_cell[      34] = 32'h0;  // 32'h687a2353;
    ram_cell[      35] = 32'h0;  // 32'ha2693e98;
    ram_cell[      36] = 32'h0;  // 32'hda0f5895;
    ram_cell[      37] = 32'h0;  // 32'h787436e1;
    ram_cell[      38] = 32'h0;  // 32'hc98a7b18;
    ram_cell[      39] = 32'h0;  // 32'h55cbc6ac;
    ram_cell[      40] = 32'h0;  // 32'h9a6bd8f3;
    ram_cell[      41] = 32'h0;  // 32'hddea0b38;
    ram_cell[      42] = 32'h0;  // 32'h214982cc;
    ram_cell[      43] = 32'h0;  // 32'h48822389;
    ram_cell[      44] = 32'h0;  // 32'h8a257fba;
    ram_cell[      45] = 32'h0;  // 32'h46188a21;
    ram_cell[      46] = 32'h0;  // 32'hb3621b68;
    ram_cell[      47] = 32'h0;  // 32'h284f58c4;
    ram_cell[      48] = 32'h0;  // 32'h6d098e93;
    ram_cell[      49] = 32'h0;  // 32'h422b795c;
    ram_cell[      50] = 32'h0;  // 32'hc3b38a09;
    ram_cell[      51] = 32'h0;  // 32'h2af0d391;
    ram_cell[      52] = 32'h0;  // 32'h56ac24be;
    ram_cell[      53] = 32'h0;  // 32'hc3a6d6b8;
    ram_cell[      54] = 32'h0;  // 32'hcd887e06;
    ram_cell[      55] = 32'h0;  // 32'h807043db;
    ram_cell[      56] = 32'h0;  // 32'h1273178f;
    ram_cell[      57] = 32'h0;  // 32'h0e0d6157;
    ram_cell[      58] = 32'h0;  // 32'h11c38499;
    ram_cell[      59] = 32'h0;  // 32'hb29e0614;
    ram_cell[      60] = 32'h0;  // 32'hf3631ee8;
    ram_cell[      61] = 32'h0;  // 32'hf55dcf1a;
    ram_cell[      62] = 32'h0;  // 32'h31a94790;
    ram_cell[      63] = 32'h0;  // 32'hbba16e84;
    ram_cell[      64] = 32'h0;  // 32'h3bfb5834;
    ram_cell[      65] = 32'h0;  // 32'h467d0e1f;
    ram_cell[      66] = 32'h0;  // 32'h1452385d;
    ram_cell[      67] = 32'h0;  // 32'hcd0e7d36;
    ram_cell[      68] = 32'h0;  // 32'he1e48cd3;
    ram_cell[      69] = 32'h0;  // 32'hdf5771e3;
    ram_cell[      70] = 32'h0;  // 32'h1b99bc7c;
    ram_cell[      71] = 32'h0;  // 32'h8b17710a;
    ram_cell[      72] = 32'h0;  // 32'hbffef6df;
    ram_cell[      73] = 32'h0;  // 32'h7685b7b4;
    ram_cell[      74] = 32'h0;  // 32'h7526be56;
    ram_cell[      75] = 32'h0;  // 32'hc46789cf;
    ram_cell[      76] = 32'h0;  // 32'hfaddc6ec;
    ram_cell[      77] = 32'h0;  // 32'h410a875b;
    ram_cell[      78] = 32'h0;  // 32'haca87b1c;
    ram_cell[      79] = 32'h0;  // 32'h0d9bf880;
    ram_cell[      80] = 32'h0;  // 32'h84c00f8a;
    ram_cell[      81] = 32'h0;  // 32'h8d5fe7e6;
    ram_cell[      82] = 32'h0;  // 32'h1984e7d8;
    ram_cell[      83] = 32'h0;  // 32'h50ebafdf;
    ram_cell[      84] = 32'h0;  // 32'h61590d1b;
    ram_cell[      85] = 32'h0;  // 32'h2b316c86;
    ram_cell[      86] = 32'h0;  // 32'h417c7b32;
    ram_cell[      87] = 32'h0;  // 32'h2ab9437e;
    ram_cell[      88] = 32'h0;  // 32'hdef7150c;
    ram_cell[      89] = 32'h0;  // 32'h8dbe4563;
    ram_cell[      90] = 32'h0;  // 32'hb7eb6bc6;
    ram_cell[      91] = 32'h0;  // 32'h182ef961;
    ram_cell[      92] = 32'h0;  // 32'h28e8693c;
    ram_cell[      93] = 32'h0;  // 32'hf61a2225;
    ram_cell[      94] = 32'h0;  // 32'ha0693404;
    ram_cell[      95] = 32'h0;  // 32'ha8af07ea;
    ram_cell[      96] = 32'h0;  // 32'ha5aa762c;
    ram_cell[      97] = 32'h0;  // 32'h1b0bd043;
    ram_cell[      98] = 32'h0;  // 32'h74f3351a;
    ram_cell[      99] = 32'h0;  // 32'h0f6d5664;
    ram_cell[     100] = 32'h0;  // 32'h7b3a17fd;
    ram_cell[     101] = 32'h0;  // 32'h8ba90397;
    ram_cell[     102] = 32'h0;  // 32'ha8ee1e2a;
    ram_cell[     103] = 32'h0;  // 32'h85eac693;
    ram_cell[     104] = 32'h0;  // 32'he75500b3;
    ram_cell[     105] = 32'h0;  // 32'h66363317;
    ram_cell[     106] = 32'h0;  // 32'h5dc4737d;
    ram_cell[     107] = 32'h0;  // 32'h7efe9895;
    ram_cell[     108] = 32'h0;  // 32'h12adbb48;
    ram_cell[     109] = 32'h0;  // 32'hf2684dbd;
    ram_cell[     110] = 32'h0;  // 32'h4ef0f521;
    ram_cell[     111] = 32'h0;  // 32'h3067d267;
    ram_cell[     112] = 32'h0;  // 32'h36bb9301;
    ram_cell[     113] = 32'h0;  // 32'hcd931de1;
    ram_cell[     114] = 32'h0;  // 32'h7604fc97;
    ram_cell[     115] = 32'h0;  // 32'h9b413a56;
    ram_cell[     116] = 32'h0;  // 32'hbf46ae19;
    ram_cell[     117] = 32'h0;  // 32'h2fad20d6;
    ram_cell[     118] = 32'h0;  // 32'h2211bf45;
    ram_cell[     119] = 32'h0;  // 32'h8dadd34b;
    ram_cell[     120] = 32'h0;  // 32'h9484d848;
    ram_cell[     121] = 32'h0;  // 32'h71dcfdbb;
    ram_cell[     122] = 32'h0;  // 32'h90d8487d;
    ram_cell[     123] = 32'h0;  // 32'h5f6da8b1;
    ram_cell[     124] = 32'h0;  // 32'h4901f138;
    ram_cell[     125] = 32'h0;  // 32'h03692341;
    ram_cell[     126] = 32'h0;  // 32'h5bfe3e21;
    ram_cell[     127] = 32'h0;  // 32'h02821040;
    ram_cell[     128] = 32'h0;  // 32'heafc9b67;
    ram_cell[     129] = 32'h0;  // 32'h82eca1bd;
    ram_cell[     130] = 32'h0;  // 32'h274b771f;
    ram_cell[     131] = 32'h0;  // 32'hcb6582b3;
    ram_cell[     132] = 32'h0;  // 32'h75dccab0;
    ram_cell[     133] = 32'h0;  // 32'hb6f54c47;
    ram_cell[     134] = 32'h0;  // 32'h3ca13a51;
    ram_cell[     135] = 32'h0;  // 32'hf6b02130;
    ram_cell[     136] = 32'h0;  // 32'h5f91b598;
    ram_cell[     137] = 32'h0;  // 32'haf5731ad;
    ram_cell[     138] = 32'h0;  // 32'h86841a5a;
    ram_cell[     139] = 32'h0;  // 32'h2909639a;
    ram_cell[     140] = 32'h0;  // 32'ha159d17b;
    ram_cell[     141] = 32'h0;  // 32'he332412d;
    ram_cell[     142] = 32'h0;  // 32'h7ebc7d27;
    ram_cell[     143] = 32'h0;  // 32'h7afcb9f8;
    ram_cell[     144] = 32'h0;  // 32'h31b58c05;
    ram_cell[     145] = 32'h0;  // 32'hc5fc2637;
    ram_cell[     146] = 32'h0;  // 32'hfbef1def;
    ram_cell[     147] = 32'h0;  // 32'h727fd008;
    ram_cell[     148] = 32'h0;  // 32'ha57199ca;
    ram_cell[     149] = 32'h0;  // 32'h3a4f4fce;
    ram_cell[     150] = 32'h0;  // 32'he1a87d7d;
    ram_cell[     151] = 32'h0;  // 32'hed706cf0;
    ram_cell[     152] = 32'h0;  // 32'h9bc1f463;
    ram_cell[     153] = 32'h0;  // 32'hab49a469;
    ram_cell[     154] = 32'h0;  // 32'hf0885c33;
    ram_cell[     155] = 32'h0;  // 32'hee24573e;
    ram_cell[     156] = 32'h0;  // 32'hc26edf0f;
    ram_cell[     157] = 32'h0;  // 32'he7122d9c;
    ram_cell[     158] = 32'h0;  // 32'h0a9f1c1c;
    ram_cell[     159] = 32'h0;  // 32'h0d5a9623;
    ram_cell[     160] = 32'h0;  // 32'h887ddeab;
    ram_cell[     161] = 32'h0;  // 32'h0be3d4a9;
    ram_cell[     162] = 32'h0;  // 32'hb1259506;
    ram_cell[     163] = 32'h0;  // 32'hf4221469;
    ram_cell[     164] = 32'h0;  // 32'ha5e4480b;
    ram_cell[     165] = 32'h0;  // 32'h0a76fa4b;
    ram_cell[     166] = 32'h0;  // 32'hdcd3e5df;
    ram_cell[     167] = 32'h0;  // 32'hdcd26ad8;
    ram_cell[     168] = 32'h0;  // 32'h1416772f;
    ram_cell[     169] = 32'h0;  // 32'hc468043c;
    ram_cell[     170] = 32'h0;  // 32'h74d5a891;
    ram_cell[     171] = 32'h0;  // 32'h8f86f7cd;
    ram_cell[     172] = 32'h0;  // 32'h686b7466;
    ram_cell[     173] = 32'h0;  // 32'h1aa2632b;
    ram_cell[     174] = 32'h0;  // 32'hab05f71e;
    ram_cell[     175] = 32'h0;  // 32'h05d6cc8d;
    ram_cell[     176] = 32'h0;  // 32'h271044e6;
    ram_cell[     177] = 32'h0;  // 32'h4baa746b;
    ram_cell[     178] = 32'h0;  // 32'h52ed854a;
    ram_cell[     179] = 32'h0;  // 32'h7ca8f361;
    ram_cell[     180] = 32'h0;  // 32'h73c68e45;
    ram_cell[     181] = 32'h0;  // 32'h16a312cb;
    ram_cell[     182] = 32'h0;  // 32'hf5128fd4;
    ram_cell[     183] = 32'h0;  // 32'hc9d8b863;
    ram_cell[     184] = 32'h0;  // 32'hb1a5d0fd;
    ram_cell[     185] = 32'h0;  // 32'hf5c7017a;
    ram_cell[     186] = 32'h0;  // 32'he357696c;
    ram_cell[     187] = 32'h0;  // 32'h08a6a8ae;
    ram_cell[     188] = 32'h0;  // 32'ha5bd6e9b;
    ram_cell[     189] = 32'h0;  // 32'hfd003cc0;
    ram_cell[     190] = 32'h0;  // 32'h10eb5c81;
    ram_cell[     191] = 32'h0;  // 32'hcde8b598;
    ram_cell[     192] = 32'h0;  // 32'h8b1907ae;
    ram_cell[     193] = 32'h0;  // 32'he13785c2;
    ram_cell[     194] = 32'h0;  // 32'hc6d4667e;
    ram_cell[     195] = 32'h0;  // 32'h82b3c4df;
    ram_cell[     196] = 32'h0;  // 32'ha3d82642;
    ram_cell[     197] = 32'h0;  // 32'h9bf1a645;
    ram_cell[     198] = 32'h0;  // 32'h9c51823d;
    ram_cell[     199] = 32'h0;  // 32'h4250e147;
    ram_cell[     200] = 32'h0;  // 32'h40ea6a46;
    ram_cell[     201] = 32'h0;  // 32'h7eb87f36;
    ram_cell[     202] = 32'h0;  // 32'h74ae8908;
    ram_cell[     203] = 32'h0;  // 32'hf7ddb51c;
    ram_cell[     204] = 32'h0;  // 32'h7b2092c4;
    ram_cell[     205] = 32'h0;  // 32'h0f158739;
    ram_cell[     206] = 32'h0;  // 32'h61679ac2;
    ram_cell[     207] = 32'h0;  // 32'h76d4989d;
    ram_cell[     208] = 32'h0;  // 32'hef124ecd;
    ram_cell[     209] = 32'h0;  // 32'h2abd1661;
    ram_cell[     210] = 32'h0;  // 32'h05414d56;
    ram_cell[     211] = 32'h0;  // 32'h4618d87d;
    ram_cell[     212] = 32'h0;  // 32'ha90439fe;
    ram_cell[     213] = 32'h0;  // 32'h1440b16e;
    ram_cell[     214] = 32'h0;  // 32'h526cf005;
    ram_cell[     215] = 32'h0;  // 32'h9a7e471b;
    ram_cell[     216] = 32'h0;  // 32'h61f24a20;
    ram_cell[     217] = 32'h0;  // 32'ha6a23c27;
    ram_cell[     218] = 32'h0;  // 32'h48d4f021;
    ram_cell[     219] = 32'h0;  // 32'hc843f3bf;
    ram_cell[     220] = 32'h0;  // 32'h3fef1389;
    ram_cell[     221] = 32'h0;  // 32'h29151f34;
    ram_cell[     222] = 32'h0;  // 32'h5a177484;
    ram_cell[     223] = 32'h0;  // 32'h7cc20703;
    ram_cell[     224] = 32'h0;  // 32'hcb402e14;
    ram_cell[     225] = 32'h0;  // 32'h42bb059f;
    ram_cell[     226] = 32'h0;  // 32'h9c1c06af;
    ram_cell[     227] = 32'h0;  // 32'h10ad7a6e;
    ram_cell[     228] = 32'h0;  // 32'h80dfff5a;
    ram_cell[     229] = 32'h0;  // 32'he14461f3;
    ram_cell[     230] = 32'h0;  // 32'hafc547a6;
    ram_cell[     231] = 32'h0;  // 32'h425d1fb0;
    ram_cell[     232] = 32'h0;  // 32'he1848f0a;
    ram_cell[     233] = 32'h0;  // 32'h625bd8cd;
    ram_cell[     234] = 32'h0;  // 32'hb668673c;
    ram_cell[     235] = 32'h0;  // 32'h90b2ff36;
    ram_cell[     236] = 32'h0;  // 32'h6049d1bd;
    ram_cell[     237] = 32'h0;  // 32'h16dadf67;
    ram_cell[     238] = 32'h0;  // 32'hf44f9ff4;
    ram_cell[     239] = 32'h0;  // 32'h596514c0;
    ram_cell[     240] = 32'h0;  // 32'h6d99d9a0;
    ram_cell[     241] = 32'h0;  // 32'h6f361f1c;
    ram_cell[     242] = 32'h0;  // 32'h2fa331f6;
    ram_cell[     243] = 32'h0;  // 32'h3905706e;
    ram_cell[     244] = 32'h0;  // 32'h2f14e0f9;
    ram_cell[     245] = 32'h0;  // 32'hed32540f;
    ram_cell[     246] = 32'h0;  // 32'h60d0d112;
    ram_cell[     247] = 32'h0;  // 32'hd96e2ba3;
    ram_cell[     248] = 32'h0;  // 32'hc5f565a1;
    ram_cell[     249] = 32'h0;  // 32'h4497afaf;
    ram_cell[     250] = 32'h0;  // 32'h584a075a;
    ram_cell[     251] = 32'h0;  // 32'h761f4828;
    ram_cell[     252] = 32'h0;  // 32'h7596bf9b;
    ram_cell[     253] = 32'h0;  // 32'h678e54cf;
    ram_cell[     254] = 32'h0;  // 32'ha2626c13;
    ram_cell[     255] = 32'h0;  // 32'h86a59710;
    ram_cell[     256] = 32'h0;  // 32'h7c091f55;
    ram_cell[     257] = 32'h0;  // 32'h3adb9701;
    ram_cell[     258] = 32'h0;  // 32'h2bbf0edc;
    ram_cell[     259] = 32'h0;  // 32'hbef4f218;
    ram_cell[     260] = 32'h0;  // 32'h1db747d4;
    ram_cell[     261] = 32'h0;  // 32'h7ecdf36f;
    ram_cell[     262] = 32'h0;  // 32'h9349ca1e;
    ram_cell[     263] = 32'h0;  // 32'h6dd5a79c;
    ram_cell[     264] = 32'h0;  // 32'h4f10f2e1;
    ram_cell[     265] = 32'h0;  // 32'h24ded3a1;
    ram_cell[     266] = 32'h0;  // 32'h48020259;
    ram_cell[     267] = 32'h0;  // 32'h57bb43c5;
    ram_cell[     268] = 32'h0;  // 32'h0b798279;
    ram_cell[     269] = 32'h0;  // 32'h788ed019;
    ram_cell[     270] = 32'h0;  // 32'h662a2037;
    ram_cell[     271] = 32'h0;  // 32'h0039e821;
    ram_cell[     272] = 32'h0;  // 32'h32b97ef1;
    ram_cell[     273] = 32'h0;  // 32'h5dca3745;
    ram_cell[     274] = 32'h0;  // 32'h61485327;
    ram_cell[     275] = 32'h0;  // 32'h3e1c6a74;
    ram_cell[     276] = 32'h0;  // 32'hb57d2759;
    ram_cell[     277] = 32'h0;  // 32'h06b4f2d4;
    ram_cell[     278] = 32'h0;  // 32'h2261a35c;
    ram_cell[     279] = 32'h0;  // 32'h3135fd8f;
    ram_cell[     280] = 32'h0;  // 32'h01fed23a;
    ram_cell[     281] = 32'h0;  // 32'h27937b6b;
    ram_cell[     282] = 32'h0;  // 32'h4dbaadfc;
    ram_cell[     283] = 32'h0;  // 32'h9d884ff4;
    ram_cell[     284] = 32'h0;  // 32'h3768b6d9;
    ram_cell[     285] = 32'h0;  // 32'heff74a47;
    ram_cell[     286] = 32'h0;  // 32'h7531d904;
    ram_cell[     287] = 32'h0;  // 32'h839a9c03;
    ram_cell[     288] = 32'h0;  // 32'h28c529f7;
    ram_cell[     289] = 32'h0;  // 32'h0fb5cda2;
    ram_cell[     290] = 32'h0;  // 32'h2a475afc;
    ram_cell[     291] = 32'h0;  // 32'h02f2fb07;
    ram_cell[     292] = 32'h0;  // 32'h4060d455;
    ram_cell[     293] = 32'h0;  // 32'h761f9544;
    ram_cell[     294] = 32'h0;  // 32'hcbc21491;
    ram_cell[     295] = 32'h0;  // 32'hbc74f51f;
    ram_cell[     296] = 32'h0;  // 32'h81de672c;
    ram_cell[     297] = 32'h0;  // 32'he248680b;
    ram_cell[     298] = 32'h0;  // 32'hec8f27ff;
    ram_cell[     299] = 32'h0;  // 32'h44f60cf8;
    ram_cell[     300] = 32'h0;  // 32'h7c375a00;
    ram_cell[     301] = 32'h0;  // 32'h2f80f56f;
    ram_cell[     302] = 32'h0;  // 32'ha987ed0e;
    ram_cell[     303] = 32'h0;  // 32'hfe0b7748;
    ram_cell[     304] = 32'h0;  // 32'hf5b35f80;
    ram_cell[     305] = 32'h0;  // 32'h5e9b9b30;
    ram_cell[     306] = 32'h0;  // 32'hde8e1e13;
    ram_cell[     307] = 32'h0;  // 32'ha21f69ed;
    ram_cell[     308] = 32'h0;  // 32'h33e0f36b;
    ram_cell[     309] = 32'h0;  // 32'h149504d8;
    ram_cell[     310] = 32'h0;  // 32'h12ab2118;
    ram_cell[     311] = 32'h0;  // 32'he3343d2b;
    ram_cell[     312] = 32'h0;  // 32'hc6bda3a3;
    ram_cell[     313] = 32'h0;  // 32'h8527db15;
    ram_cell[     314] = 32'h0;  // 32'hd6a8ea2c;
    ram_cell[     315] = 32'h0;  // 32'h160275cf;
    ram_cell[     316] = 32'h0;  // 32'hdb0bf639;
    ram_cell[     317] = 32'h0;  // 32'h094c7adc;
    ram_cell[     318] = 32'h0;  // 32'h0d16d7e8;
    ram_cell[     319] = 32'h0;  // 32'h0548f7c4;
    ram_cell[     320] = 32'h0;  // 32'h2457a585;
    ram_cell[     321] = 32'h0;  // 32'h4ec7a836;
    ram_cell[     322] = 32'h0;  // 32'h26b07792;
    ram_cell[     323] = 32'h0;  // 32'hdf6757e8;
    ram_cell[     324] = 32'h0;  // 32'hc3cf46a1;
    ram_cell[     325] = 32'h0;  // 32'h81a82ec8;
    ram_cell[     326] = 32'h0;  // 32'hddb36cef;
    ram_cell[     327] = 32'h0;  // 32'h674a12be;
    ram_cell[     328] = 32'h0;  // 32'h17214421;
    ram_cell[     329] = 32'h0;  // 32'h9d21eb4a;
    ram_cell[     330] = 32'h0;  // 32'hf5622d69;
    ram_cell[     331] = 32'h0;  // 32'h9d3b5171;
    ram_cell[     332] = 32'h0;  // 32'hb2ca8292;
    ram_cell[     333] = 32'h0;  // 32'h94d81777;
    ram_cell[     334] = 32'h0;  // 32'hee671bc4;
    ram_cell[     335] = 32'h0;  // 32'hed404d88;
    ram_cell[     336] = 32'h0;  // 32'hed6b8710;
    ram_cell[     337] = 32'h0;  // 32'hfae7a628;
    ram_cell[     338] = 32'h0;  // 32'h028515f3;
    ram_cell[     339] = 32'h0;  // 32'had0c34ca;
    ram_cell[     340] = 32'h0;  // 32'hefecb4fe;
    ram_cell[     341] = 32'h0;  // 32'hb4fb1fd1;
    ram_cell[     342] = 32'h0;  // 32'he2ada1a9;
    ram_cell[     343] = 32'h0;  // 32'he91ae967;
    ram_cell[     344] = 32'h0;  // 32'hfe97ac5e;
    ram_cell[     345] = 32'h0;  // 32'h8c9b544c;
    ram_cell[     346] = 32'h0;  // 32'hfd76d0c4;
    ram_cell[     347] = 32'h0;  // 32'h138a19f9;
    ram_cell[     348] = 32'h0;  // 32'h2901c130;
    ram_cell[     349] = 32'h0;  // 32'h88cc0167;
    ram_cell[     350] = 32'h0;  // 32'hceac22f5;
    ram_cell[     351] = 32'h0;  // 32'h5866799d;
    ram_cell[     352] = 32'h0;  // 32'hb233b1cb;
    ram_cell[     353] = 32'h0;  // 32'h585dbe1e;
    ram_cell[     354] = 32'h0;  // 32'ha886dfe9;
    ram_cell[     355] = 32'h0;  // 32'hc6de4585;
    ram_cell[     356] = 32'h0;  // 32'hb970c228;
    ram_cell[     357] = 32'h0;  // 32'hee348ac0;
    ram_cell[     358] = 32'h0;  // 32'h5c859db0;
    ram_cell[     359] = 32'h0;  // 32'hd0ddbbba;
    ram_cell[     360] = 32'h0;  // 32'h68820e15;
    ram_cell[     361] = 32'h0;  // 32'ha9c56230;
    ram_cell[     362] = 32'h0;  // 32'hf91d0dcb;
    ram_cell[     363] = 32'h0;  // 32'hb22de4f3;
    ram_cell[     364] = 32'h0;  // 32'h07101e9e;
    ram_cell[     365] = 32'h0;  // 32'hef83f554;
    ram_cell[     366] = 32'h0;  // 32'h37f9ab2d;
    ram_cell[     367] = 32'h0;  // 32'hca6d6559;
    ram_cell[     368] = 32'h0;  // 32'ha7185d03;
    ram_cell[     369] = 32'h0;  // 32'h39001701;
    ram_cell[     370] = 32'h0;  // 32'h1f5eb657;
    ram_cell[     371] = 32'h0;  // 32'h52f80ed7;
    ram_cell[     372] = 32'h0;  // 32'h29f95fc2;
    ram_cell[     373] = 32'h0;  // 32'h5bea27ad;
    ram_cell[     374] = 32'h0;  // 32'hd0fef7f8;
    ram_cell[     375] = 32'h0;  // 32'h06fd0b4c;
    ram_cell[     376] = 32'h0;  // 32'h0d85ef3a;
    ram_cell[     377] = 32'h0;  // 32'h820091db;
    ram_cell[     378] = 32'h0;  // 32'hc2dcd41f;
    ram_cell[     379] = 32'h0;  // 32'h10adc5eb;
    ram_cell[     380] = 32'h0;  // 32'hb14ec4f4;
    ram_cell[     381] = 32'h0;  // 32'hdef6233b;
    ram_cell[     382] = 32'h0;  // 32'h977481c4;
    ram_cell[     383] = 32'h0;  // 32'hf4bf76ed;
    ram_cell[     384] = 32'h0;  // 32'hda5a8156;
    ram_cell[     385] = 32'h0;  // 32'hf40409b0;
    ram_cell[     386] = 32'h0;  // 32'h8e17bac4;
    ram_cell[     387] = 32'h0;  // 32'hd520a7ea;
    ram_cell[     388] = 32'h0;  // 32'h1b1ebd3b;
    ram_cell[     389] = 32'h0;  // 32'h2c3b39a8;
    ram_cell[     390] = 32'h0;  // 32'hb5cb3154;
    ram_cell[     391] = 32'h0;  // 32'h2599c42a;
    ram_cell[     392] = 32'h0;  // 32'h1c72fd5b;
    ram_cell[     393] = 32'h0;  // 32'h424d9b0f;
    ram_cell[     394] = 32'h0;  // 32'hb5d23cd1;
    ram_cell[     395] = 32'h0;  // 32'h3d1c87e6;
    ram_cell[     396] = 32'h0;  // 32'h39b9bd6e;
    ram_cell[     397] = 32'h0;  // 32'h23e6d86a;
    ram_cell[     398] = 32'h0;  // 32'h429d3051;
    ram_cell[     399] = 32'h0;  // 32'h17a8cd02;
    ram_cell[     400] = 32'h0;  // 32'h9c57d3de;
    ram_cell[     401] = 32'h0;  // 32'he445a280;
    ram_cell[     402] = 32'h0;  // 32'h983f3385;
    ram_cell[     403] = 32'h0;  // 32'h08b77822;
    ram_cell[     404] = 32'h0;  // 32'ha1d684f0;
    ram_cell[     405] = 32'h0;  // 32'h0a23fbca;
    ram_cell[     406] = 32'h0;  // 32'h15843c64;
    ram_cell[     407] = 32'h0;  // 32'h692a324c;
    ram_cell[     408] = 32'h0;  // 32'h48905660;
    ram_cell[     409] = 32'h0;  // 32'h85afff8b;
    ram_cell[     410] = 32'h0;  // 32'h79b31db7;
    ram_cell[     411] = 32'h0;  // 32'h36acd1a9;
    ram_cell[     412] = 32'h0;  // 32'had2873dc;
    ram_cell[     413] = 32'h0;  // 32'h53f79960;
    ram_cell[     414] = 32'h0;  // 32'hbf050ef9;
    ram_cell[     415] = 32'h0;  // 32'ha75e8d3d;
    ram_cell[     416] = 32'h0;  // 32'hb367447e;
    ram_cell[     417] = 32'h0;  // 32'h681300cd;
    ram_cell[     418] = 32'h0;  // 32'hff3b3900;
    ram_cell[     419] = 32'h0;  // 32'hd1a70df5;
    ram_cell[     420] = 32'h0;  // 32'ha2518567;
    ram_cell[     421] = 32'h0;  // 32'h53893786;
    ram_cell[     422] = 32'h0;  // 32'hfd902aa1;
    ram_cell[     423] = 32'h0;  // 32'hfff6d8b6;
    ram_cell[     424] = 32'h0;  // 32'h04d8877a;
    ram_cell[     425] = 32'h0;  // 32'h3eb98d75;
    ram_cell[     426] = 32'h0;  // 32'h0c81a6f1;
    ram_cell[     427] = 32'h0;  // 32'h4e03eb2e;
    ram_cell[     428] = 32'h0;  // 32'ha0ca17a1;
    ram_cell[     429] = 32'h0;  // 32'hc63f1af8;
    ram_cell[     430] = 32'h0;  // 32'h30219a40;
    ram_cell[     431] = 32'h0;  // 32'h731a82fe;
    ram_cell[     432] = 32'h0;  // 32'h6caaf934;
    ram_cell[     433] = 32'h0;  // 32'h57a93651;
    ram_cell[     434] = 32'h0;  // 32'h14337196;
    ram_cell[     435] = 32'h0;  // 32'h44b9ddad;
    ram_cell[     436] = 32'h0;  // 32'h4150ff0e;
    ram_cell[     437] = 32'h0;  // 32'h700baf10;
    ram_cell[     438] = 32'h0;  // 32'h9a2d8732;
    ram_cell[     439] = 32'h0;  // 32'h0c90fb55;
    ram_cell[     440] = 32'h0;  // 32'h522a924a;
    ram_cell[     441] = 32'h0;  // 32'hf3df7c40;
    ram_cell[     442] = 32'h0;  // 32'h5fd9a010;
    ram_cell[     443] = 32'h0;  // 32'haeec62b5;
    ram_cell[     444] = 32'h0;  // 32'hbd6cc033;
    ram_cell[     445] = 32'h0;  // 32'h945c6aaa;
    ram_cell[     446] = 32'h0;  // 32'h3271b30b;
    ram_cell[     447] = 32'h0;  // 32'h38fbc0a6;
    ram_cell[     448] = 32'h0;  // 32'hfeb76819;
    ram_cell[     449] = 32'h0;  // 32'h8cff508c;
    ram_cell[     450] = 32'h0;  // 32'h52547145;
    ram_cell[     451] = 32'h0;  // 32'h85306e59;
    ram_cell[     452] = 32'h0;  // 32'hb42ae923;
    ram_cell[     453] = 32'h0;  // 32'h86a8dc6a;
    ram_cell[     454] = 32'h0;  // 32'he49a614f;
    ram_cell[     455] = 32'h0;  // 32'h7061b0f6;
    ram_cell[     456] = 32'h0;  // 32'h521a9014;
    ram_cell[     457] = 32'h0;  // 32'h15e21684;
    ram_cell[     458] = 32'h0;  // 32'h2cc8958c;
    ram_cell[     459] = 32'h0;  // 32'h9f839b8c;
    ram_cell[     460] = 32'h0;  // 32'hd169624d;
    ram_cell[     461] = 32'h0;  // 32'h60779561;
    ram_cell[     462] = 32'h0;  // 32'h09b2f739;
    ram_cell[     463] = 32'h0;  // 32'h3cefaa80;
    ram_cell[     464] = 32'h0;  // 32'h76b70658;
    ram_cell[     465] = 32'h0;  // 32'h00f95b07;
    ram_cell[     466] = 32'h0;  // 32'hf9f0479a;
    ram_cell[     467] = 32'h0;  // 32'h94eb134d;
    ram_cell[     468] = 32'h0;  // 32'hd608a236;
    ram_cell[     469] = 32'h0;  // 32'ha0473bfd;
    ram_cell[     470] = 32'h0;  // 32'h11f80446;
    ram_cell[     471] = 32'h0;  // 32'h33150a72;
    ram_cell[     472] = 32'h0;  // 32'h96134468;
    ram_cell[     473] = 32'h0;  // 32'h32316275;
    ram_cell[     474] = 32'h0;  // 32'h2b48b47a;
    ram_cell[     475] = 32'h0;  // 32'h4a309ba8;
    ram_cell[     476] = 32'h0;  // 32'hbb6170cd;
    ram_cell[     477] = 32'h0;  // 32'h31996c0d;
    ram_cell[     478] = 32'h0;  // 32'h51390702;
    ram_cell[     479] = 32'h0;  // 32'hc43da6da;
    ram_cell[     480] = 32'h0;  // 32'h6172e375;
    ram_cell[     481] = 32'h0;  // 32'h6e701c2f;
    ram_cell[     482] = 32'h0;  // 32'h66bb9816;
    ram_cell[     483] = 32'h0;  // 32'hb0134628;
    ram_cell[     484] = 32'h0;  // 32'hdd0cc769;
    ram_cell[     485] = 32'h0;  // 32'h9e36b985;
    ram_cell[     486] = 32'h0;  // 32'hf80c3f0f;
    ram_cell[     487] = 32'h0;  // 32'h70f3b9c1;
    ram_cell[     488] = 32'h0;  // 32'hfbe6c42d;
    ram_cell[     489] = 32'h0;  // 32'h8cddb12a;
    ram_cell[     490] = 32'h0;  // 32'h9fb3e216;
    ram_cell[     491] = 32'h0;  // 32'hc4aa7c5e;
    ram_cell[     492] = 32'h0;  // 32'hb16d8052;
    ram_cell[     493] = 32'h0;  // 32'h52260977;
    ram_cell[     494] = 32'h0;  // 32'hd61a3fb8;
    ram_cell[     495] = 32'h0;  // 32'hb28a938b;
    ram_cell[     496] = 32'h0;  // 32'h01379cfe;
    ram_cell[     497] = 32'h0;  // 32'hd63d32b9;
    ram_cell[     498] = 32'h0;  // 32'had2b6e9b;
    ram_cell[     499] = 32'h0;  // 32'h23380bc5;
    ram_cell[     500] = 32'h0;  // 32'h518e039b;
    ram_cell[     501] = 32'h0;  // 32'hccb5ec51;
    ram_cell[     502] = 32'h0;  // 32'h7727784e;
    ram_cell[     503] = 32'h0;  // 32'he6c7be1b;
    ram_cell[     504] = 32'h0;  // 32'h6796eabe;
    ram_cell[     505] = 32'h0;  // 32'he816e5fe;
    ram_cell[     506] = 32'h0;  // 32'h964fff8d;
    ram_cell[     507] = 32'h0;  // 32'hc31df44a;
    ram_cell[     508] = 32'h0;  // 32'he774ac19;
    ram_cell[     509] = 32'h0;  // 32'ha8be7b4a;
    ram_cell[     510] = 32'h0;  // 32'h66146642;
    ram_cell[     511] = 32'h0;  // 32'hc3ce2bd7;
    ram_cell[     512] = 32'h0;  // 32'h58e3cc73;
    ram_cell[     513] = 32'h0;  // 32'hccedc4ce;
    ram_cell[     514] = 32'h0;  // 32'h75ad351c;
    ram_cell[     515] = 32'h0;  // 32'h17190139;
    ram_cell[     516] = 32'h0;  // 32'h66e4b800;
    ram_cell[     517] = 32'h0;  // 32'h1d67fb3a;
    ram_cell[     518] = 32'h0;  // 32'h34c97357;
    ram_cell[     519] = 32'h0;  // 32'h17dbd460;
    ram_cell[     520] = 32'h0;  // 32'hf2a21aa0;
    ram_cell[     521] = 32'h0;  // 32'h46259800;
    ram_cell[     522] = 32'h0;  // 32'h392078a2;
    ram_cell[     523] = 32'h0;  // 32'hc76ee3cf;
    ram_cell[     524] = 32'h0;  // 32'hb0121466;
    ram_cell[     525] = 32'h0;  // 32'h86fff9e6;
    ram_cell[     526] = 32'h0;  // 32'h95723596;
    ram_cell[     527] = 32'h0;  // 32'h65c9c985;
    ram_cell[     528] = 32'h0;  // 32'h2f27197b;
    ram_cell[     529] = 32'h0;  // 32'hdfe2babd;
    ram_cell[     530] = 32'h0;  // 32'hb5f73169;
    ram_cell[     531] = 32'h0;  // 32'h24185e77;
    ram_cell[     532] = 32'h0;  // 32'hd2ff40e7;
    ram_cell[     533] = 32'h0;  // 32'h7413cdee;
    ram_cell[     534] = 32'h0;  // 32'h4d3487e2;
    ram_cell[     535] = 32'h0;  // 32'h4724066c;
    ram_cell[     536] = 32'h0;  // 32'h36096627;
    ram_cell[     537] = 32'h0;  // 32'h7a007cbe;
    ram_cell[     538] = 32'h0;  // 32'hb03f5d6a;
    ram_cell[     539] = 32'h0;  // 32'h63c7bc7f;
    ram_cell[     540] = 32'h0;  // 32'h6c4fe4a6;
    ram_cell[     541] = 32'h0;  // 32'hce7728db;
    ram_cell[     542] = 32'h0;  // 32'h806b9a5e;
    ram_cell[     543] = 32'h0;  // 32'h2c866537;
    ram_cell[     544] = 32'h0;  // 32'hc69d2eae;
    ram_cell[     545] = 32'h0;  // 32'h7701b790;
    ram_cell[     546] = 32'h0;  // 32'hf271327f;
    ram_cell[     547] = 32'h0;  // 32'hf3a06e11;
    ram_cell[     548] = 32'h0;  // 32'h206934fc;
    ram_cell[     549] = 32'h0;  // 32'h0454b094;
    ram_cell[     550] = 32'h0;  // 32'h5abeaeaa;
    ram_cell[     551] = 32'h0;  // 32'h90db9444;
    ram_cell[     552] = 32'h0;  // 32'he4bc5f2e;
    ram_cell[     553] = 32'h0;  // 32'h76b24442;
    ram_cell[     554] = 32'h0;  // 32'h7c3e7bb4;
    ram_cell[     555] = 32'h0;  // 32'h5696f778;
    ram_cell[     556] = 32'h0;  // 32'hfc99883e;
    ram_cell[     557] = 32'h0;  // 32'h1f163267;
    ram_cell[     558] = 32'h0;  // 32'hae7c0ed6;
    ram_cell[     559] = 32'h0;  // 32'hdb367f9e;
    ram_cell[     560] = 32'h0;  // 32'hc8c9eab5;
    ram_cell[     561] = 32'h0;  // 32'h426e9e98;
    ram_cell[     562] = 32'h0;  // 32'h2875090b;
    ram_cell[     563] = 32'h0;  // 32'h1f4f0ff6;
    ram_cell[     564] = 32'h0;  // 32'h43c294eb;
    ram_cell[     565] = 32'h0;  // 32'h5513f1bf;
    ram_cell[     566] = 32'h0;  // 32'h70370b4b;
    ram_cell[     567] = 32'h0;  // 32'hd5391c54;
    ram_cell[     568] = 32'h0;  // 32'hd20b61e7;
    ram_cell[     569] = 32'h0;  // 32'hfe51baee;
    ram_cell[     570] = 32'h0;  // 32'hd4002338;
    ram_cell[     571] = 32'h0;  // 32'h9320a84d;
    ram_cell[     572] = 32'h0;  // 32'h6bc134ca;
    ram_cell[     573] = 32'h0;  // 32'h6d5d7ece;
    ram_cell[     574] = 32'h0;  // 32'he71b7df1;
    ram_cell[     575] = 32'h0;  // 32'h82e53c0c;
    ram_cell[     576] = 32'h0;  // 32'hba335ab8;
    ram_cell[     577] = 32'h0;  // 32'hc85cbc50;
    ram_cell[     578] = 32'h0;  // 32'hc8598f4e;
    ram_cell[     579] = 32'h0;  // 32'ha1e37a19;
    ram_cell[     580] = 32'h0;  // 32'h90417b1f;
    ram_cell[     581] = 32'h0;  // 32'h2b0ae0c2;
    ram_cell[     582] = 32'h0;  // 32'hbc289bca;
    ram_cell[     583] = 32'h0;  // 32'h6f6e3a4d;
    ram_cell[     584] = 32'h0;  // 32'h809af71b;
    ram_cell[     585] = 32'h0;  // 32'h0cab4ac2;
    ram_cell[     586] = 32'h0;  // 32'ha761788e;
    ram_cell[     587] = 32'h0;  // 32'he0ac9ec0;
    ram_cell[     588] = 32'h0;  // 32'h9058c5cd;
    ram_cell[     589] = 32'h0;  // 32'hbf4d9bd2;
    ram_cell[     590] = 32'h0;  // 32'h3edecfe4;
    ram_cell[     591] = 32'h0;  // 32'h35ee0176;
    ram_cell[     592] = 32'h0;  // 32'h3861d197;
    ram_cell[     593] = 32'h0;  // 32'h4eff0725;
    ram_cell[     594] = 32'h0;  // 32'h69a0a2d7;
    ram_cell[     595] = 32'h0;  // 32'he72b9460;
    ram_cell[     596] = 32'h0;  // 32'hbad05323;
    ram_cell[     597] = 32'h0;  // 32'h302db0ea;
    ram_cell[     598] = 32'h0;  // 32'h557a44bf;
    ram_cell[     599] = 32'h0;  // 32'hea7878c3;
    ram_cell[     600] = 32'h0;  // 32'hec5f8d3d;
    ram_cell[     601] = 32'h0;  // 32'h4774951c;
    ram_cell[     602] = 32'h0;  // 32'h4e30343e;
    ram_cell[     603] = 32'h0;  // 32'hdabd7223;
    ram_cell[     604] = 32'h0;  // 32'h50271577;
    ram_cell[     605] = 32'h0;  // 32'h4270c9d9;
    ram_cell[     606] = 32'h0;  // 32'h9fe0ff83;
    ram_cell[     607] = 32'h0;  // 32'h46f3f075;
    ram_cell[     608] = 32'h0;  // 32'h9371bbbd;
    ram_cell[     609] = 32'h0;  // 32'hfe77e262;
    ram_cell[     610] = 32'h0;  // 32'h5f067701;
    ram_cell[     611] = 32'h0;  // 32'h43e3118b;
    ram_cell[     612] = 32'h0;  // 32'h4ef31347;
    ram_cell[     613] = 32'h0;  // 32'h7113a8d8;
    ram_cell[     614] = 32'h0;  // 32'hb1c0ead7;
    ram_cell[     615] = 32'h0;  // 32'h86513d89;
    ram_cell[     616] = 32'h0;  // 32'hbc36015e;
    ram_cell[     617] = 32'h0;  // 32'h5a006db8;
    ram_cell[     618] = 32'h0;  // 32'hb4535e39;
    ram_cell[     619] = 32'h0;  // 32'h20a75fc8;
    ram_cell[     620] = 32'h0;  // 32'he5e6a7ee;
    ram_cell[     621] = 32'h0;  // 32'h76730ee7;
    ram_cell[     622] = 32'h0;  // 32'hef04f362;
    ram_cell[     623] = 32'h0;  // 32'h2d2e05c0;
    ram_cell[     624] = 32'h0;  // 32'h6c5a46d9;
    ram_cell[     625] = 32'h0;  // 32'haa8f05d6;
    ram_cell[     626] = 32'h0;  // 32'h9038bd63;
    ram_cell[     627] = 32'h0;  // 32'hd77f7226;
    ram_cell[     628] = 32'h0;  // 32'h235fbfb2;
    ram_cell[     629] = 32'h0;  // 32'hab8383ed;
    ram_cell[     630] = 32'h0;  // 32'h0b09a1a1;
    ram_cell[     631] = 32'h0;  // 32'h95b036a2;
    ram_cell[     632] = 32'h0;  // 32'haf8956cd;
    ram_cell[     633] = 32'h0;  // 32'hdea8d1f5;
    ram_cell[     634] = 32'h0;  // 32'he1d284a9;
    ram_cell[     635] = 32'h0;  // 32'h1755b56a;
    ram_cell[     636] = 32'h0;  // 32'h00b60fa9;
    ram_cell[     637] = 32'h0;  // 32'h4809d907;
    ram_cell[     638] = 32'h0;  // 32'hd7ea3c35;
    ram_cell[     639] = 32'h0;  // 32'hb7da6ff6;
    ram_cell[     640] = 32'h0;  // 32'haeb992a9;
    ram_cell[     641] = 32'h0;  // 32'h29e91990;
    ram_cell[     642] = 32'h0;  // 32'h28d6f7ee;
    ram_cell[     643] = 32'h0;  // 32'hce3d648f;
    ram_cell[     644] = 32'h0;  // 32'h3c6650df;
    ram_cell[     645] = 32'h0;  // 32'hdad257a0;
    ram_cell[     646] = 32'h0;  // 32'h37503b62;
    ram_cell[     647] = 32'h0;  // 32'h3fa92701;
    ram_cell[     648] = 32'h0;  // 32'h9ace48d0;
    ram_cell[     649] = 32'h0;  // 32'h5e39642a;
    ram_cell[     650] = 32'h0;  // 32'h28fbb0c9;
    ram_cell[     651] = 32'h0;  // 32'h2f145add;
    ram_cell[     652] = 32'h0;  // 32'h8cdc708e;
    ram_cell[     653] = 32'h0;  // 32'hf5894010;
    ram_cell[     654] = 32'h0;  // 32'h05f94790;
    ram_cell[     655] = 32'h0;  // 32'hf0fb3a9b;
    ram_cell[     656] = 32'h0;  // 32'h50265610;
    ram_cell[     657] = 32'h0;  // 32'hb95d8bbd;
    ram_cell[     658] = 32'h0;  // 32'h4e7a2fb7;
    ram_cell[     659] = 32'h0;  // 32'h21c13dc9;
    ram_cell[     660] = 32'h0;  // 32'hde9721d5;
    ram_cell[     661] = 32'h0;  // 32'hfbbf93cd;
    ram_cell[     662] = 32'h0;  // 32'hc9016d1f;
    ram_cell[     663] = 32'h0;  // 32'hba67a4df;
    ram_cell[     664] = 32'h0;  // 32'h09546189;
    ram_cell[     665] = 32'h0;  // 32'h28b9d361;
    ram_cell[     666] = 32'h0;  // 32'he63cda3f;
    ram_cell[     667] = 32'h0;  // 32'he1e2302c;
    ram_cell[     668] = 32'h0;  // 32'h3ef2aba7;
    ram_cell[     669] = 32'h0;  // 32'hb1d7b15f;
    ram_cell[     670] = 32'h0;  // 32'h4d26378a;
    ram_cell[     671] = 32'h0;  // 32'h7d8c7bd9;
    ram_cell[     672] = 32'h0;  // 32'h2c6d5372;
    ram_cell[     673] = 32'h0;  // 32'h8a198d10;
    ram_cell[     674] = 32'h0;  // 32'hb28530c9;
    ram_cell[     675] = 32'h0;  // 32'h1a0621cd;
    ram_cell[     676] = 32'h0;  // 32'h6a5aeadd;
    ram_cell[     677] = 32'h0;  // 32'hec0a6219;
    ram_cell[     678] = 32'h0;  // 32'h445d31dc;
    ram_cell[     679] = 32'h0;  // 32'ha7f9e83b;
    ram_cell[     680] = 32'h0;  // 32'h83e36b7a;
    ram_cell[     681] = 32'h0;  // 32'h6d10aa63;
    ram_cell[     682] = 32'h0;  // 32'h4e174009;
    ram_cell[     683] = 32'h0;  // 32'hc9746e49;
    ram_cell[     684] = 32'h0;  // 32'hf82a056a;
    ram_cell[     685] = 32'h0;  // 32'hf0f00015;
    ram_cell[     686] = 32'h0;  // 32'hd7f56f5f;
    ram_cell[     687] = 32'h0;  // 32'h42fba786;
    ram_cell[     688] = 32'h0;  // 32'h6debf81f;
    ram_cell[     689] = 32'h0;  // 32'hdfae8dd8;
    ram_cell[     690] = 32'h0;  // 32'h82530fa2;
    ram_cell[     691] = 32'h0;  // 32'he2d38b5d;
    ram_cell[     692] = 32'h0;  // 32'hebf3ffc9;
    ram_cell[     693] = 32'h0;  // 32'hd2cf5d68;
    ram_cell[     694] = 32'h0;  // 32'he72d98a8;
    ram_cell[     695] = 32'h0;  // 32'hc493457c;
    ram_cell[     696] = 32'h0;  // 32'h892ba896;
    ram_cell[     697] = 32'h0;  // 32'h0dcdc6f0;
    ram_cell[     698] = 32'h0;  // 32'h769656a7;
    ram_cell[     699] = 32'h0;  // 32'hacd3ec15;
    ram_cell[     700] = 32'h0;  // 32'hd8b31bbe;
    ram_cell[     701] = 32'h0;  // 32'ha34ec475;
    ram_cell[     702] = 32'h0;  // 32'h0ca3fc97;
    ram_cell[     703] = 32'h0;  // 32'hd164f714;
    ram_cell[     704] = 32'h0;  // 32'h775fc7d0;
    ram_cell[     705] = 32'h0;  // 32'he9648fb4;
    ram_cell[     706] = 32'h0;  // 32'hd6a4f2af;
    ram_cell[     707] = 32'h0;  // 32'hd963408d;
    ram_cell[     708] = 32'h0;  // 32'h081844fb;
    ram_cell[     709] = 32'h0;  // 32'h42b9cc06;
    ram_cell[     710] = 32'h0;  // 32'hb5dd7b94;
    ram_cell[     711] = 32'h0;  // 32'hbfc1d00c;
    ram_cell[     712] = 32'h0;  // 32'h58932147;
    ram_cell[     713] = 32'h0;  // 32'h1af3175e;
    ram_cell[     714] = 32'h0;  // 32'hbae8767a;
    ram_cell[     715] = 32'h0;  // 32'h182c85c8;
    ram_cell[     716] = 32'h0;  // 32'he6dbfb14;
    ram_cell[     717] = 32'h0;  // 32'h49a68fd6;
    ram_cell[     718] = 32'h0;  // 32'hf593ecee;
    ram_cell[     719] = 32'h0;  // 32'h2bb494eb;
    ram_cell[     720] = 32'h0;  // 32'hcff9643a;
    ram_cell[     721] = 32'h0;  // 32'hcd679e17;
    ram_cell[     722] = 32'h0;  // 32'hea9c3fa8;
    ram_cell[     723] = 32'h0;  // 32'h48e3a6ba;
    ram_cell[     724] = 32'h0;  // 32'hccd83738;
    ram_cell[     725] = 32'h0;  // 32'h977c4152;
    ram_cell[     726] = 32'h0;  // 32'hf32a9b8a;
    ram_cell[     727] = 32'h0;  // 32'h969f96d1;
    ram_cell[     728] = 32'h0;  // 32'h5b84920b;
    ram_cell[     729] = 32'h0;  // 32'hb6a117c8;
    ram_cell[     730] = 32'h0;  // 32'hb4d0040d;
    ram_cell[     731] = 32'h0;  // 32'hce2e5a29;
    ram_cell[     732] = 32'h0;  // 32'h90348ff1;
    ram_cell[     733] = 32'h0;  // 32'h3840e3b0;
    ram_cell[     734] = 32'h0;  // 32'h6361cb59;
    ram_cell[     735] = 32'h0;  // 32'h1ad0615a;
    ram_cell[     736] = 32'h0;  // 32'hcd1cc6fc;
    ram_cell[     737] = 32'h0;  // 32'hd2ac67fe;
    ram_cell[     738] = 32'h0;  // 32'hf38877f4;
    ram_cell[     739] = 32'h0;  // 32'hc5bcda86;
    ram_cell[     740] = 32'h0;  // 32'h70767b28;
    ram_cell[     741] = 32'h0;  // 32'h3412dc92;
    ram_cell[     742] = 32'h0;  // 32'h73108934;
    ram_cell[     743] = 32'h0;  // 32'h8ff173db;
    ram_cell[     744] = 32'h0;  // 32'ha65e4d81;
    ram_cell[     745] = 32'h0;  // 32'h9dbfe65d;
    ram_cell[     746] = 32'h0;  // 32'h338ee261;
    ram_cell[     747] = 32'h0;  // 32'ha7daa690;
    ram_cell[     748] = 32'h0;  // 32'h4e11a9c3;
    ram_cell[     749] = 32'h0;  // 32'ha6e3f853;
    ram_cell[     750] = 32'h0;  // 32'h603c8a22;
    ram_cell[     751] = 32'h0;  // 32'h2d04cfea;
    ram_cell[     752] = 32'h0;  // 32'h439bbb26;
    ram_cell[     753] = 32'h0;  // 32'hf876b3ef;
    ram_cell[     754] = 32'h0;  // 32'h72538189;
    ram_cell[     755] = 32'h0;  // 32'h9fbb8a8e;
    ram_cell[     756] = 32'h0;  // 32'h75adaeb7;
    ram_cell[     757] = 32'h0;  // 32'h72b63f37;
    ram_cell[     758] = 32'h0;  // 32'h90f68f66;
    ram_cell[     759] = 32'h0;  // 32'hc327f0a6;
    ram_cell[     760] = 32'h0;  // 32'h17d79c53;
    ram_cell[     761] = 32'h0;  // 32'h7315c30b;
    ram_cell[     762] = 32'h0;  // 32'hf9672969;
    ram_cell[     763] = 32'h0;  // 32'h2cdd1d62;
    ram_cell[     764] = 32'h0;  // 32'h86ef05eb;
    ram_cell[     765] = 32'h0;  // 32'hec501802;
    ram_cell[     766] = 32'h0;  // 32'h50c0cd4d;
    ram_cell[     767] = 32'h0;  // 32'hfc42f0ae;
    ram_cell[     768] = 32'h0;  // 32'h951c6cba;
    ram_cell[     769] = 32'h0;  // 32'h397f8ed2;
    ram_cell[     770] = 32'h0;  // 32'h5b802955;
    ram_cell[     771] = 32'h0;  // 32'h90962327;
    ram_cell[     772] = 32'h0;  // 32'h53d59b54;
    ram_cell[     773] = 32'h0;  // 32'h2d7129f1;
    ram_cell[     774] = 32'h0;  // 32'h20f39a17;
    ram_cell[     775] = 32'h0;  // 32'h86fe3f61;
    ram_cell[     776] = 32'h0;  // 32'hba337c5c;
    ram_cell[     777] = 32'h0;  // 32'h786aab1f;
    ram_cell[     778] = 32'h0;  // 32'h708b98f4;
    ram_cell[     779] = 32'h0;  // 32'h6199cad7;
    ram_cell[     780] = 32'h0;  // 32'hf402420e;
    ram_cell[     781] = 32'h0;  // 32'h7e10cbb5;
    ram_cell[     782] = 32'h0;  // 32'h5815c60f;
    ram_cell[     783] = 32'h0;  // 32'hcfe304cd;
    ram_cell[     784] = 32'h0;  // 32'h42cf637d;
    ram_cell[     785] = 32'h0;  // 32'heb002354;
    ram_cell[     786] = 32'h0;  // 32'h09f52a49;
    ram_cell[     787] = 32'h0;  // 32'h2f47deb0;
    ram_cell[     788] = 32'h0;  // 32'h8597e564;
    ram_cell[     789] = 32'h0;  // 32'hbb1efc2c;
    ram_cell[     790] = 32'h0;  // 32'hfabedff2;
    ram_cell[     791] = 32'h0;  // 32'hc8989b42;
    ram_cell[     792] = 32'h0;  // 32'h7f4c773b;
    ram_cell[     793] = 32'h0;  // 32'he3f2ae5f;
    ram_cell[     794] = 32'h0;  // 32'h22f8e112;
    ram_cell[     795] = 32'h0;  // 32'h8329468b;
    ram_cell[     796] = 32'h0;  // 32'h87b1eed0;
    ram_cell[     797] = 32'h0;  // 32'h9f93ab05;
    ram_cell[     798] = 32'h0;  // 32'h2be25744;
    ram_cell[     799] = 32'h0;  // 32'h3730bb55;
    ram_cell[     800] = 32'h0;  // 32'h08de0795;
    ram_cell[     801] = 32'h0;  // 32'hae9daa66;
    ram_cell[     802] = 32'h0;  // 32'h658c343c;
    ram_cell[     803] = 32'h0;  // 32'hc9b18793;
    ram_cell[     804] = 32'h0;  // 32'h6e89f00c;
    ram_cell[     805] = 32'h0;  // 32'h8fcbe7e9;
    ram_cell[     806] = 32'h0;  // 32'hd0ee0dc9;
    ram_cell[     807] = 32'h0;  // 32'h91195aea;
    ram_cell[     808] = 32'h0;  // 32'h50ee7da4;
    ram_cell[     809] = 32'h0;  // 32'h87402ed1;
    ram_cell[     810] = 32'h0;  // 32'h9391079d;
    ram_cell[     811] = 32'h0;  // 32'h62742e30;
    ram_cell[     812] = 32'h0;  // 32'hdd56acda;
    ram_cell[     813] = 32'h0;  // 32'h3bb0b2f8;
    ram_cell[     814] = 32'h0;  // 32'h046f5bbe;
    ram_cell[     815] = 32'h0;  // 32'hd8763019;
    ram_cell[     816] = 32'h0;  // 32'hdc3a65c7;
    ram_cell[     817] = 32'h0;  // 32'h39e93ed9;
    ram_cell[     818] = 32'h0;  // 32'hd048cfcb;
    ram_cell[     819] = 32'h0;  // 32'h3f50fd3a;
    ram_cell[     820] = 32'h0;  // 32'h1b93a622;
    ram_cell[     821] = 32'h0;  // 32'h7ffbeb5d;
    ram_cell[     822] = 32'h0;  // 32'hd34640cc;
    ram_cell[     823] = 32'h0;  // 32'hcc043eb0;
    ram_cell[     824] = 32'h0;  // 32'h81575c07;
    ram_cell[     825] = 32'h0;  // 32'h3a384f4c;
    ram_cell[     826] = 32'h0;  // 32'hf7749f6b;
    ram_cell[     827] = 32'h0;  // 32'h26291936;
    ram_cell[     828] = 32'h0;  // 32'h28db992b;
    ram_cell[     829] = 32'h0;  // 32'h9e355409;
    ram_cell[     830] = 32'h0;  // 32'he74e7aba;
    ram_cell[     831] = 32'h0;  // 32'h24b5f656;
    ram_cell[     832] = 32'h0;  // 32'he8cca287;
    ram_cell[     833] = 32'h0;  // 32'h56fe196f;
    ram_cell[     834] = 32'h0;  // 32'h6e98ec8f;
    ram_cell[     835] = 32'h0;  // 32'h9ee6a166;
    ram_cell[     836] = 32'h0;  // 32'h5a61c2b6;
    ram_cell[     837] = 32'h0;  // 32'h938a7aad;
    ram_cell[     838] = 32'h0;  // 32'h556dec49;
    ram_cell[     839] = 32'h0;  // 32'hd0e345b9;
    ram_cell[     840] = 32'h0;  // 32'hbfd1bac0;
    ram_cell[     841] = 32'h0;  // 32'h295f56fd;
    ram_cell[     842] = 32'h0;  // 32'ha6165fc9;
    ram_cell[     843] = 32'h0;  // 32'h087de5de;
    ram_cell[     844] = 32'h0;  // 32'h6158ad0d;
    ram_cell[     845] = 32'h0;  // 32'h19c6f5b1;
    ram_cell[     846] = 32'h0;  // 32'h9cca3c4b;
    ram_cell[     847] = 32'h0;  // 32'h5f02490d;
    ram_cell[     848] = 32'h0;  // 32'h98246d03;
    ram_cell[     849] = 32'h0;  // 32'h8967f510;
    ram_cell[     850] = 32'h0;  // 32'haa92d60c;
    ram_cell[     851] = 32'h0;  // 32'h7161de9e;
    ram_cell[     852] = 32'h0;  // 32'h300d0160;
    ram_cell[     853] = 32'h0;  // 32'hc88242d4;
    ram_cell[     854] = 32'h0;  // 32'hb7811cfe;
    ram_cell[     855] = 32'h0;  // 32'h0171ab82;
    ram_cell[     856] = 32'h0;  // 32'h96644a4e;
    ram_cell[     857] = 32'h0;  // 32'hba224ec3;
    ram_cell[     858] = 32'h0;  // 32'h120d25c5;
    ram_cell[     859] = 32'h0;  // 32'h1e32c99d;
    ram_cell[     860] = 32'h0;  // 32'h099f6414;
    ram_cell[     861] = 32'h0;  // 32'h9aecc18d;
    ram_cell[     862] = 32'h0;  // 32'h2b7c7246;
    ram_cell[     863] = 32'h0;  // 32'he011df09;
    ram_cell[     864] = 32'h0;  // 32'h91b84231;
    ram_cell[     865] = 32'h0;  // 32'h85fc07d0;
    ram_cell[     866] = 32'h0;  // 32'h435ccbce;
    ram_cell[     867] = 32'h0;  // 32'ha0a92bfe;
    ram_cell[     868] = 32'h0;  // 32'h0da83915;
    ram_cell[     869] = 32'h0;  // 32'h819fa720;
    ram_cell[     870] = 32'h0;  // 32'hb723200b;
    ram_cell[     871] = 32'h0;  // 32'h56d0c423;
    ram_cell[     872] = 32'h0;  // 32'h36b51a7e;
    ram_cell[     873] = 32'h0;  // 32'h9b71d080;
    ram_cell[     874] = 32'h0;  // 32'h606d0c06;
    ram_cell[     875] = 32'h0;  // 32'hf13d38d2;
    ram_cell[     876] = 32'h0;  // 32'h28edb79d;
    ram_cell[     877] = 32'h0;  // 32'h152d1916;
    ram_cell[     878] = 32'h0;  // 32'h7b3b2191;
    ram_cell[     879] = 32'h0;  // 32'he1ad13e8;
    ram_cell[     880] = 32'h0;  // 32'hd30941fc;
    ram_cell[     881] = 32'h0;  // 32'h313de7a1;
    ram_cell[     882] = 32'h0;  // 32'ha9f1edfa;
    ram_cell[     883] = 32'h0;  // 32'h3957f0c7;
    ram_cell[     884] = 32'h0;  // 32'hbe55f025;
    ram_cell[     885] = 32'h0;  // 32'h0cdce44f;
    ram_cell[     886] = 32'h0;  // 32'h759bea57;
    ram_cell[     887] = 32'h0;  // 32'ha39cc271;
    ram_cell[     888] = 32'h0;  // 32'h4ebea84c;
    ram_cell[     889] = 32'h0;  // 32'hbad325ba;
    ram_cell[     890] = 32'h0;  // 32'h12a065e7;
    ram_cell[     891] = 32'h0;  // 32'h16e5c417;
    ram_cell[     892] = 32'h0;  // 32'h77f6e907;
    ram_cell[     893] = 32'h0;  // 32'h8b4d9917;
    ram_cell[     894] = 32'h0;  // 32'h58c7b91d;
    ram_cell[     895] = 32'h0;  // 32'h6bd843d5;
    ram_cell[     896] = 32'h0;  // 32'hd1cc5424;
    ram_cell[     897] = 32'h0;  // 32'h06a75cec;
    ram_cell[     898] = 32'h0;  // 32'h403b208b;
    ram_cell[     899] = 32'h0;  // 32'h4f012c53;
    ram_cell[     900] = 32'h0;  // 32'h4bf46c74;
    ram_cell[     901] = 32'h0;  // 32'h1390a3a5;
    ram_cell[     902] = 32'h0;  // 32'h4faf2e10;
    ram_cell[     903] = 32'h0;  // 32'ha9b16daa;
    ram_cell[     904] = 32'h0;  // 32'h772aa31b;
    ram_cell[     905] = 32'h0;  // 32'h01467f4f;
    ram_cell[     906] = 32'h0;  // 32'hdd3228e2;
    ram_cell[     907] = 32'h0;  // 32'h5cea9c3d;
    ram_cell[     908] = 32'h0;  // 32'hefac61aa;
    ram_cell[     909] = 32'h0;  // 32'h9d249f1a;
    ram_cell[     910] = 32'h0;  // 32'h2b73e826;
    ram_cell[     911] = 32'h0;  // 32'hf552f4d6;
    ram_cell[     912] = 32'h0;  // 32'h4cde6c2a;
    ram_cell[     913] = 32'h0;  // 32'h2d10966c;
    ram_cell[     914] = 32'h0;  // 32'h49f04d30;
    ram_cell[     915] = 32'h0;  // 32'h950ee305;
    ram_cell[     916] = 32'h0;  // 32'h92e1025e;
    ram_cell[     917] = 32'h0;  // 32'he71f4af1;
    ram_cell[     918] = 32'h0;  // 32'h63d9cf7c;
    ram_cell[     919] = 32'h0;  // 32'h99cdedc8;
    ram_cell[     920] = 32'h0;  // 32'hc36bf7c1;
    ram_cell[     921] = 32'h0;  // 32'h7f540c3c;
    ram_cell[     922] = 32'h0;  // 32'h2d96bb78;
    ram_cell[     923] = 32'h0;  // 32'h3f9629f2;
    ram_cell[     924] = 32'h0;  // 32'h0644bea4;
    ram_cell[     925] = 32'h0;  // 32'h11d8e72d;
    ram_cell[     926] = 32'h0;  // 32'hf6d9de7e;
    ram_cell[     927] = 32'h0;  // 32'hde112b2a;
    ram_cell[     928] = 32'h0;  // 32'ha5825a68;
    ram_cell[     929] = 32'h0;  // 32'h4b749c46;
    ram_cell[     930] = 32'h0;  // 32'hbdeb2a85;
    ram_cell[     931] = 32'h0;  // 32'hd731842d;
    ram_cell[     932] = 32'h0;  // 32'h875e2d57;
    ram_cell[     933] = 32'h0;  // 32'h9bfe60ec;
    ram_cell[     934] = 32'h0;  // 32'hd680e9ea;
    ram_cell[     935] = 32'h0;  // 32'hd246e4a6;
    ram_cell[     936] = 32'h0;  // 32'hb638ff14;
    ram_cell[     937] = 32'h0;  // 32'he656a4b6;
    ram_cell[     938] = 32'h0;  // 32'h2d2c9c05;
    ram_cell[     939] = 32'h0;  // 32'h4156d49d;
    ram_cell[     940] = 32'h0;  // 32'hf1067516;
    ram_cell[     941] = 32'h0;  // 32'h567a43cc;
    ram_cell[     942] = 32'h0;  // 32'h46eb22df;
    ram_cell[     943] = 32'h0;  // 32'h312bc6f4;
    ram_cell[     944] = 32'h0;  // 32'h527b26be;
    ram_cell[     945] = 32'h0;  // 32'h7aa4b69f;
    ram_cell[     946] = 32'h0;  // 32'h1c54934e;
    ram_cell[     947] = 32'h0;  // 32'hb43409e9;
    ram_cell[     948] = 32'h0;  // 32'h6bb8af3a;
    ram_cell[     949] = 32'h0;  // 32'h012057fb;
    ram_cell[     950] = 32'h0;  // 32'hd1e6032f;
    ram_cell[     951] = 32'h0;  // 32'hebd0bace;
    ram_cell[     952] = 32'h0;  // 32'hf764fadb;
    ram_cell[     953] = 32'h0;  // 32'hde60c2f8;
    ram_cell[     954] = 32'h0;  // 32'hff6b1aab;
    ram_cell[     955] = 32'h0;  // 32'hf8a01a58;
    ram_cell[     956] = 32'h0;  // 32'hb5e0ae42;
    ram_cell[     957] = 32'h0;  // 32'hde4f541a;
    ram_cell[     958] = 32'h0;  // 32'hb8eb9b35;
    ram_cell[     959] = 32'h0;  // 32'hcb4ca317;
    ram_cell[     960] = 32'h0;  // 32'h091179b4;
    ram_cell[     961] = 32'h0;  // 32'ha942cf57;
    ram_cell[     962] = 32'h0;  // 32'hcff8a948;
    ram_cell[     963] = 32'h0;  // 32'h5c4efb60;
    ram_cell[     964] = 32'h0;  // 32'h96cf0377;
    ram_cell[     965] = 32'h0;  // 32'h94673d3b;
    ram_cell[     966] = 32'h0;  // 32'h5a04d62a;
    ram_cell[     967] = 32'h0;  // 32'h93dc6901;
    ram_cell[     968] = 32'h0;  // 32'he7449e27;
    ram_cell[     969] = 32'h0;  // 32'heceb5e6a;
    ram_cell[     970] = 32'h0;  // 32'h54c7b71d;
    ram_cell[     971] = 32'h0;  // 32'h32634ed0;
    ram_cell[     972] = 32'h0;  // 32'h4b1ab702;
    ram_cell[     973] = 32'h0;  // 32'h60c94dd2;
    ram_cell[     974] = 32'h0;  // 32'h90b3cb51;
    ram_cell[     975] = 32'h0;  // 32'h22e27422;
    ram_cell[     976] = 32'h0;  // 32'h067979e2;
    ram_cell[     977] = 32'h0;  // 32'h9837f4a2;
    ram_cell[     978] = 32'h0;  // 32'he00f2a37;
    ram_cell[     979] = 32'h0;  // 32'he445e381;
    ram_cell[     980] = 32'h0;  // 32'h9c3d61f0;
    ram_cell[     981] = 32'h0;  // 32'h38a1e442;
    ram_cell[     982] = 32'h0;  // 32'h4b9cfbf0;
    ram_cell[     983] = 32'h0;  // 32'h4ba1314c;
    ram_cell[     984] = 32'h0;  // 32'h26d37d4d;
    ram_cell[     985] = 32'h0;  // 32'hb7ffcfe0;
    ram_cell[     986] = 32'h0;  // 32'h0e9bb437;
    ram_cell[     987] = 32'h0;  // 32'h42a38b75;
    ram_cell[     988] = 32'h0;  // 32'hcf7450f9;
    ram_cell[     989] = 32'h0;  // 32'hc2ac01d1;
    ram_cell[     990] = 32'h0;  // 32'h034fdc62;
    ram_cell[     991] = 32'h0;  // 32'h807e9d14;
    ram_cell[     992] = 32'h0;  // 32'hc7bcbac6;
    ram_cell[     993] = 32'h0;  // 32'he18a4117;
    ram_cell[     994] = 32'h0;  // 32'hece635f7;
    ram_cell[     995] = 32'h0;  // 32'hcd551f10;
    ram_cell[     996] = 32'h0;  // 32'h2df404db;
    ram_cell[     997] = 32'h0;  // 32'hd149574f;
    ram_cell[     998] = 32'h0;  // 32'h6c1d7102;
    ram_cell[     999] = 32'h0;  // 32'ha62fae62;
    ram_cell[    1000] = 32'h0;  // 32'h9446a0c3;
    ram_cell[    1001] = 32'h0;  // 32'h87585f46;
    ram_cell[    1002] = 32'h0;  // 32'h1c63f9c0;
    ram_cell[    1003] = 32'h0;  // 32'h7f34e1d4;
    ram_cell[    1004] = 32'h0;  // 32'hc0a8e971;
    ram_cell[    1005] = 32'h0;  // 32'h859b5eee;
    ram_cell[    1006] = 32'h0;  // 32'hdf0299fb;
    ram_cell[    1007] = 32'h0;  // 32'h1a4e6531;
    ram_cell[    1008] = 32'h0;  // 32'h9c7cd166;
    ram_cell[    1009] = 32'h0;  // 32'h86a3f4bd;
    ram_cell[    1010] = 32'h0;  // 32'h79d3ccd8;
    ram_cell[    1011] = 32'h0;  // 32'h96f127bd;
    ram_cell[    1012] = 32'h0;  // 32'he9eed389;
    ram_cell[    1013] = 32'h0;  // 32'h9bf33ffd;
    ram_cell[    1014] = 32'h0;  // 32'hf5081800;
    ram_cell[    1015] = 32'h0;  // 32'h0e484f2e;
    ram_cell[    1016] = 32'h0;  // 32'h1a539aa8;
    ram_cell[    1017] = 32'h0;  // 32'h800a5f11;
    ram_cell[    1018] = 32'h0;  // 32'h80ec29d1;
    ram_cell[    1019] = 32'h0;  // 32'h8f572012;
    ram_cell[    1020] = 32'h0;  // 32'h0b85e1de;
    ram_cell[    1021] = 32'h0;  // 32'h76ce46cf;
    ram_cell[    1022] = 32'h0;  // 32'h6e6a2a4f;
    ram_cell[    1023] = 32'h0;  // 32'h8541f91a;
    // src matrix A
    ram_cell[    1024] = 32'hbee8d368;
    ram_cell[    1025] = 32'he66f569c;
    ram_cell[    1026] = 32'h2074437b;
    ram_cell[    1027] = 32'h54d1db17;
    ram_cell[    1028] = 32'h18b05ce8;
    ram_cell[    1029] = 32'hf533f3a8;
    ram_cell[    1030] = 32'haf567915;
    ram_cell[    1031] = 32'h9cc1da9b;
    ram_cell[    1032] = 32'h8d1dcbad;
    ram_cell[    1033] = 32'h46120669;
    ram_cell[    1034] = 32'h7e7310dd;
    ram_cell[    1035] = 32'h28384869;
    ram_cell[    1036] = 32'he79eaffc;
    ram_cell[    1037] = 32'hf0c603e7;
    ram_cell[    1038] = 32'h84b45b0c;
    ram_cell[    1039] = 32'h9b26f238;
    ram_cell[    1040] = 32'hd75d7267;
    ram_cell[    1041] = 32'ha5ca018a;
    ram_cell[    1042] = 32'h8a0d0e3d;
    ram_cell[    1043] = 32'h25a453b4;
    ram_cell[    1044] = 32'h60c534bc;
    ram_cell[    1045] = 32'h162348dd;
    ram_cell[    1046] = 32'hb40fc6e9;
    ram_cell[    1047] = 32'hfa18c51f;
    ram_cell[    1048] = 32'hd81a450c;
    ram_cell[    1049] = 32'hde313028;
    ram_cell[    1050] = 32'hefe0d327;
    ram_cell[    1051] = 32'hf743bba7;
    ram_cell[    1052] = 32'hd3699e82;
    ram_cell[    1053] = 32'hb306ee77;
    ram_cell[    1054] = 32'h425bc2cf;
    ram_cell[    1055] = 32'h9b7ca2dc;
    ram_cell[    1056] = 32'h2a061609;
    ram_cell[    1057] = 32'h72c5a2a9;
    ram_cell[    1058] = 32'h4a1b495b;
    ram_cell[    1059] = 32'ha2b89520;
    ram_cell[    1060] = 32'h6e302d7f;
    ram_cell[    1061] = 32'he2d95684;
    ram_cell[    1062] = 32'hc49a180f;
    ram_cell[    1063] = 32'h07289384;
    ram_cell[    1064] = 32'h6f305f56;
    ram_cell[    1065] = 32'hcf250733;
    ram_cell[    1066] = 32'h12c9e33a;
    ram_cell[    1067] = 32'hbe050cce;
    ram_cell[    1068] = 32'h1b02f91c;
    ram_cell[    1069] = 32'hf214d46a;
    ram_cell[    1070] = 32'h559ce023;
    ram_cell[    1071] = 32'ha1efc5e5;
    ram_cell[    1072] = 32'h5271311e;
    ram_cell[    1073] = 32'h2623efea;
    ram_cell[    1074] = 32'hfc538caa;
    ram_cell[    1075] = 32'h4c754fb9;
    ram_cell[    1076] = 32'h9836add0;
    ram_cell[    1077] = 32'h588759cb;
    ram_cell[    1078] = 32'h4bffc078;
    ram_cell[    1079] = 32'hd530ea64;
    ram_cell[    1080] = 32'h30fb0f3d;
    ram_cell[    1081] = 32'h0de71b5d;
    ram_cell[    1082] = 32'h5a5e4c3e;
    ram_cell[    1083] = 32'h4dfeb9c1;
    ram_cell[    1084] = 32'h85e59591;
    ram_cell[    1085] = 32'ha2a7d56c;
    ram_cell[    1086] = 32'h60231094;
    ram_cell[    1087] = 32'h7b40f71d;
    ram_cell[    1088] = 32'ha569d1b1;
    ram_cell[    1089] = 32'h63d7854f;
    ram_cell[    1090] = 32'hfc07e046;
    ram_cell[    1091] = 32'hfe9be7b1;
    ram_cell[    1092] = 32'h74db1d9a;
    ram_cell[    1093] = 32'haf9e3071;
    ram_cell[    1094] = 32'h0838b87d;
    ram_cell[    1095] = 32'h66a88f3f;
    ram_cell[    1096] = 32'hf3d46067;
    ram_cell[    1097] = 32'h25bb643e;
    ram_cell[    1098] = 32'h290510c9;
    ram_cell[    1099] = 32'h6c8e7d29;
    ram_cell[    1100] = 32'h1fcb5889;
    ram_cell[    1101] = 32'hc7eb65f2;
    ram_cell[    1102] = 32'hccee22c2;
    ram_cell[    1103] = 32'h28abe882;
    ram_cell[    1104] = 32'hfccf35de;
    ram_cell[    1105] = 32'hcf9b2a89;
    ram_cell[    1106] = 32'hc6ca9789;
    ram_cell[    1107] = 32'hbcb85e40;
    ram_cell[    1108] = 32'h0ac4da70;
    ram_cell[    1109] = 32'hee24fcbd;
    ram_cell[    1110] = 32'h9a2ee56d;
    ram_cell[    1111] = 32'hf8f9703c;
    ram_cell[    1112] = 32'h2d2b0241;
    ram_cell[    1113] = 32'hb599c2f7;
    ram_cell[    1114] = 32'hd0ac4aea;
    ram_cell[    1115] = 32'h56ad210b;
    ram_cell[    1116] = 32'h24642e24;
    ram_cell[    1117] = 32'hdee29d41;
    ram_cell[    1118] = 32'hc5fc3081;
    ram_cell[    1119] = 32'h4df7ee2a;
    ram_cell[    1120] = 32'h9ac4949e;
    ram_cell[    1121] = 32'hac834808;
    ram_cell[    1122] = 32'h61a4cec6;
    ram_cell[    1123] = 32'h6dd94839;
    ram_cell[    1124] = 32'h9e49f523;
    ram_cell[    1125] = 32'h902e1236;
    ram_cell[    1126] = 32'h67f557ed;
    ram_cell[    1127] = 32'had90dc82;
    ram_cell[    1128] = 32'h4c4a08f6;
    ram_cell[    1129] = 32'ha31e19fe;
    ram_cell[    1130] = 32'h8b6c6854;
    ram_cell[    1131] = 32'haf13753b;
    ram_cell[    1132] = 32'h9b1a7938;
    ram_cell[    1133] = 32'ha60fd19b;
    ram_cell[    1134] = 32'h961bcbb9;
    ram_cell[    1135] = 32'h0aca2654;
    ram_cell[    1136] = 32'hec8641c2;
    ram_cell[    1137] = 32'hbaf7f680;
    ram_cell[    1138] = 32'hba0e6e4f;
    ram_cell[    1139] = 32'h7e9ae4c7;
    ram_cell[    1140] = 32'he92d255d;
    ram_cell[    1141] = 32'hc2fecd61;
    ram_cell[    1142] = 32'h3c1ca0f4;
    ram_cell[    1143] = 32'h3238fbc1;
    ram_cell[    1144] = 32'h05ba584a;
    ram_cell[    1145] = 32'h49a1615b;
    ram_cell[    1146] = 32'h1dfbc294;
    ram_cell[    1147] = 32'h5cd7fb77;
    ram_cell[    1148] = 32'h9498f538;
    ram_cell[    1149] = 32'ha032968c;
    ram_cell[    1150] = 32'h039a947f;
    ram_cell[    1151] = 32'h0110bdd7;
    ram_cell[    1152] = 32'h1b48f219;
    ram_cell[    1153] = 32'h66f707b8;
    ram_cell[    1154] = 32'h5608d834;
    ram_cell[    1155] = 32'h287e5b41;
    ram_cell[    1156] = 32'h018384c7;
    ram_cell[    1157] = 32'hf3cec7a5;
    ram_cell[    1158] = 32'hb76c7afd;
    ram_cell[    1159] = 32'h67753420;
    ram_cell[    1160] = 32'h5812b0b1;
    ram_cell[    1161] = 32'h2b7054cc;
    ram_cell[    1162] = 32'hf66fc0b1;
    ram_cell[    1163] = 32'hf84da533;
    ram_cell[    1164] = 32'h732d38c2;
    ram_cell[    1165] = 32'hf59c8e71;
    ram_cell[    1166] = 32'h84728239;
    ram_cell[    1167] = 32'hd5b672e2;
    ram_cell[    1168] = 32'h662c05fa;
    ram_cell[    1169] = 32'h0eb03ece;
    ram_cell[    1170] = 32'hd659c23d;
    ram_cell[    1171] = 32'hdbdcb435;
    ram_cell[    1172] = 32'hd254372f;
    ram_cell[    1173] = 32'h0e5cd41a;
    ram_cell[    1174] = 32'h023b50e6;
    ram_cell[    1175] = 32'hd9b4be15;
    ram_cell[    1176] = 32'h6d9cb3b0;
    ram_cell[    1177] = 32'h58b295df;
    ram_cell[    1178] = 32'hc1efbf29;
    ram_cell[    1179] = 32'h3db38b29;
    ram_cell[    1180] = 32'hd4ee525b;
    ram_cell[    1181] = 32'ha71cc215;
    ram_cell[    1182] = 32'h019dd985;
    ram_cell[    1183] = 32'h6a9c3146;
    ram_cell[    1184] = 32'h6a32bbd6;
    ram_cell[    1185] = 32'h1740a0dc;
    ram_cell[    1186] = 32'h9c57be88;
    ram_cell[    1187] = 32'h9503d0c9;
    ram_cell[    1188] = 32'h5b99d051;
    ram_cell[    1189] = 32'h189ff10e;
    ram_cell[    1190] = 32'h32d55da5;
    ram_cell[    1191] = 32'hcb8d8f55;
    ram_cell[    1192] = 32'h9dde1372;
    ram_cell[    1193] = 32'h989c5d8b;
    ram_cell[    1194] = 32'h2605e4bd;
    ram_cell[    1195] = 32'h7052f279;
    ram_cell[    1196] = 32'h34c2b6ed;
    ram_cell[    1197] = 32'h56ec5f08;
    ram_cell[    1198] = 32'hde7d5d32;
    ram_cell[    1199] = 32'h020c8123;
    ram_cell[    1200] = 32'h9f4d961e;
    ram_cell[    1201] = 32'h40a781fe;
    ram_cell[    1202] = 32'h6df481fa;
    ram_cell[    1203] = 32'he8dc5e6e;
    ram_cell[    1204] = 32'hde809812;
    ram_cell[    1205] = 32'hf9e8c7f2;
    ram_cell[    1206] = 32'h7145ff13;
    ram_cell[    1207] = 32'h734276af;
    ram_cell[    1208] = 32'h8cdca45b;
    ram_cell[    1209] = 32'he76db252;
    ram_cell[    1210] = 32'hc438f7b6;
    ram_cell[    1211] = 32'h2643c13e;
    ram_cell[    1212] = 32'h310e7826;
    ram_cell[    1213] = 32'hefb7240b;
    ram_cell[    1214] = 32'h29fa6fab;
    ram_cell[    1215] = 32'hc47eedc5;
    ram_cell[    1216] = 32'hf5a766d4;
    ram_cell[    1217] = 32'h9c87777f;
    ram_cell[    1218] = 32'ha4807d32;
    ram_cell[    1219] = 32'h7d4dc191;
    ram_cell[    1220] = 32'h122e692c;
    ram_cell[    1221] = 32'hda16a1b3;
    ram_cell[    1222] = 32'hc2015898;
    ram_cell[    1223] = 32'hdca4dcbd;
    ram_cell[    1224] = 32'h0432e155;
    ram_cell[    1225] = 32'h558a8c8e;
    ram_cell[    1226] = 32'hc3daf2a1;
    ram_cell[    1227] = 32'hac6f68a3;
    ram_cell[    1228] = 32'h0c964f3d;
    ram_cell[    1229] = 32'h928f4e21;
    ram_cell[    1230] = 32'h700e2055;
    ram_cell[    1231] = 32'he759ad33;
    ram_cell[    1232] = 32'h5dc5b076;
    ram_cell[    1233] = 32'hb05c2cd3;
    ram_cell[    1234] = 32'hff9b02f6;
    ram_cell[    1235] = 32'h3a840e70;
    ram_cell[    1236] = 32'h4f406ce7;
    ram_cell[    1237] = 32'h5b19ef0b;
    ram_cell[    1238] = 32'h4070bced;
    ram_cell[    1239] = 32'h51a04cb0;
    ram_cell[    1240] = 32'hb9ea16a2;
    ram_cell[    1241] = 32'h0bda8e7b;
    ram_cell[    1242] = 32'h5495c634;
    ram_cell[    1243] = 32'h7474e1d7;
    ram_cell[    1244] = 32'h37f29e14;
    ram_cell[    1245] = 32'h3bb576c2;
    ram_cell[    1246] = 32'hc1b83e6c;
    ram_cell[    1247] = 32'h5bcb9df1;
    ram_cell[    1248] = 32'h8549dc1c;
    ram_cell[    1249] = 32'h1ddc8023;
    ram_cell[    1250] = 32'h6d04e95c;
    ram_cell[    1251] = 32'h2eb764cb;
    ram_cell[    1252] = 32'h9e59b1a8;
    ram_cell[    1253] = 32'hc5cba65b;
    ram_cell[    1254] = 32'h5e7b2a37;
    ram_cell[    1255] = 32'hce87f367;
    ram_cell[    1256] = 32'h05a543ed;
    ram_cell[    1257] = 32'ha2c98a80;
    ram_cell[    1258] = 32'h098311c9;
    ram_cell[    1259] = 32'h1b29dc2b;
    ram_cell[    1260] = 32'h74dd4e3c;
    ram_cell[    1261] = 32'h99c8d6ff;
    ram_cell[    1262] = 32'he266b410;
    ram_cell[    1263] = 32'h00f91b26;
    ram_cell[    1264] = 32'he840dda2;
    ram_cell[    1265] = 32'h37d7d5c9;
    ram_cell[    1266] = 32'hc17d442d;
    ram_cell[    1267] = 32'h8fd3ba5d;
    ram_cell[    1268] = 32'hca0f293d;
    ram_cell[    1269] = 32'h72669e79;
    ram_cell[    1270] = 32'h2fac9b18;
    ram_cell[    1271] = 32'h89247f5d;
    ram_cell[    1272] = 32'hbd5cdbf7;
    ram_cell[    1273] = 32'h4f5f4d76;
    ram_cell[    1274] = 32'h1a5cd8ef;
    ram_cell[    1275] = 32'hedcb9299;
    ram_cell[    1276] = 32'h21033c7b;
    ram_cell[    1277] = 32'ha8875edb;
    ram_cell[    1278] = 32'h57c451de;
    ram_cell[    1279] = 32'h560939cd;
    ram_cell[    1280] = 32'h53d95a63;
    ram_cell[    1281] = 32'h5cea9498;
    ram_cell[    1282] = 32'h5be35cb7;
    ram_cell[    1283] = 32'h79924712;
    ram_cell[    1284] = 32'h3d58e963;
    ram_cell[    1285] = 32'h26db3b40;
    ram_cell[    1286] = 32'hd2953d09;
    ram_cell[    1287] = 32'h60c821b2;
    ram_cell[    1288] = 32'ha29b5e4b;
    ram_cell[    1289] = 32'ha7a4e739;
    ram_cell[    1290] = 32'h1a229c8c;
    ram_cell[    1291] = 32'hbcbcc861;
    ram_cell[    1292] = 32'hb1f4f677;
    ram_cell[    1293] = 32'h4ba1c30f;
    ram_cell[    1294] = 32'h2ab074dc;
    ram_cell[    1295] = 32'h9db88852;
    ram_cell[    1296] = 32'hc5a5cadc;
    ram_cell[    1297] = 32'h6c47ac30;
    ram_cell[    1298] = 32'h0d448fca;
    ram_cell[    1299] = 32'h0d0a345e;
    ram_cell[    1300] = 32'h5b5541d3;
    ram_cell[    1301] = 32'h357c2589;
    ram_cell[    1302] = 32'hbd19b260;
    ram_cell[    1303] = 32'h27c11d73;
    ram_cell[    1304] = 32'hb56aaa1f;
    ram_cell[    1305] = 32'h9d1a9529;
    ram_cell[    1306] = 32'hfe26e1e6;
    ram_cell[    1307] = 32'hb3034b39;
    ram_cell[    1308] = 32'heb5ca979;
    ram_cell[    1309] = 32'h260d28fb;
    ram_cell[    1310] = 32'h824eaab8;
    ram_cell[    1311] = 32'h5ffacd23;
    ram_cell[    1312] = 32'h6100f86f;
    ram_cell[    1313] = 32'h9df3fe67;
    ram_cell[    1314] = 32'h47cba8f4;
    ram_cell[    1315] = 32'h032df9d8;
    ram_cell[    1316] = 32'h494de145;
    ram_cell[    1317] = 32'hf6abd005;
    ram_cell[    1318] = 32'hae73377f;
    ram_cell[    1319] = 32'h2ed2538b;
    ram_cell[    1320] = 32'h818ce903;
    ram_cell[    1321] = 32'h26751b82;
    ram_cell[    1322] = 32'h4cc1992e;
    ram_cell[    1323] = 32'hc984fcc0;
    ram_cell[    1324] = 32'h27cc2b67;
    ram_cell[    1325] = 32'h1155033a;
    ram_cell[    1326] = 32'hf4a413b5;
    ram_cell[    1327] = 32'hac8c8f2e;
    ram_cell[    1328] = 32'h961aceee;
    ram_cell[    1329] = 32'h4100f751;
    ram_cell[    1330] = 32'hce35c6d5;
    ram_cell[    1331] = 32'hf45380fe;
    ram_cell[    1332] = 32'h9b5a0d6b;
    ram_cell[    1333] = 32'h2dce6d25;
    ram_cell[    1334] = 32'hdeb0c086;
    ram_cell[    1335] = 32'h69efc3f3;
    ram_cell[    1336] = 32'he979e19e;
    ram_cell[    1337] = 32'h5d1b8dcf;
    ram_cell[    1338] = 32'hac8d0f59;
    ram_cell[    1339] = 32'h34ff3285;
    ram_cell[    1340] = 32'hd6ac00d2;
    ram_cell[    1341] = 32'h7b3ad6d5;
    ram_cell[    1342] = 32'h5f4d2ce2;
    ram_cell[    1343] = 32'h78243c8b;
    ram_cell[    1344] = 32'h295d18ac;
    ram_cell[    1345] = 32'h8d826b94;
    ram_cell[    1346] = 32'ha6a5bc9d;
    ram_cell[    1347] = 32'hf3e9c777;
    ram_cell[    1348] = 32'h298c7cf2;
    ram_cell[    1349] = 32'hca998084;
    ram_cell[    1350] = 32'hd53c68a8;
    ram_cell[    1351] = 32'h5070bb65;
    ram_cell[    1352] = 32'h3dd8c937;
    ram_cell[    1353] = 32'hf5ae55f5;
    ram_cell[    1354] = 32'h111d7d7c;
    ram_cell[    1355] = 32'h0a97256c;
    ram_cell[    1356] = 32'h605fcbec;
    ram_cell[    1357] = 32'h40d7145f;
    ram_cell[    1358] = 32'h7430a3ed;
    ram_cell[    1359] = 32'h379c5c2c;
    ram_cell[    1360] = 32'h510611c8;
    ram_cell[    1361] = 32'h17e576c5;
    ram_cell[    1362] = 32'hca3d80f8;
    ram_cell[    1363] = 32'h0fa90093;
    ram_cell[    1364] = 32'h65ccda9c;
    ram_cell[    1365] = 32'hb1976853;
    ram_cell[    1366] = 32'ha0d2e7d3;
    ram_cell[    1367] = 32'h8a1abb16;
    ram_cell[    1368] = 32'h334c7fb2;
    ram_cell[    1369] = 32'he606cdd1;
    ram_cell[    1370] = 32'he2dc694e;
    ram_cell[    1371] = 32'hc00f983b;
    ram_cell[    1372] = 32'ha5272f5d;
    ram_cell[    1373] = 32'h44aaaf7d;
    ram_cell[    1374] = 32'h7b63d3a7;
    ram_cell[    1375] = 32'h0062294c;
    ram_cell[    1376] = 32'ha48c5f27;
    ram_cell[    1377] = 32'h40acba03;
    ram_cell[    1378] = 32'hea1cf260;
    ram_cell[    1379] = 32'h0b65809e;
    ram_cell[    1380] = 32'h7596adff;
    ram_cell[    1381] = 32'hc8510236;
    ram_cell[    1382] = 32'h2e7bfb77;
    ram_cell[    1383] = 32'h68c3744b;
    ram_cell[    1384] = 32'h45b9b012;
    ram_cell[    1385] = 32'h08e1a932;
    ram_cell[    1386] = 32'h06ea1e1c;
    ram_cell[    1387] = 32'h2f1992d4;
    ram_cell[    1388] = 32'ha9cfddf2;
    ram_cell[    1389] = 32'hd9fa2177;
    ram_cell[    1390] = 32'h689fb50f;
    ram_cell[    1391] = 32'hffc87d48;
    ram_cell[    1392] = 32'h5101c5c1;
    ram_cell[    1393] = 32'h735fd0c9;
    ram_cell[    1394] = 32'h0b9fd362;
    ram_cell[    1395] = 32'h667d248b;
    ram_cell[    1396] = 32'hb2417da2;
    ram_cell[    1397] = 32'h5b9b8194;
    ram_cell[    1398] = 32'hacee7e3e;
    ram_cell[    1399] = 32'h34e40d18;
    ram_cell[    1400] = 32'h74f02bc8;
    ram_cell[    1401] = 32'hf2ca4414;
    ram_cell[    1402] = 32'hf996e88b;
    ram_cell[    1403] = 32'he092ede3;
    ram_cell[    1404] = 32'h9ac8bc22;
    ram_cell[    1405] = 32'h118c1717;
    ram_cell[    1406] = 32'hc396156e;
    ram_cell[    1407] = 32'h9aa83fcb;
    ram_cell[    1408] = 32'hdea2d548;
    ram_cell[    1409] = 32'hd7f6d3d4;
    ram_cell[    1410] = 32'h038e167e;
    ram_cell[    1411] = 32'hb3800983;
    ram_cell[    1412] = 32'haf5593d6;
    ram_cell[    1413] = 32'h1ee81344;
    ram_cell[    1414] = 32'hba45295e;
    ram_cell[    1415] = 32'hf05e0a81;
    ram_cell[    1416] = 32'h657c02b3;
    ram_cell[    1417] = 32'h52b14747;
    ram_cell[    1418] = 32'h1520cec9;
    ram_cell[    1419] = 32'hb4d444af;
    ram_cell[    1420] = 32'h1d0d804b;
    ram_cell[    1421] = 32'h9d34bf17;
    ram_cell[    1422] = 32'h3206ac7c;
    ram_cell[    1423] = 32'h9f97058e;
    ram_cell[    1424] = 32'h7e182f1c;
    ram_cell[    1425] = 32'h6a867afc;
    ram_cell[    1426] = 32'hf963b7d0;
    ram_cell[    1427] = 32'h8bb75bd1;
    ram_cell[    1428] = 32'h3b3cad65;
    ram_cell[    1429] = 32'h2143a2c6;
    ram_cell[    1430] = 32'hed8bdeb3;
    ram_cell[    1431] = 32'h055d1033;
    ram_cell[    1432] = 32'h9aed74a7;
    ram_cell[    1433] = 32'h2da10971;
    ram_cell[    1434] = 32'h154660f7;
    ram_cell[    1435] = 32'hbb8ecf6d;
    ram_cell[    1436] = 32'h4f3b10a9;
    ram_cell[    1437] = 32'h75879786;
    ram_cell[    1438] = 32'h8c4542c4;
    ram_cell[    1439] = 32'h20fb3e70;
    ram_cell[    1440] = 32'h8d628ea1;
    ram_cell[    1441] = 32'hf2a40304;
    ram_cell[    1442] = 32'h4440ee3f;
    ram_cell[    1443] = 32'hea49dc72;
    ram_cell[    1444] = 32'h1ff3bf90;
    ram_cell[    1445] = 32'ha1974bd5;
    ram_cell[    1446] = 32'hacb2ef18;
    ram_cell[    1447] = 32'he94fca2d;
    ram_cell[    1448] = 32'h509b9c79;
    ram_cell[    1449] = 32'h489d13d6;
    ram_cell[    1450] = 32'h0006b264;
    ram_cell[    1451] = 32'hce15e1b4;
    ram_cell[    1452] = 32'h74baa35c;
    ram_cell[    1453] = 32'ha3dd2b1c;
    ram_cell[    1454] = 32'h0d2b1c2c;
    ram_cell[    1455] = 32'hc0eaa73c;
    ram_cell[    1456] = 32'h3ddfe92e;
    ram_cell[    1457] = 32'h1ca13c75;
    ram_cell[    1458] = 32'h3413b78e;
    ram_cell[    1459] = 32'hae0687c2;
    ram_cell[    1460] = 32'h15477729;
    ram_cell[    1461] = 32'h4f40a49a;
    ram_cell[    1462] = 32'h9ed4f0d1;
    ram_cell[    1463] = 32'hf9e2f895;
    ram_cell[    1464] = 32'hdeb82a05;
    ram_cell[    1465] = 32'hb1c27250;
    ram_cell[    1466] = 32'h015aaabc;
    ram_cell[    1467] = 32'ha04b9197;
    ram_cell[    1468] = 32'h0a5d9f4f;
    ram_cell[    1469] = 32'h5039d86c;
    ram_cell[    1470] = 32'h28d059ab;
    ram_cell[    1471] = 32'h3c2920f0;
    ram_cell[    1472] = 32'h2c0a1e1c;
    ram_cell[    1473] = 32'h1518da64;
    ram_cell[    1474] = 32'hdc6bb69b;
    ram_cell[    1475] = 32'h0592bfa8;
    ram_cell[    1476] = 32'h4c7ae9e5;
    ram_cell[    1477] = 32'h2d570793;
    ram_cell[    1478] = 32'h89875151;
    ram_cell[    1479] = 32'h0972342f;
    ram_cell[    1480] = 32'hf6ee942b;
    ram_cell[    1481] = 32'ha44f150c;
    ram_cell[    1482] = 32'h873b5db8;
    ram_cell[    1483] = 32'hf74b80f6;
    ram_cell[    1484] = 32'h028b39dd;
    ram_cell[    1485] = 32'h6c5f85e3;
    ram_cell[    1486] = 32'h749f1d53;
    ram_cell[    1487] = 32'ha8bc8647;
    ram_cell[    1488] = 32'hd959e225;
    ram_cell[    1489] = 32'hda26996e;
    ram_cell[    1490] = 32'h546bab05;
    ram_cell[    1491] = 32'hf62d4906;
    ram_cell[    1492] = 32'h7dcd59ab;
    ram_cell[    1493] = 32'h48c31024;
    ram_cell[    1494] = 32'h950f3227;
    ram_cell[    1495] = 32'hde31ba38;
    ram_cell[    1496] = 32'h5165c6de;
    ram_cell[    1497] = 32'h8ac76fa8;
    ram_cell[    1498] = 32'h9d520442;
    ram_cell[    1499] = 32'hbe1d1e35;
    ram_cell[    1500] = 32'h76c49b7c;
    ram_cell[    1501] = 32'hebd0a3ee;
    ram_cell[    1502] = 32'h666b4641;
    ram_cell[    1503] = 32'h9e74c2ab;
    ram_cell[    1504] = 32'h38952c83;
    ram_cell[    1505] = 32'hfa61c11f;
    ram_cell[    1506] = 32'haaa1a33b;
    ram_cell[    1507] = 32'ha34da04c;
    ram_cell[    1508] = 32'h97d38702;
    ram_cell[    1509] = 32'hc9c77500;
    ram_cell[    1510] = 32'ha0e0ae15;
    ram_cell[    1511] = 32'h6fde3f17;
    ram_cell[    1512] = 32'h7856a8d7;
    ram_cell[    1513] = 32'hfd959b6c;
    ram_cell[    1514] = 32'h817e7811;
    ram_cell[    1515] = 32'h4065d5b6;
    ram_cell[    1516] = 32'h9e9b9f63;
    ram_cell[    1517] = 32'hdc531742;
    ram_cell[    1518] = 32'h123c3ceb;
    ram_cell[    1519] = 32'h61c15790;
    ram_cell[    1520] = 32'hed4c20ef;
    ram_cell[    1521] = 32'h9329ef42;
    ram_cell[    1522] = 32'h71ad4574;
    ram_cell[    1523] = 32'h3cf0258b;
    ram_cell[    1524] = 32'h7cf7a39a;
    ram_cell[    1525] = 32'h03648586;
    ram_cell[    1526] = 32'hdb73a173;
    ram_cell[    1527] = 32'h9598ca94;
    ram_cell[    1528] = 32'h36b983f8;
    ram_cell[    1529] = 32'h466e2d75;
    ram_cell[    1530] = 32'h9e822f21;
    ram_cell[    1531] = 32'ha0671c49;
    ram_cell[    1532] = 32'h11819ca9;
    ram_cell[    1533] = 32'h7ecc17dd;
    ram_cell[    1534] = 32'h5b9a7917;
    ram_cell[    1535] = 32'hf4d3943b;
    ram_cell[    1536] = 32'hf43c19da;
    ram_cell[    1537] = 32'h6e3c395d;
    ram_cell[    1538] = 32'hf264c69f;
    ram_cell[    1539] = 32'h8b71ad79;
    ram_cell[    1540] = 32'ha896e197;
    ram_cell[    1541] = 32'hee59136a;
    ram_cell[    1542] = 32'h2e0d51a8;
    ram_cell[    1543] = 32'h1a146805;
    ram_cell[    1544] = 32'h25855fa8;
    ram_cell[    1545] = 32'h62d90a86;
    ram_cell[    1546] = 32'h6f590d6d;
    ram_cell[    1547] = 32'h6151544a;
    ram_cell[    1548] = 32'h278b1a26;
    ram_cell[    1549] = 32'hbcd4e6e5;
    ram_cell[    1550] = 32'h8b194032;
    ram_cell[    1551] = 32'ha5fd972d;
    ram_cell[    1552] = 32'h3cdafaf2;
    ram_cell[    1553] = 32'hc9555388;
    ram_cell[    1554] = 32'hf1a82bf9;
    ram_cell[    1555] = 32'h1e4bc91f;
    ram_cell[    1556] = 32'hcba115a4;
    ram_cell[    1557] = 32'ha8709707;
    ram_cell[    1558] = 32'h50f9508a;
    ram_cell[    1559] = 32'h1a31ca08;
    ram_cell[    1560] = 32'hbf528ba9;
    ram_cell[    1561] = 32'hac47e81f;
    ram_cell[    1562] = 32'hdbc2dd45;
    ram_cell[    1563] = 32'hff261fff;
    ram_cell[    1564] = 32'h1d9cad02;
    ram_cell[    1565] = 32'h0ec3b0ca;
    ram_cell[    1566] = 32'h7a1fdb39;
    ram_cell[    1567] = 32'h7e2c61c4;
    ram_cell[    1568] = 32'ha228a8fe;
    ram_cell[    1569] = 32'h922e56d6;
    ram_cell[    1570] = 32'h0d8ab644;
    ram_cell[    1571] = 32'he71b7f30;
    ram_cell[    1572] = 32'h8688d944;
    ram_cell[    1573] = 32'h2c105c9d;
    ram_cell[    1574] = 32'ha4554112;
    ram_cell[    1575] = 32'h1a44e857;
    ram_cell[    1576] = 32'h73b402e1;
    ram_cell[    1577] = 32'hf380bce2;
    ram_cell[    1578] = 32'hefb3576f;
    ram_cell[    1579] = 32'hfc5196ad;
    ram_cell[    1580] = 32'h923a418f;
    ram_cell[    1581] = 32'hd943c5a1;
    ram_cell[    1582] = 32'hf4633648;
    ram_cell[    1583] = 32'h695848d3;
    ram_cell[    1584] = 32'h2eed2b4c;
    ram_cell[    1585] = 32'hdd29c792;
    ram_cell[    1586] = 32'hf79c682f;
    ram_cell[    1587] = 32'h528492d5;
    ram_cell[    1588] = 32'h19778c3b;
    ram_cell[    1589] = 32'hb7703384;
    ram_cell[    1590] = 32'h65cc44c7;
    ram_cell[    1591] = 32'h9c4b1c00;
    ram_cell[    1592] = 32'hb44025fd;
    ram_cell[    1593] = 32'h5057fc88;
    ram_cell[    1594] = 32'ha9c77eb2;
    ram_cell[    1595] = 32'h970989f4;
    ram_cell[    1596] = 32'hd023c270;
    ram_cell[    1597] = 32'hca66894d;
    ram_cell[    1598] = 32'h2cdaac48;
    ram_cell[    1599] = 32'haed48b1c;
    ram_cell[    1600] = 32'h240a833b;
    ram_cell[    1601] = 32'h61a36492;
    ram_cell[    1602] = 32'h85ba2132;
    ram_cell[    1603] = 32'h5baeb480;
    ram_cell[    1604] = 32'h2de0157a;
    ram_cell[    1605] = 32'hb40e6f19;
    ram_cell[    1606] = 32'h7f07f400;
    ram_cell[    1607] = 32'h4a619569;
    ram_cell[    1608] = 32'h63d01932;
    ram_cell[    1609] = 32'h6bc9c077;
    ram_cell[    1610] = 32'h6b905a0f;
    ram_cell[    1611] = 32'hae7275d6;
    ram_cell[    1612] = 32'h9b902797;
    ram_cell[    1613] = 32'h225eb0a6;
    ram_cell[    1614] = 32'hdc3d62f8;
    ram_cell[    1615] = 32'hd710c644;
    ram_cell[    1616] = 32'h29e12367;
    ram_cell[    1617] = 32'h7d1cd24a;
    ram_cell[    1618] = 32'ha8b3801b;
    ram_cell[    1619] = 32'h4aaca761;
    ram_cell[    1620] = 32'hc4e1e0ad;
    ram_cell[    1621] = 32'ha7e7e705;
    ram_cell[    1622] = 32'h75843f96;
    ram_cell[    1623] = 32'hecdb4b16;
    ram_cell[    1624] = 32'h032cfd5c;
    ram_cell[    1625] = 32'hc3f858d5;
    ram_cell[    1626] = 32'h5a2f79ed;
    ram_cell[    1627] = 32'h1be4c748;
    ram_cell[    1628] = 32'h759ccdc4;
    ram_cell[    1629] = 32'h07c201ae;
    ram_cell[    1630] = 32'h8c441057;
    ram_cell[    1631] = 32'h9feb2f22;
    ram_cell[    1632] = 32'h0e7a1785;
    ram_cell[    1633] = 32'h277aff15;
    ram_cell[    1634] = 32'h4776f9ec;
    ram_cell[    1635] = 32'hea16c70f;
    ram_cell[    1636] = 32'h986803fc;
    ram_cell[    1637] = 32'h040f408a;
    ram_cell[    1638] = 32'h74743214;
    ram_cell[    1639] = 32'h6fd8a940;
    ram_cell[    1640] = 32'h4f9e69e5;
    ram_cell[    1641] = 32'h273f288f;
    ram_cell[    1642] = 32'h2ff1d3bf;
    ram_cell[    1643] = 32'hebd1c8e6;
    ram_cell[    1644] = 32'hb1b1e5a9;
    ram_cell[    1645] = 32'hde77353c;
    ram_cell[    1646] = 32'h1a0cc1e6;
    ram_cell[    1647] = 32'h347ef320;
    ram_cell[    1648] = 32'h66a553eb;
    ram_cell[    1649] = 32'hca13cf61;
    ram_cell[    1650] = 32'h623e31c3;
    ram_cell[    1651] = 32'h4a9dc0f8;
    ram_cell[    1652] = 32'h66a3ebe0;
    ram_cell[    1653] = 32'h4aa9479d;
    ram_cell[    1654] = 32'hc49e131e;
    ram_cell[    1655] = 32'h07df7c41;
    ram_cell[    1656] = 32'h0c518c03;
    ram_cell[    1657] = 32'hbc6a5d0a;
    ram_cell[    1658] = 32'h4b8ef4fb;
    ram_cell[    1659] = 32'h02e78dcb;
    ram_cell[    1660] = 32'h6128695d;
    ram_cell[    1661] = 32'h53397e9c;
    ram_cell[    1662] = 32'hc6d92e25;
    ram_cell[    1663] = 32'h0cb51e7e;
    ram_cell[    1664] = 32'h23d3918b;
    ram_cell[    1665] = 32'h1814d020;
    ram_cell[    1666] = 32'hf11244c1;
    ram_cell[    1667] = 32'h40dba8e1;
    ram_cell[    1668] = 32'h188a1552;
    ram_cell[    1669] = 32'h5920b8e9;
    ram_cell[    1670] = 32'h0e557e0f;
    ram_cell[    1671] = 32'h668cd835;
    ram_cell[    1672] = 32'ha361ed72;
    ram_cell[    1673] = 32'h6e493d48;
    ram_cell[    1674] = 32'h9f5765e7;
    ram_cell[    1675] = 32'hb5e4239f;
    ram_cell[    1676] = 32'h948c463d;
    ram_cell[    1677] = 32'hcbf549b9;
    ram_cell[    1678] = 32'h3bec7e28;
    ram_cell[    1679] = 32'hf810c449;
    ram_cell[    1680] = 32'h1d16e53b;
    ram_cell[    1681] = 32'hd523c537;
    ram_cell[    1682] = 32'h8becc828;
    ram_cell[    1683] = 32'h45c7aca7;
    ram_cell[    1684] = 32'h6fd94dfc;
    ram_cell[    1685] = 32'h32b42755;
    ram_cell[    1686] = 32'h51ffcf3c;
    ram_cell[    1687] = 32'h3a30b3e6;
    ram_cell[    1688] = 32'h23ee53bd;
    ram_cell[    1689] = 32'he2332059;
    ram_cell[    1690] = 32'hf44b77ca;
    ram_cell[    1691] = 32'h5a225d5e;
    ram_cell[    1692] = 32'h87fedd8b;
    ram_cell[    1693] = 32'hb9df47a6;
    ram_cell[    1694] = 32'h368bb363;
    ram_cell[    1695] = 32'h0472b7ae;
    ram_cell[    1696] = 32'hab8926a2;
    ram_cell[    1697] = 32'h9dcdbc42;
    ram_cell[    1698] = 32'h846be3e0;
    ram_cell[    1699] = 32'h1b485486;
    ram_cell[    1700] = 32'hea424f12;
    ram_cell[    1701] = 32'h04b8163d;
    ram_cell[    1702] = 32'h7b0c03e2;
    ram_cell[    1703] = 32'he9d3143b;
    ram_cell[    1704] = 32'hca237e1f;
    ram_cell[    1705] = 32'hbd966954;
    ram_cell[    1706] = 32'hd453dbd9;
    ram_cell[    1707] = 32'h8bf0f439;
    ram_cell[    1708] = 32'h03ee8a22;
    ram_cell[    1709] = 32'hd1cfc7ad;
    ram_cell[    1710] = 32'hbc890013;
    ram_cell[    1711] = 32'h13fab017;
    ram_cell[    1712] = 32'h42483aa9;
    ram_cell[    1713] = 32'hd453e402;
    ram_cell[    1714] = 32'hcd649ad2;
    ram_cell[    1715] = 32'h2d35977e;
    ram_cell[    1716] = 32'h87d063e5;
    ram_cell[    1717] = 32'h4ad3ae57;
    ram_cell[    1718] = 32'h2d28e96c;
    ram_cell[    1719] = 32'h22401f23;
    ram_cell[    1720] = 32'h94a68b26;
    ram_cell[    1721] = 32'hbf7ae50a;
    ram_cell[    1722] = 32'hefdc619d;
    ram_cell[    1723] = 32'haa27695f;
    ram_cell[    1724] = 32'he6e3e301;
    ram_cell[    1725] = 32'h23a6557f;
    ram_cell[    1726] = 32'h7455f9ed;
    ram_cell[    1727] = 32'hbbe11865;
    ram_cell[    1728] = 32'he2d3e74f;
    ram_cell[    1729] = 32'h65f85b84;
    ram_cell[    1730] = 32'h0479b039;
    ram_cell[    1731] = 32'h5a0d8974;
    ram_cell[    1732] = 32'h1dc42001;
    ram_cell[    1733] = 32'haa40596a;
    ram_cell[    1734] = 32'h73b0064f;
    ram_cell[    1735] = 32'hef387d7c;
    ram_cell[    1736] = 32'h98934f4e;
    ram_cell[    1737] = 32'h26d4f3a3;
    ram_cell[    1738] = 32'hdcb6df6c;
    ram_cell[    1739] = 32'hc58d794b;
    ram_cell[    1740] = 32'hf11e06f1;
    ram_cell[    1741] = 32'haccb44dc;
    ram_cell[    1742] = 32'hc34f5f08;
    ram_cell[    1743] = 32'h5f193e46;
    ram_cell[    1744] = 32'h5d1fbbc0;
    ram_cell[    1745] = 32'h369e7deb;
    ram_cell[    1746] = 32'h75f9b7ec;
    ram_cell[    1747] = 32'h17e904bb;
    ram_cell[    1748] = 32'h21cc0773;
    ram_cell[    1749] = 32'ha77a038c;
    ram_cell[    1750] = 32'hf02601bf;
    ram_cell[    1751] = 32'h09a4dbde;
    ram_cell[    1752] = 32'hb57aa5d2;
    ram_cell[    1753] = 32'h52ea7520;
    ram_cell[    1754] = 32'h482c4ec3;
    ram_cell[    1755] = 32'hb5190bf7;
    ram_cell[    1756] = 32'hf4b8cbcc;
    ram_cell[    1757] = 32'h9e2cf6ff;
    ram_cell[    1758] = 32'h671c4df9;
    ram_cell[    1759] = 32'h21fd16ae;
    ram_cell[    1760] = 32'h4cf7e2b8;
    ram_cell[    1761] = 32'h02f27baa;
    ram_cell[    1762] = 32'ha298ad17;
    ram_cell[    1763] = 32'hb8552d83;
    ram_cell[    1764] = 32'h74987b3c;
    ram_cell[    1765] = 32'h2a9eb923;
    ram_cell[    1766] = 32'he3e80c25;
    ram_cell[    1767] = 32'hdcd0e77f;
    ram_cell[    1768] = 32'h7335c735;
    ram_cell[    1769] = 32'h7bf2230d;
    ram_cell[    1770] = 32'h0ca224ce;
    ram_cell[    1771] = 32'h2f959fe8;
    ram_cell[    1772] = 32'h5f853cb7;
    ram_cell[    1773] = 32'h2f8c9f8c;
    ram_cell[    1774] = 32'hb70b6db4;
    ram_cell[    1775] = 32'h679dfaaa;
    ram_cell[    1776] = 32'hce47be19;
    ram_cell[    1777] = 32'h1adf0c9c;
    ram_cell[    1778] = 32'hdf2ff44d;
    ram_cell[    1779] = 32'h5cd9c523;
    ram_cell[    1780] = 32'h4a39da00;
    ram_cell[    1781] = 32'hffdc178e;
    ram_cell[    1782] = 32'h46ec9493;
    ram_cell[    1783] = 32'h34a8a1cd;
    ram_cell[    1784] = 32'h67153289;
    ram_cell[    1785] = 32'he2f25487;
    ram_cell[    1786] = 32'h1c80a23f;
    ram_cell[    1787] = 32'h904d41da;
    ram_cell[    1788] = 32'hf2b2bcb0;
    ram_cell[    1789] = 32'h966d9f82;
    ram_cell[    1790] = 32'h27fa26d1;
    ram_cell[    1791] = 32'h3ef426ce;
    ram_cell[    1792] = 32'h3b15e27f;
    ram_cell[    1793] = 32'hb3e1b162;
    ram_cell[    1794] = 32'h3d143a49;
    ram_cell[    1795] = 32'hfc219ffd;
    ram_cell[    1796] = 32'h1441f161;
    ram_cell[    1797] = 32'had4f4dd8;
    ram_cell[    1798] = 32'h0ed3ba2c;
    ram_cell[    1799] = 32'h635050db;
    ram_cell[    1800] = 32'h5d0635da;
    ram_cell[    1801] = 32'hc000bb60;
    ram_cell[    1802] = 32'h9684245b;
    ram_cell[    1803] = 32'h9c77865b;
    ram_cell[    1804] = 32'h95085324;
    ram_cell[    1805] = 32'h28d452cb;
    ram_cell[    1806] = 32'h77c64f90;
    ram_cell[    1807] = 32'ha88a8b46;
    ram_cell[    1808] = 32'hb4d7a3dc;
    ram_cell[    1809] = 32'h89771a02;
    ram_cell[    1810] = 32'h1ccbf803;
    ram_cell[    1811] = 32'h46ea84ca;
    ram_cell[    1812] = 32'h64e4ab9a;
    ram_cell[    1813] = 32'h43acd4d4;
    ram_cell[    1814] = 32'h659cdaa6;
    ram_cell[    1815] = 32'h562ba12e;
    ram_cell[    1816] = 32'he4e7ff5d;
    ram_cell[    1817] = 32'h5f291084;
    ram_cell[    1818] = 32'h501ed45e;
    ram_cell[    1819] = 32'h6fe5a3ca;
    ram_cell[    1820] = 32'h2492cc53;
    ram_cell[    1821] = 32'hafc8433c;
    ram_cell[    1822] = 32'hb361b755;
    ram_cell[    1823] = 32'hcca402ba;
    ram_cell[    1824] = 32'h2603fd0e;
    ram_cell[    1825] = 32'habd09c73;
    ram_cell[    1826] = 32'h7c87f4d5;
    ram_cell[    1827] = 32'h8c3c201d;
    ram_cell[    1828] = 32'hfeaaec2f;
    ram_cell[    1829] = 32'h40c371d5;
    ram_cell[    1830] = 32'h5c136b60;
    ram_cell[    1831] = 32'hb2f545d5;
    ram_cell[    1832] = 32'h31951c98;
    ram_cell[    1833] = 32'hc9d073d8;
    ram_cell[    1834] = 32'h3779872c;
    ram_cell[    1835] = 32'h513522b3;
    ram_cell[    1836] = 32'hde77f16f;
    ram_cell[    1837] = 32'h4273c7d6;
    ram_cell[    1838] = 32'h9edb8bbd;
    ram_cell[    1839] = 32'h179d8739;
    ram_cell[    1840] = 32'h23102e08;
    ram_cell[    1841] = 32'h72f4cb72;
    ram_cell[    1842] = 32'hbb1c55c3;
    ram_cell[    1843] = 32'he8e39d4c;
    ram_cell[    1844] = 32'h5f858f5c;
    ram_cell[    1845] = 32'h7e24ef18;
    ram_cell[    1846] = 32'hb6254dd8;
    ram_cell[    1847] = 32'hffd4a231;
    ram_cell[    1848] = 32'hc20bff4d;
    ram_cell[    1849] = 32'h6c707859;
    ram_cell[    1850] = 32'h2f7808a1;
    ram_cell[    1851] = 32'h732ab965;
    ram_cell[    1852] = 32'h58fa5240;
    ram_cell[    1853] = 32'h8e91a9df;
    ram_cell[    1854] = 32'hd9c68538;
    ram_cell[    1855] = 32'h66b82323;
    ram_cell[    1856] = 32'h6bb50267;
    ram_cell[    1857] = 32'hc5e10b57;
    ram_cell[    1858] = 32'h15ec861f;
    ram_cell[    1859] = 32'hdfba8851;
    ram_cell[    1860] = 32'h8f25fd35;
    ram_cell[    1861] = 32'h8925874b;
    ram_cell[    1862] = 32'h8092042d;
    ram_cell[    1863] = 32'hd0a9a684;
    ram_cell[    1864] = 32'h8e72873a;
    ram_cell[    1865] = 32'h91d6aa9a;
    ram_cell[    1866] = 32'hbeb3776b;
    ram_cell[    1867] = 32'h63a89f47;
    ram_cell[    1868] = 32'h5e399cb1;
    ram_cell[    1869] = 32'h95ec34f3;
    ram_cell[    1870] = 32'hcd14747d;
    ram_cell[    1871] = 32'h3ac6a332;
    ram_cell[    1872] = 32'h8248249c;
    ram_cell[    1873] = 32'ha651c051;
    ram_cell[    1874] = 32'h28ca337f;
    ram_cell[    1875] = 32'h36419990;
    ram_cell[    1876] = 32'h73a3a3a9;
    ram_cell[    1877] = 32'h0a9aed0f;
    ram_cell[    1878] = 32'hfb6f22f5;
    ram_cell[    1879] = 32'h412572d4;
    ram_cell[    1880] = 32'h6a3e9c7f;
    ram_cell[    1881] = 32'h81f362d7;
    ram_cell[    1882] = 32'h0f247685;
    ram_cell[    1883] = 32'haebaf745;
    ram_cell[    1884] = 32'h327e1cbb;
    ram_cell[    1885] = 32'hd37e8bf5;
    ram_cell[    1886] = 32'h06727438;
    ram_cell[    1887] = 32'hf3c55217;
    ram_cell[    1888] = 32'h69e76faf;
    ram_cell[    1889] = 32'h38e92a37;
    ram_cell[    1890] = 32'h2be103f0;
    ram_cell[    1891] = 32'hf2cbc4c9;
    ram_cell[    1892] = 32'hb4f9d65a;
    ram_cell[    1893] = 32'h8a9fe417;
    ram_cell[    1894] = 32'haa062da6;
    ram_cell[    1895] = 32'h88236062;
    ram_cell[    1896] = 32'hf022c031;
    ram_cell[    1897] = 32'h4252eada;
    ram_cell[    1898] = 32'h1de544c4;
    ram_cell[    1899] = 32'h4dc54697;
    ram_cell[    1900] = 32'h05b2042a;
    ram_cell[    1901] = 32'h1e8ef155;
    ram_cell[    1902] = 32'h4d466f1b;
    ram_cell[    1903] = 32'h44d57ed9;
    ram_cell[    1904] = 32'h4012aa2f;
    ram_cell[    1905] = 32'h911b598f;
    ram_cell[    1906] = 32'h3edfb980;
    ram_cell[    1907] = 32'hc733b09d;
    ram_cell[    1908] = 32'h1356fdf3;
    ram_cell[    1909] = 32'h8e22c250;
    ram_cell[    1910] = 32'h6a467ec8;
    ram_cell[    1911] = 32'h25c4a7e5;
    ram_cell[    1912] = 32'hc562a4b7;
    ram_cell[    1913] = 32'h71fa2e9d;
    ram_cell[    1914] = 32'h3b0a9066;
    ram_cell[    1915] = 32'h752dc00e;
    ram_cell[    1916] = 32'h95ee6564;
    ram_cell[    1917] = 32'h6e3ea938;
    ram_cell[    1918] = 32'h5378bda0;
    ram_cell[    1919] = 32'heaaf8d1b;
    ram_cell[    1920] = 32'hd1f321e1;
    ram_cell[    1921] = 32'hc66b881c;
    ram_cell[    1922] = 32'h6b81dd7e;
    ram_cell[    1923] = 32'h2456a740;
    ram_cell[    1924] = 32'h837a6904;
    ram_cell[    1925] = 32'h4f54f57b;
    ram_cell[    1926] = 32'h299ce651;
    ram_cell[    1927] = 32'h5c77a50f;
    ram_cell[    1928] = 32'h4ff55508;
    ram_cell[    1929] = 32'hd2bfc34d;
    ram_cell[    1930] = 32'haa1152c0;
    ram_cell[    1931] = 32'hb45f1829;
    ram_cell[    1932] = 32'h17c503ac;
    ram_cell[    1933] = 32'h38e3e4d3;
    ram_cell[    1934] = 32'hc54274cb;
    ram_cell[    1935] = 32'h8f399476;
    ram_cell[    1936] = 32'h72b2c4cf;
    ram_cell[    1937] = 32'h27522df9;
    ram_cell[    1938] = 32'h1c64cbc4;
    ram_cell[    1939] = 32'h908d95bb;
    ram_cell[    1940] = 32'hf7a6e393;
    ram_cell[    1941] = 32'h26ec0de2;
    ram_cell[    1942] = 32'h8e675e28;
    ram_cell[    1943] = 32'hdbb43a40;
    ram_cell[    1944] = 32'h78c833f4;
    ram_cell[    1945] = 32'hbbde89b8;
    ram_cell[    1946] = 32'hf23ac774;
    ram_cell[    1947] = 32'hafcac352;
    ram_cell[    1948] = 32'h619f186c;
    ram_cell[    1949] = 32'h2a5ae9f8;
    ram_cell[    1950] = 32'h94ff94ea;
    ram_cell[    1951] = 32'h33105166;
    ram_cell[    1952] = 32'h9eb4efc6;
    ram_cell[    1953] = 32'hd12a1ef8;
    ram_cell[    1954] = 32'h6621082f;
    ram_cell[    1955] = 32'h3b29b362;
    ram_cell[    1956] = 32'h98c63c92;
    ram_cell[    1957] = 32'habb2b572;
    ram_cell[    1958] = 32'ha67e2ad5;
    ram_cell[    1959] = 32'h0b35c997;
    ram_cell[    1960] = 32'hbd626fd4;
    ram_cell[    1961] = 32'h460cc0fe;
    ram_cell[    1962] = 32'h15aaae1d;
    ram_cell[    1963] = 32'h2953c6b7;
    ram_cell[    1964] = 32'h8a7095c0;
    ram_cell[    1965] = 32'h3256ae8d;
    ram_cell[    1966] = 32'haa6565f1;
    ram_cell[    1967] = 32'hda040669;
    ram_cell[    1968] = 32'h539438c1;
    ram_cell[    1969] = 32'ha447a69b;
    ram_cell[    1970] = 32'hf23ec1c4;
    ram_cell[    1971] = 32'h5981bd17;
    ram_cell[    1972] = 32'h5629dead;
    ram_cell[    1973] = 32'h7fbee031;
    ram_cell[    1974] = 32'he2cb4e76;
    ram_cell[    1975] = 32'hed5b3013;
    ram_cell[    1976] = 32'hf6b94acf;
    ram_cell[    1977] = 32'h1a6f2e6c;
    ram_cell[    1978] = 32'h0abb9d8e;
    ram_cell[    1979] = 32'h8b30e501;
    ram_cell[    1980] = 32'hd9cdeb75;
    ram_cell[    1981] = 32'h5cb5cee6;
    ram_cell[    1982] = 32'hb5df64af;
    ram_cell[    1983] = 32'h47230a50;
    ram_cell[    1984] = 32'h5080f6ca;
    ram_cell[    1985] = 32'h1352ef95;
    ram_cell[    1986] = 32'h36503e42;
    ram_cell[    1987] = 32'h29d17f48;
    ram_cell[    1988] = 32'hece1fb38;
    ram_cell[    1989] = 32'h4bf869ac;
    ram_cell[    1990] = 32'h35aca757;
    ram_cell[    1991] = 32'h08501d85;
    ram_cell[    1992] = 32'h12e77a22;
    ram_cell[    1993] = 32'hc793cddb;
    ram_cell[    1994] = 32'hc0d7c892;
    ram_cell[    1995] = 32'he640b958;
    ram_cell[    1996] = 32'hcde09daf;
    ram_cell[    1997] = 32'hfc41da19;
    ram_cell[    1998] = 32'hec0dfeed;
    ram_cell[    1999] = 32'h6e86ec72;
    ram_cell[    2000] = 32'hec46823d;
    ram_cell[    2001] = 32'hf8a5e77e;
    ram_cell[    2002] = 32'hcb8de426;
    ram_cell[    2003] = 32'h4dbd25da;
    ram_cell[    2004] = 32'h8bab10d8;
    ram_cell[    2005] = 32'h4e1c3324;
    ram_cell[    2006] = 32'h4e6d8be4;
    ram_cell[    2007] = 32'h3ebd7cf2;
    ram_cell[    2008] = 32'h3e5bfe02;
    ram_cell[    2009] = 32'h85215035;
    ram_cell[    2010] = 32'he52f2b42;
    ram_cell[    2011] = 32'hf48cace0;
    ram_cell[    2012] = 32'h7c3927da;
    ram_cell[    2013] = 32'h3da4cc4f;
    ram_cell[    2014] = 32'hdfb4cf26;
    ram_cell[    2015] = 32'h7975730f;
    ram_cell[    2016] = 32'hef355805;
    ram_cell[    2017] = 32'h5e8c6cdc;
    ram_cell[    2018] = 32'h63b3eb62;
    ram_cell[    2019] = 32'h25a37213;
    ram_cell[    2020] = 32'hf2b61a7c;
    ram_cell[    2021] = 32'h6ce19d12;
    ram_cell[    2022] = 32'hb03904eb;
    ram_cell[    2023] = 32'h77c592a0;
    ram_cell[    2024] = 32'h15ac2693;
    ram_cell[    2025] = 32'h272cfad4;
    ram_cell[    2026] = 32'hfe99d8bd;
    ram_cell[    2027] = 32'hfc294287;
    ram_cell[    2028] = 32'hc94fd2fe;
    ram_cell[    2029] = 32'hb1f27dcf;
    ram_cell[    2030] = 32'h63c5f270;
    ram_cell[    2031] = 32'h0283227b;
    ram_cell[    2032] = 32'h66d4ef4a;
    ram_cell[    2033] = 32'h2a9b49ab;
    ram_cell[    2034] = 32'h25495d0c;
    ram_cell[    2035] = 32'h8d9c5a41;
    ram_cell[    2036] = 32'h0a2be637;
    ram_cell[    2037] = 32'h4311ce54;
    ram_cell[    2038] = 32'ha0b4d264;
    ram_cell[    2039] = 32'h758b608f;
    ram_cell[    2040] = 32'h04e792c8;
    ram_cell[    2041] = 32'h9d37e55f;
    ram_cell[    2042] = 32'h437ba589;
    ram_cell[    2043] = 32'h1f3b7616;
    ram_cell[    2044] = 32'h6b0df10f;
    ram_cell[    2045] = 32'hd88e514a;
    ram_cell[    2046] = 32'h3836aeda;
    ram_cell[    2047] = 32'h61d0af2d;
    // src matrix B
    ram_cell[    2048] = 32'h103c4e1d;
    ram_cell[    2049] = 32'h368fe3f5;
    ram_cell[    2050] = 32'h23ddb475;
    ram_cell[    2051] = 32'hf39455ec;
    ram_cell[    2052] = 32'h8e95d359;
    ram_cell[    2053] = 32'h7dfa8d74;
    ram_cell[    2054] = 32'had2e222f;
    ram_cell[    2055] = 32'hf25ebe9b;
    ram_cell[    2056] = 32'hb655fc4d;
    ram_cell[    2057] = 32'h14f396b0;
    ram_cell[    2058] = 32'h09de2985;
    ram_cell[    2059] = 32'h6557410d;
    ram_cell[    2060] = 32'h97641256;
    ram_cell[    2061] = 32'h88949b18;
    ram_cell[    2062] = 32'hb180b0c7;
    ram_cell[    2063] = 32'h769aedbe;
    ram_cell[    2064] = 32'h3b3c91f5;
    ram_cell[    2065] = 32'hf9219726;
    ram_cell[    2066] = 32'hbab914d3;
    ram_cell[    2067] = 32'h6cbdbb1f;
    ram_cell[    2068] = 32'h4d3a5aa2;
    ram_cell[    2069] = 32'h9ed9381b;
    ram_cell[    2070] = 32'h68082d95;
    ram_cell[    2071] = 32'h9cf05257;
    ram_cell[    2072] = 32'hc7c41ebc;
    ram_cell[    2073] = 32'h852b3120;
    ram_cell[    2074] = 32'hf3052f2f;
    ram_cell[    2075] = 32'h4dfb2ce6;
    ram_cell[    2076] = 32'hf1200a6d;
    ram_cell[    2077] = 32'hc5be822e;
    ram_cell[    2078] = 32'h01199d5e;
    ram_cell[    2079] = 32'h3aa490f6;
    ram_cell[    2080] = 32'h72c5ea97;
    ram_cell[    2081] = 32'h5d524eb6;
    ram_cell[    2082] = 32'hef02948d;
    ram_cell[    2083] = 32'h2be9a8dc;
    ram_cell[    2084] = 32'h54aa9816;
    ram_cell[    2085] = 32'h6a716e2a;
    ram_cell[    2086] = 32'ha9916a59;
    ram_cell[    2087] = 32'h01d867c8;
    ram_cell[    2088] = 32'hd03d3e06;
    ram_cell[    2089] = 32'he1a553ab;
    ram_cell[    2090] = 32'h41c8242b;
    ram_cell[    2091] = 32'h168f9708;
    ram_cell[    2092] = 32'ha6899545;
    ram_cell[    2093] = 32'h25ecc053;
    ram_cell[    2094] = 32'h91b6c1f1;
    ram_cell[    2095] = 32'h85d005b2;
    ram_cell[    2096] = 32'h2032ee44;
    ram_cell[    2097] = 32'hb7697bab;
    ram_cell[    2098] = 32'he5f43e54;
    ram_cell[    2099] = 32'h7f6746b9;
    ram_cell[    2100] = 32'h322726fa;
    ram_cell[    2101] = 32'hcb3c1f56;
    ram_cell[    2102] = 32'hbc2c2b99;
    ram_cell[    2103] = 32'h608604a7;
    ram_cell[    2104] = 32'h63f3c5d5;
    ram_cell[    2105] = 32'h3a421838;
    ram_cell[    2106] = 32'h39ce85a5;
    ram_cell[    2107] = 32'h552ffea1;
    ram_cell[    2108] = 32'hc1a1481d;
    ram_cell[    2109] = 32'hde62a0fc;
    ram_cell[    2110] = 32'h5ad15771;
    ram_cell[    2111] = 32'hdbe03c11;
    ram_cell[    2112] = 32'he33c3f16;
    ram_cell[    2113] = 32'hdc8e8740;
    ram_cell[    2114] = 32'hfbc6203e;
    ram_cell[    2115] = 32'hfb800ce3;
    ram_cell[    2116] = 32'h52c4c077;
    ram_cell[    2117] = 32'ha8daf4e9;
    ram_cell[    2118] = 32'h89776db9;
    ram_cell[    2119] = 32'h2fe208af;
    ram_cell[    2120] = 32'hf92889ba;
    ram_cell[    2121] = 32'h3f12f4a9;
    ram_cell[    2122] = 32'h23c54227;
    ram_cell[    2123] = 32'h2f7d93bc;
    ram_cell[    2124] = 32'h1ecb9057;
    ram_cell[    2125] = 32'h4dcedcc0;
    ram_cell[    2126] = 32'h1660e4f3;
    ram_cell[    2127] = 32'haffd2daa;
    ram_cell[    2128] = 32'h1151c967;
    ram_cell[    2129] = 32'h81565e08;
    ram_cell[    2130] = 32'h06d8c2cb;
    ram_cell[    2131] = 32'h1515846a;
    ram_cell[    2132] = 32'h0e494ada;
    ram_cell[    2133] = 32'h2dd4b9ab;
    ram_cell[    2134] = 32'h13b52c49;
    ram_cell[    2135] = 32'hc02224de;
    ram_cell[    2136] = 32'h539dc38a;
    ram_cell[    2137] = 32'h9cf0de05;
    ram_cell[    2138] = 32'hde44f148;
    ram_cell[    2139] = 32'h1302e1cf;
    ram_cell[    2140] = 32'h634822ae;
    ram_cell[    2141] = 32'h3f4f290e;
    ram_cell[    2142] = 32'h69856e18;
    ram_cell[    2143] = 32'h1eb0ad90;
    ram_cell[    2144] = 32'hfd8a623e;
    ram_cell[    2145] = 32'hacd4b9b2;
    ram_cell[    2146] = 32'he7c53ae5;
    ram_cell[    2147] = 32'he7da8182;
    ram_cell[    2148] = 32'h5dc5aefb;
    ram_cell[    2149] = 32'h92a83460;
    ram_cell[    2150] = 32'h18fa49da;
    ram_cell[    2151] = 32'hbaf6a54b;
    ram_cell[    2152] = 32'ha35f32f2;
    ram_cell[    2153] = 32'hfd3c4e1d;
    ram_cell[    2154] = 32'h26d3e39a;
    ram_cell[    2155] = 32'h879f1cc8;
    ram_cell[    2156] = 32'h3e714cc2;
    ram_cell[    2157] = 32'he402aafc;
    ram_cell[    2158] = 32'hb16dc9a2;
    ram_cell[    2159] = 32'h2f679bbd;
    ram_cell[    2160] = 32'h007f5518;
    ram_cell[    2161] = 32'h2bfaf850;
    ram_cell[    2162] = 32'hfeff8d9e;
    ram_cell[    2163] = 32'h6f431de4;
    ram_cell[    2164] = 32'h6dd1b6e7;
    ram_cell[    2165] = 32'he3796db3;
    ram_cell[    2166] = 32'h1df7c5d2;
    ram_cell[    2167] = 32'h7ea113aa;
    ram_cell[    2168] = 32'h40e80d99;
    ram_cell[    2169] = 32'hdc3ea43d;
    ram_cell[    2170] = 32'hd6e270a2;
    ram_cell[    2171] = 32'hec281ebc;
    ram_cell[    2172] = 32'h19c053fb;
    ram_cell[    2173] = 32'h89fbead7;
    ram_cell[    2174] = 32'h69aa02b2;
    ram_cell[    2175] = 32'hb5b58575;
    ram_cell[    2176] = 32'hc6228618;
    ram_cell[    2177] = 32'hf429efde;
    ram_cell[    2178] = 32'h17ce39f8;
    ram_cell[    2179] = 32'h0ff68df5;
    ram_cell[    2180] = 32'h069136a6;
    ram_cell[    2181] = 32'h1f3aaf19;
    ram_cell[    2182] = 32'h8eb1e5c8;
    ram_cell[    2183] = 32'h2893718a;
    ram_cell[    2184] = 32'h30f8d6ac;
    ram_cell[    2185] = 32'hf69d711f;
    ram_cell[    2186] = 32'h6db3a211;
    ram_cell[    2187] = 32'he59f1806;
    ram_cell[    2188] = 32'h1df3fc91;
    ram_cell[    2189] = 32'h7722465d;
    ram_cell[    2190] = 32'h3a40e4df;
    ram_cell[    2191] = 32'h303111cd;
    ram_cell[    2192] = 32'h6ba17c15;
    ram_cell[    2193] = 32'hae0a8730;
    ram_cell[    2194] = 32'h0f131632;
    ram_cell[    2195] = 32'h9d438ea5;
    ram_cell[    2196] = 32'h7dd3b421;
    ram_cell[    2197] = 32'h58ed48ce;
    ram_cell[    2198] = 32'h7abfde7b;
    ram_cell[    2199] = 32'h42bafbff;
    ram_cell[    2200] = 32'h8883cedf;
    ram_cell[    2201] = 32'hd4d0daa9;
    ram_cell[    2202] = 32'ha1b3fbee;
    ram_cell[    2203] = 32'h1ff54388;
    ram_cell[    2204] = 32'h0c719c8f;
    ram_cell[    2205] = 32'h488098e9;
    ram_cell[    2206] = 32'hbd10fc60;
    ram_cell[    2207] = 32'habe49f47;
    ram_cell[    2208] = 32'h186a4a0e;
    ram_cell[    2209] = 32'hb4cc38d9;
    ram_cell[    2210] = 32'h22a7cee7;
    ram_cell[    2211] = 32'h6418e0c4;
    ram_cell[    2212] = 32'h47b49628;
    ram_cell[    2213] = 32'h851c53a6;
    ram_cell[    2214] = 32'h8d74536a;
    ram_cell[    2215] = 32'he98e37e7;
    ram_cell[    2216] = 32'had62a4ad;
    ram_cell[    2217] = 32'h269fcab8;
    ram_cell[    2218] = 32'he7719295;
    ram_cell[    2219] = 32'h7611fd28;
    ram_cell[    2220] = 32'h242089a9;
    ram_cell[    2221] = 32'hda0dbc4c;
    ram_cell[    2222] = 32'h3319d2dc;
    ram_cell[    2223] = 32'h02cfd24f;
    ram_cell[    2224] = 32'hcb4f8451;
    ram_cell[    2225] = 32'hcbdfde0a;
    ram_cell[    2226] = 32'hd0072327;
    ram_cell[    2227] = 32'h4ba4115e;
    ram_cell[    2228] = 32'h6e83501d;
    ram_cell[    2229] = 32'hfb221d57;
    ram_cell[    2230] = 32'h85de4187;
    ram_cell[    2231] = 32'h25a26b25;
    ram_cell[    2232] = 32'hcebe2847;
    ram_cell[    2233] = 32'h3d9940f7;
    ram_cell[    2234] = 32'h8b71ed2f;
    ram_cell[    2235] = 32'h00eaa746;
    ram_cell[    2236] = 32'h93983606;
    ram_cell[    2237] = 32'hffed4578;
    ram_cell[    2238] = 32'hbda22876;
    ram_cell[    2239] = 32'h77823b4e;
    ram_cell[    2240] = 32'h8a2e5155;
    ram_cell[    2241] = 32'ha5f26dec;
    ram_cell[    2242] = 32'h1116c642;
    ram_cell[    2243] = 32'h60c4e6b9;
    ram_cell[    2244] = 32'h8e82499c;
    ram_cell[    2245] = 32'hefd44c62;
    ram_cell[    2246] = 32'hae2e1fb4;
    ram_cell[    2247] = 32'ha4dc666c;
    ram_cell[    2248] = 32'hf0f0f2a5;
    ram_cell[    2249] = 32'hd7e70f97;
    ram_cell[    2250] = 32'hb5145f00;
    ram_cell[    2251] = 32'h0fd4b0af;
    ram_cell[    2252] = 32'hf164a236;
    ram_cell[    2253] = 32'h8753ccf9;
    ram_cell[    2254] = 32'hc580b6be;
    ram_cell[    2255] = 32'he3199ae4;
    ram_cell[    2256] = 32'h46215271;
    ram_cell[    2257] = 32'hbc4d56b8;
    ram_cell[    2258] = 32'h58be509d;
    ram_cell[    2259] = 32'h920bb45a;
    ram_cell[    2260] = 32'h29dd20c9;
    ram_cell[    2261] = 32'hdf881ee5;
    ram_cell[    2262] = 32'hb7e50d6e;
    ram_cell[    2263] = 32'h7f107657;
    ram_cell[    2264] = 32'h1d9fa4bc;
    ram_cell[    2265] = 32'hb03837be;
    ram_cell[    2266] = 32'hbf90c768;
    ram_cell[    2267] = 32'hbf848f9c;
    ram_cell[    2268] = 32'hb1919f05;
    ram_cell[    2269] = 32'hb3bd9356;
    ram_cell[    2270] = 32'h5ec82060;
    ram_cell[    2271] = 32'h880f3854;
    ram_cell[    2272] = 32'hc708a24f;
    ram_cell[    2273] = 32'hdba4dd39;
    ram_cell[    2274] = 32'hccd6216a;
    ram_cell[    2275] = 32'hd97ae13d;
    ram_cell[    2276] = 32'h0cee9d9c;
    ram_cell[    2277] = 32'h68149712;
    ram_cell[    2278] = 32'hb512e6f1;
    ram_cell[    2279] = 32'h2a583d86;
    ram_cell[    2280] = 32'h299fd7b1;
    ram_cell[    2281] = 32'h75790b06;
    ram_cell[    2282] = 32'hc26168bc;
    ram_cell[    2283] = 32'h73a4fabe;
    ram_cell[    2284] = 32'h9b526c8a;
    ram_cell[    2285] = 32'ha701ef49;
    ram_cell[    2286] = 32'h865edce2;
    ram_cell[    2287] = 32'h2729507f;
    ram_cell[    2288] = 32'h735fefa3;
    ram_cell[    2289] = 32'hbc4beb68;
    ram_cell[    2290] = 32'hec67c42f;
    ram_cell[    2291] = 32'h611ff291;
    ram_cell[    2292] = 32'h9d850072;
    ram_cell[    2293] = 32'h66faf342;
    ram_cell[    2294] = 32'h198dd754;
    ram_cell[    2295] = 32'hd1fff098;
    ram_cell[    2296] = 32'he73c288a;
    ram_cell[    2297] = 32'hf6d1e036;
    ram_cell[    2298] = 32'h738f1d83;
    ram_cell[    2299] = 32'hb85a465b;
    ram_cell[    2300] = 32'h3d77ef1b;
    ram_cell[    2301] = 32'h21dde37f;
    ram_cell[    2302] = 32'hafcd2139;
    ram_cell[    2303] = 32'ha650c098;
    ram_cell[    2304] = 32'h0332e0f4;
    ram_cell[    2305] = 32'hef06a9cd;
    ram_cell[    2306] = 32'h6205b36b;
    ram_cell[    2307] = 32'haf97de92;
    ram_cell[    2308] = 32'hfb315297;
    ram_cell[    2309] = 32'h6b1d3576;
    ram_cell[    2310] = 32'haff60297;
    ram_cell[    2311] = 32'h8aaf75f4;
    ram_cell[    2312] = 32'hcb5acee4;
    ram_cell[    2313] = 32'hf2a83da9;
    ram_cell[    2314] = 32'ha528c36a;
    ram_cell[    2315] = 32'h13a86890;
    ram_cell[    2316] = 32'h8aee5424;
    ram_cell[    2317] = 32'hc652f69e;
    ram_cell[    2318] = 32'hfdfb1fbe;
    ram_cell[    2319] = 32'hcc177eee;
    ram_cell[    2320] = 32'hc585aad6;
    ram_cell[    2321] = 32'h2551e899;
    ram_cell[    2322] = 32'h9cfa88de;
    ram_cell[    2323] = 32'h850bf22b;
    ram_cell[    2324] = 32'hfcc33263;
    ram_cell[    2325] = 32'h0e903db9;
    ram_cell[    2326] = 32'h3e300324;
    ram_cell[    2327] = 32'h8ed83b9f;
    ram_cell[    2328] = 32'hb5d5565f;
    ram_cell[    2329] = 32'h3ed60055;
    ram_cell[    2330] = 32'he6bbb81f;
    ram_cell[    2331] = 32'h2b67150f;
    ram_cell[    2332] = 32'h5e123bda;
    ram_cell[    2333] = 32'hc9f8c8ec;
    ram_cell[    2334] = 32'he4ab70c5;
    ram_cell[    2335] = 32'hd172c044;
    ram_cell[    2336] = 32'h90601a13;
    ram_cell[    2337] = 32'hcd3ccf68;
    ram_cell[    2338] = 32'h1f4f5d5a;
    ram_cell[    2339] = 32'h5670f658;
    ram_cell[    2340] = 32'h7cfdead3;
    ram_cell[    2341] = 32'h304c64ea;
    ram_cell[    2342] = 32'hc3c2278c;
    ram_cell[    2343] = 32'hea50e617;
    ram_cell[    2344] = 32'h3c8afa71;
    ram_cell[    2345] = 32'h2c8e609b;
    ram_cell[    2346] = 32'h4cd54042;
    ram_cell[    2347] = 32'hd179e184;
    ram_cell[    2348] = 32'h571927ba;
    ram_cell[    2349] = 32'h6c245235;
    ram_cell[    2350] = 32'h21b19dcf;
    ram_cell[    2351] = 32'hbe909463;
    ram_cell[    2352] = 32'h283c3856;
    ram_cell[    2353] = 32'h5f47169e;
    ram_cell[    2354] = 32'h327dbb06;
    ram_cell[    2355] = 32'h3bb9d0e5;
    ram_cell[    2356] = 32'h09f9c052;
    ram_cell[    2357] = 32'h014f21a4;
    ram_cell[    2358] = 32'hac6d73d3;
    ram_cell[    2359] = 32'h2092b03e;
    ram_cell[    2360] = 32'h1c98cb3c;
    ram_cell[    2361] = 32'h7e1ded7f;
    ram_cell[    2362] = 32'hb2bf6491;
    ram_cell[    2363] = 32'hc1509818;
    ram_cell[    2364] = 32'h51e840f1;
    ram_cell[    2365] = 32'h91b54a06;
    ram_cell[    2366] = 32'h3b8246b9;
    ram_cell[    2367] = 32'hedd8d379;
    ram_cell[    2368] = 32'hcdd88c37;
    ram_cell[    2369] = 32'h9b4767bf;
    ram_cell[    2370] = 32'h80f738f1;
    ram_cell[    2371] = 32'heb9324dc;
    ram_cell[    2372] = 32'h3e8f0dd6;
    ram_cell[    2373] = 32'h820a1b58;
    ram_cell[    2374] = 32'hdacc927b;
    ram_cell[    2375] = 32'hc4bc5ba6;
    ram_cell[    2376] = 32'h3a4c9129;
    ram_cell[    2377] = 32'hda156bca;
    ram_cell[    2378] = 32'h02317b98;
    ram_cell[    2379] = 32'h1ed6066e;
    ram_cell[    2380] = 32'h67cfe5df;
    ram_cell[    2381] = 32'h5b9ad7de;
    ram_cell[    2382] = 32'h3d0c184e;
    ram_cell[    2383] = 32'hf32ad8bc;
    ram_cell[    2384] = 32'h5895d54f;
    ram_cell[    2385] = 32'hdfdcb062;
    ram_cell[    2386] = 32'hd287abb7;
    ram_cell[    2387] = 32'h3713a249;
    ram_cell[    2388] = 32'h01e2f622;
    ram_cell[    2389] = 32'hf46006cd;
    ram_cell[    2390] = 32'h279332d3;
    ram_cell[    2391] = 32'h11651232;
    ram_cell[    2392] = 32'h51864148;
    ram_cell[    2393] = 32'h50386c17;
    ram_cell[    2394] = 32'h37662bf3;
    ram_cell[    2395] = 32'ha23be20d;
    ram_cell[    2396] = 32'h1cbc7cf1;
    ram_cell[    2397] = 32'h5230e287;
    ram_cell[    2398] = 32'h879b6316;
    ram_cell[    2399] = 32'h2420545d;
    ram_cell[    2400] = 32'hda7dad83;
    ram_cell[    2401] = 32'hcac110c5;
    ram_cell[    2402] = 32'h8a0b3ade;
    ram_cell[    2403] = 32'h426e0560;
    ram_cell[    2404] = 32'hb8152b9a;
    ram_cell[    2405] = 32'h3d0b1a88;
    ram_cell[    2406] = 32'hde041e09;
    ram_cell[    2407] = 32'h057c60a3;
    ram_cell[    2408] = 32'h7ec6aa2b;
    ram_cell[    2409] = 32'h0bfad378;
    ram_cell[    2410] = 32'h314e915b;
    ram_cell[    2411] = 32'hb3868f76;
    ram_cell[    2412] = 32'h8687bf6a;
    ram_cell[    2413] = 32'h6f1de3dd;
    ram_cell[    2414] = 32'h13bb2af4;
    ram_cell[    2415] = 32'hb8c8e174;
    ram_cell[    2416] = 32'he9e00c9a;
    ram_cell[    2417] = 32'he1ce193e;
    ram_cell[    2418] = 32'h86cef0a5;
    ram_cell[    2419] = 32'h3a22d27a;
    ram_cell[    2420] = 32'h37a51e34;
    ram_cell[    2421] = 32'hbe3f7d8c;
    ram_cell[    2422] = 32'hbcac03bb;
    ram_cell[    2423] = 32'h82eb7184;
    ram_cell[    2424] = 32'h8a5b29b2;
    ram_cell[    2425] = 32'h9e68ed6b;
    ram_cell[    2426] = 32'h9145ebfa;
    ram_cell[    2427] = 32'h0f05589e;
    ram_cell[    2428] = 32'h3583ad98;
    ram_cell[    2429] = 32'hf7939fbf;
    ram_cell[    2430] = 32'h83cc03e4;
    ram_cell[    2431] = 32'h841e9d23;
    ram_cell[    2432] = 32'h304b041c;
    ram_cell[    2433] = 32'h4ed1750f;
    ram_cell[    2434] = 32'h93e147fa;
    ram_cell[    2435] = 32'h27bb9871;
    ram_cell[    2436] = 32'hff5d7b88;
    ram_cell[    2437] = 32'h097aeaf8;
    ram_cell[    2438] = 32'hfd5e93ba;
    ram_cell[    2439] = 32'h19a78d1b;
    ram_cell[    2440] = 32'h34086555;
    ram_cell[    2441] = 32'h741b36cb;
    ram_cell[    2442] = 32'h4ee4f128;
    ram_cell[    2443] = 32'h8f6ff2c9;
    ram_cell[    2444] = 32'hac2111f5;
    ram_cell[    2445] = 32'h01f2a5de;
    ram_cell[    2446] = 32'h5663f7b4;
    ram_cell[    2447] = 32'hf97f4a0c;
    ram_cell[    2448] = 32'h1083de70;
    ram_cell[    2449] = 32'h9f5edf0b;
    ram_cell[    2450] = 32'h2211ea03;
    ram_cell[    2451] = 32'hd7c918bb;
    ram_cell[    2452] = 32'h5038dd94;
    ram_cell[    2453] = 32'heaa37ad8;
    ram_cell[    2454] = 32'h87f5fa85;
    ram_cell[    2455] = 32'h8a3b008b;
    ram_cell[    2456] = 32'h13f4ee7b;
    ram_cell[    2457] = 32'h70477f07;
    ram_cell[    2458] = 32'hfd8452ea;
    ram_cell[    2459] = 32'hf0ae4828;
    ram_cell[    2460] = 32'h0efe3b56;
    ram_cell[    2461] = 32'he6c49321;
    ram_cell[    2462] = 32'hc226c655;
    ram_cell[    2463] = 32'h6813376d;
    ram_cell[    2464] = 32'ha4ac44a6;
    ram_cell[    2465] = 32'h3cd96dd3;
    ram_cell[    2466] = 32'hcfbf765a;
    ram_cell[    2467] = 32'h56951841;
    ram_cell[    2468] = 32'h334f11f5;
    ram_cell[    2469] = 32'he084b4a7;
    ram_cell[    2470] = 32'h42061a99;
    ram_cell[    2471] = 32'h68eb713d;
    ram_cell[    2472] = 32'hda22e409;
    ram_cell[    2473] = 32'hcb6f2212;
    ram_cell[    2474] = 32'hcf02e1a7;
    ram_cell[    2475] = 32'hb58d020a;
    ram_cell[    2476] = 32'h5a1290e5;
    ram_cell[    2477] = 32'haa29ca1a;
    ram_cell[    2478] = 32'h26e3b127;
    ram_cell[    2479] = 32'ha3ccc454;
    ram_cell[    2480] = 32'hc9b30742;
    ram_cell[    2481] = 32'h2536ed07;
    ram_cell[    2482] = 32'h28e62f36;
    ram_cell[    2483] = 32'hda70340a;
    ram_cell[    2484] = 32'h3db54886;
    ram_cell[    2485] = 32'h0c68cb4a;
    ram_cell[    2486] = 32'hb89eb7dc;
    ram_cell[    2487] = 32'h9acf44f8;
    ram_cell[    2488] = 32'h26a29170;
    ram_cell[    2489] = 32'ha0da8ca0;
    ram_cell[    2490] = 32'h6e5c58d1;
    ram_cell[    2491] = 32'hff9e2065;
    ram_cell[    2492] = 32'h08529207;
    ram_cell[    2493] = 32'h315e394c;
    ram_cell[    2494] = 32'h89902b1a;
    ram_cell[    2495] = 32'h70d153d9;
    ram_cell[    2496] = 32'h5cff892b;
    ram_cell[    2497] = 32'hcef658c3;
    ram_cell[    2498] = 32'hca4aed73;
    ram_cell[    2499] = 32'h8f94b3fb;
    ram_cell[    2500] = 32'he55a0837;
    ram_cell[    2501] = 32'h47171f07;
    ram_cell[    2502] = 32'hab39862d;
    ram_cell[    2503] = 32'h229e9cb6;
    ram_cell[    2504] = 32'hd55504b1;
    ram_cell[    2505] = 32'h81d16598;
    ram_cell[    2506] = 32'h4b3f2754;
    ram_cell[    2507] = 32'hff6796d6;
    ram_cell[    2508] = 32'had792b70;
    ram_cell[    2509] = 32'h7b66360d;
    ram_cell[    2510] = 32'hbe7ed4d2;
    ram_cell[    2511] = 32'ha7900b41;
    ram_cell[    2512] = 32'h6cba8968;
    ram_cell[    2513] = 32'h104883cd;
    ram_cell[    2514] = 32'h438d4c2a;
    ram_cell[    2515] = 32'h5f93fe15;
    ram_cell[    2516] = 32'h2ce27f76;
    ram_cell[    2517] = 32'h586e585b;
    ram_cell[    2518] = 32'he00bdadb;
    ram_cell[    2519] = 32'hf08992f1;
    ram_cell[    2520] = 32'h011e4be0;
    ram_cell[    2521] = 32'hdf2744eb;
    ram_cell[    2522] = 32'h0bb47fd9;
    ram_cell[    2523] = 32'h37ca1116;
    ram_cell[    2524] = 32'h7747358d;
    ram_cell[    2525] = 32'h8b57f0bb;
    ram_cell[    2526] = 32'hd55e05de;
    ram_cell[    2527] = 32'h0c34eac7;
    ram_cell[    2528] = 32'h083e5d71;
    ram_cell[    2529] = 32'h94f0810b;
    ram_cell[    2530] = 32'hfb05974e;
    ram_cell[    2531] = 32'h052f97d4;
    ram_cell[    2532] = 32'h2ab726b1;
    ram_cell[    2533] = 32'h7ce3ae6b;
    ram_cell[    2534] = 32'h270f28ec;
    ram_cell[    2535] = 32'h6e95fc1f;
    ram_cell[    2536] = 32'hc39ea790;
    ram_cell[    2537] = 32'h75735b60;
    ram_cell[    2538] = 32'h34c8f52b;
    ram_cell[    2539] = 32'hc4bd8caa;
    ram_cell[    2540] = 32'he6d5ad94;
    ram_cell[    2541] = 32'hcc82cb0a;
    ram_cell[    2542] = 32'h6c4ae6ba;
    ram_cell[    2543] = 32'h2d83e9c6;
    ram_cell[    2544] = 32'hed6982ec;
    ram_cell[    2545] = 32'h17f019aa;
    ram_cell[    2546] = 32'he16c4fdf;
    ram_cell[    2547] = 32'haf65dac7;
    ram_cell[    2548] = 32'h63638890;
    ram_cell[    2549] = 32'h6dcd9f89;
    ram_cell[    2550] = 32'h1970c5b3;
    ram_cell[    2551] = 32'h3e4cd6b2;
    ram_cell[    2552] = 32'h21cd2efc;
    ram_cell[    2553] = 32'h3c76c4a6;
    ram_cell[    2554] = 32'he36fff3a;
    ram_cell[    2555] = 32'hfa72b932;
    ram_cell[    2556] = 32'h6ed6e3b3;
    ram_cell[    2557] = 32'h00893d8d;
    ram_cell[    2558] = 32'h5be7f369;
    ram_cell[    2559] = 32'hb6e9a370;
    ram_cell[    2560] = 32'heab31cac;
    ram_cell[    2561] = 32'h6221ad3d;
    ram_cell[    2562] = 32'h4de0bcc2;
    ram_cell[    2563] = 32'h8a0c85f5;
    ram_cell[    2564] = 32'hf8690358;
    ram_cell[    2565] = 32'ha6fcfa1b;
    ram_cell[    2566] = 32'he5cf686f;
    ram_cell[    2567] = 32'h6b06ecd0;
    ram_cell[    2568] = 32'hb7534cd8;
    ram_cell[    2569] = 32'h93314bf1;
    ram_cell[    2570] = 32'h87b08e77;
    ram_cell[    2571] = 32'h6391b9bf;
    ram_cell[    2572] = 32'h3a4b0fb5;
    ram_cell[    2573] = 32'hf1a077e3;
    ram_cell[    2574] = 32'h192eeea6;
    ram_cell[    2575] = 32'h55332852;
    ram_cell[    2576] = 32'h93146b5e;
    ram_cell[    2577] = 32'ha7eb3037;
    ram_cell[    2578] = 32'h2f1f656d;
    ram_cell[    2579] = 32'hdf2da349;
    ram_cell[    2580] = 32'ha9d73033;
    ram_cell[    2581] = 32'h820c54d6;
    ram_cell[    2582] = 32'h453e28b5;
    ram_cell[    2583] = 32'h0bfe33be;
    ram_cell[    2584] = 32'h9e344417;
    ram_cell[    2585] = 32'ha523f344;
    ram_cell[    2586] = 32'hb19a5dd7;
    ram_cell[    2587] = 32'hbc6e8572;
    ram_cell[    2588] = 32'haf045492;
    ram_cell[    2589] = 32'hb9a70c82;
    ram_cell[    2590] = 32'h3d1244b1;
    ram_cell[    2591] = 32'h56d49adc;
    ram_cell[    2592] = 32'h46bb552c;
    ram_cell[    2593] = 32'hafd2d6fa;
    ram_cell[    2594] = 32'h45b6ed4d;
    ram_cell[    2595] = 32'h2abeb346;
    ram_cell[    2596] = 32'h6be0ddbb;
    ram_cell[    2597] = 32'h0684c801;
    ram_cell[    2598] = 32'h08f3ceb8;
    ram_cell[    2599] = 32'h67023a19;
    ram_cell[    2600] = 32'hb99d36de;
    ram_cell[    2601] = 32'h681f5342;
    ram_cell[    2602] = 32'h32f59934;
    ram_cell[    2603] = 32'h19dd73ef;
    ram_cell[    2604] = 32'h7d07da83;
    ram_cell[    2605] = 32'h0ae0370f;
    ram_cell[    2606] = 32'h7b3f975d;
    ram_cell[    2607] = 32'hdc5596a1;
    ram_cell[    2608] = 32'hedd8ddda;
    ram_cell[    2609] = 32'h90dee81a;
    ram_cell[    2610] = 32'h69ffe11a;
    ram_cell[    2611] = 32'hf1e26bc1;
    ram_cell[    2612] = 32'ha4bb4337;
    ram_cell[    2613] = 32'h53213089;
    ram_cell[    2614] = 32'ha1096be3;
    ram_cell[    2615] = 32'h5f3ce87f;
    ram_cell[    2616] = 32'hafe2736d;
    ram_cell[    2617] = 32'ha2ccca9e;
    ram_cell[    2618] = 32'hac70db18;
    ram_cell[    2619] = 32'h8ab14e7a;
    ram_cell[    2620] = 32'h4b3a1b2c;
    ram_cell[    2621] = 32'he47410d3;
    ram_cell[    2622] = 32'hb527d111;
    ram_cell[    2623] = 32'h607c4c4e;
    ram_cell[    2624] = 32'h5c82c006;
    ram_cell[    2625] = 32'h7b4f0465;
    ram_cell[    2626] = 32'hf48ce993;
    ram_cell[    2627] = 32'h80b1e4cc;
    ram_cell[    2628] = 32'h6ef12455;
    ram_cell[    2629] = 32'he85e749c;
    ram_cell[    2630] = 32'hc902d6e2;
    ram_cell[    2631] = 32'h066cda79;
    ram_cell[    2632] = 32'he44e1b00;
    ram_cell[    2633] = 32'hd3e3e89c;
    ram_cell[    2634] = 32'hee7ee36a;
    ram_cell[    2635] = 32'h32a8206c;
    ram_cell[    2636] = 32'hf0b1bbbc;
    ram_cell[    2637] = 32'hd64a9a98;
    ram_cell[    2638] = 32'h3287c349;
    ram_cell[    2639] = 32'h5c851ce3;
    ram_cell[    2640] = 32'h1c63f067;
    ram_cell[    2641] = 32'h1a0a2f77;
    ram_cell[    2642] = 32'h7650a354;
    ram_cell[    2643] = 32'h94b53eaa;
    ram_cell[    2644] = 32'h121d5e3b;
    ram_cell[    2645] = 32'hbe8e42c8;
    ram_cell[    2646] = 32'he764ed09;
    ram_cell[    2647] = 32'h11ddad1d;
    ram_cell[    2648] = 32'h587ff145;
    ram_cell[    2649] = 32'h42611507;
    ram_cell[    2650] = 32'h2899ac03;
    ram_cell[    2651] = 32'h761efcd4;
    ram_cell[    2652] = 32'h7da5db2c;
    ram_cell[    2653] = 32'h52acaf6d;
    ram_cell[    2654] = 32'hc965d3c2;
    ram_cell[    2655] = 32'hc493ff68;
    ram_cell[    2656] = 32'h5872fc9a;
    ram_cell[    2657] = 32'hd5552ad6;
    ram_cell[    2658] = 32'h805bbe9f;
    ram_cell[    2659] = 32'hced735fa;
    ram_cell[    2660] = 32'he000c1c5;
    ram_cell[    2661] = 32'h36df3182;
    ram_cell[    2662] = 32'heacdea08;
    ram_cell[    2663] = 32'hd699ba3e;
    ram_cell[    2664] = 32'hc3820db7;
    ram_cell[    2665] = 32'h9b8da8e9;
    ram_cell[    2666] = 32'h0614d06f;
    ram_cell[    2667] = 32'h795bb628;
    ram_cell[    2668] = 32'hd73b4498;
    ram_cell[    2669] = 32'h033a5873;
    ram_cell[    2670] = 32'h1c0ed9c6;
    ram_cell[    2671] = 32'hc02ca27b;
    ram_cell[    2672] = 32'h715e9809;
    ram_cell[    2673] = 32'hb455f7b0;
    ram_cell[    2674] = 32'h451391b0;
    ram_cell[    2675] = 32'h53b7f0f9;
    ram_cell[    2676] = 32'h119b406b;
    ram_cell[    2677] = 32'h15287c6e;
    ram_cell[    2678] = 32'hf06dcc17;
    ram_cell[    2679] = 32'h3b15b409;
    ram_cell[    2680] = 32'hfafc180a;
    ram_cell[    2681] = 32'h202265c2;
    ram_cell[    2682] = 32'h7ecee22a;
    ram_cell[    2683] = 32'h7aabb714;
    ram_cell[    2684] = 32'h166335d0;
    ram_cell[    2685] = 32'hce560d1e;
    ram_cell[    2686] = 32'h6ee1db78;
    ram_cell[    2687] = 32'h16aa1722;
    ram_cell[    2688] = 32'ha3b21196;
    ram_cell[    2689] = 32'h041db6eb;
    ram_cell[    2690] = 32'hef122c4e;
    ram_cell[    2691] = 32'h73ae09ce;
    ram_cell[    2692] = 32'h0c3c1fc4;
    ram_cell[    2693] = 32'h3cf9a7ef;
    ram_cell[    2694] = 32'h9a0d97b8;
    ram_cell[    2695] = 32'h4835d45c;
    ram_cell[    2696] = 32'h4b676988;
    ram_cell[    2697] = 32'hf968a87b;
    ram_cell[    2698] = 32'h83ae709c;
    ram_cell[    2699] = 32'h637e147d;
    ram_cell[    2700] = 32'h3083364a;
    ram_cell[    2701] = 32'h3b3c07f0;
    ram_cell[    2702] = 32'h8e771c10;
    ram_cell[    2703] = 32'h781fe998;
    ram_cell[    2704] = 32'hecb219bf;
    ram_cell[    2705] = 32'h44d34dd9;
    ram_cell[    2706] = 32'hbe709416;
    ram_cell[    2707] = 32'h40071d7a;
    ram_cell[    2708] = 32'h3e00662f;
    ram_cell[    2709] = 32'h2bbec534;
    ram_cell[    2710] = 32'h4414fa5a;
    ram_cell[    2711] = 32'h3f561d48;
    ram_cell[    2712] = 32'hbf304dd8;
    ram_cell[    2713] = 32'ha7b4d996;
    ram_cell[    2714] = 32'h997ba235;
    ram_cell[    2715] = 32'h3fb2aafe;
    ram_cell[    2716] = 32'hf2dfb308;
    ram_cell[    2717] = 32'h771b2d2f;
    ram_cell[    2718] = 32'ha9d889c0;
    ram_cell[    2719] = 32'h2c003e94;
    ram_cell[    2720] = 32'h4651bf5e;
    ram_cell[    2721] = 32'h2f46a645;
    ram_cell[    2722] = 32'hc49e7a3d;
    ram_cell[    2723] = 32'h01a1ba32;
    ram_cell[    2724] = 32'h265f7cb0;
    ram_cell[    2725] = 32'h65a97b5f;
    ram_cell[    2726] = 32'h0043f6c6;
    ram_cell[    2727] = 32'hc0d12361;
    ram_cell[    2728] = 32'h87f4c6cb;
    ram_cell[    2729] = 32'h9690c292;
    ram_cell[    2730] = 32'hf8b76db6;
    ram_cell[    2731] = 32'hdbb18db5;
    ram_cell[    2732] = 32'h859414f0;
    ram_cell[    2733] = 32'h5369e910;
    ram_cell[    2734] = 32'h458853cd;
    ram_cell[    2735] = 32'h7b997eb4;
    ram_cell[    2736] = 32'hc8bb040d;
    ram_cell[    2737] = 32'hd0369942;
    ram_cell[    2738] = 32'hf28e3d82;
    ram_cell[    2739] = 32'h9859477a;
    ram_cell[    2740] = 32'h4f7a0a6a;
    ram_cell[    2741] = 32'hfda25fd7;
    ram_cell[    2742] = 32'hb249b6f0;
    ram_cell[    2743] = 32'h052e6ee4;
    ram_cell[    2744] = 32'h233d7f43;
    ram_cell[    2745] = 32'h756151bd;
    ram_cell[    2746] = 32'h666a59fc;
    ram_cell[    2747] = 32'hd55e66a2;
    ram_cell[    2748] = 32'h5a8f642d;
    ram_cell[    2749] = 32'hd4e43457;
    ram_cell[    2750] = 32'h04764238;
    ram_cell[    2751] = 32'h024b2a45;
    ram_cell[    2752] = 32'h264c739a;
    ram_cell[    2753] = 32'h699524cf;
    ram_cell[    2754] = 32'h53cd1fca;
    ram_cell[    2755] = 32'hebce9e2a;
    ram_cell[    2756] = 32'h2725f8be;
    ram_cell[    2757] = 32'he6a89003;
    ram_cell[    2758] = 32'hbf9a97e6;
    ram_cell[    2759] = 32'h98f6b374;
    ram_cell[    2760] = 32'h18c2ea4b;
    ram_cell[    2761] = 32'h2ef826f9;
    ram_cell[    2762] = 32'hf1431e21;
    ram_cell[    2763] = 32'h102aeddb;
    ram_cell[    2764] = 32'h45381f11;
    ram_cell[    2765] = 32'hb99bdedd;
    ram_cell[    2766] = 32'h1ddc53b6;
    ram_cell[    2767] = 32'h8ebb8a69;
    ram_cell[    2768] = 32'h62b38082;
    ram_cell[    2769] = 32'h98ac750e;
    ram_cell[    2770] = 32'h8a8a0ead;
    ram_cell[    2771] = 32'hca44b407;
    ram_cell[    2772] = 32'h694960c1;
    ram_cell[    2773] = 32'h9390d1d7;
    ram_cell[    2774] = 32'h9fa05323;
    ram_cell[    2775] = 32'h9eaa2043;
    ram_cell[    2776] = 32'h33775575;
    ram_cell[    2777] = 32'hf56c64e8;
    ram_cell[    2778] = 32'hfa897c10;
    ram_cell[    2779] = 32'h980a7102;
    ram_cell[    2780] = 32'h2a0c75e0;
    ram_cell[    2781] = 32'h77b54d55;
    ram_cell[    2782] = 32'h2319e27f;
    ram_cell[    2783] = 32'hf4556098;
    ram_cell[    2784] = 32'h309fb053;
    ram_cell[    2785] = 32'h208e5820;
    ram_cell[    2786] = 32'h053526de;
    ram_cell[    2787] = 32'h855ed359;
    ram_cell[    2788] = 32'hd09d7df4;
    ram_cell[    2789] = 32'ha0f1980e;
    ram_cell[    2790] = 32'h84a2b92c;
    ram_cell[    2791] = 32'h3d38890c;
    ram_cell[    2792] = 32'h6ad3b545;
    ram_cell[    2793] = 32'h989a3bfe;
    ram_cell[    2794] = 32'h73ec2a8e;
    ram_cell[    2795] = 32'h40daaaea;
    ram_cell[    2796] = 32'hd477fb5d;
    ram_cell[    2797] = 32'h8f10abe1;
    ram_cell[    2798] = 32'h68777e91;
    ram_cell[    2799] = 32'h4b0b2455;
    ram_cell[    2800] = 32'hf0550aa3;
    ram_cell[    2801] = 32'h0cefd85f;
    ram_cell[    2802] = 32'h34ee9bde;
    ram_cell[    2803] = 32'h34813297;
    ram_cell[    2804] = 32'heb36c03b;
    ram_cell[    2805] = 32'h875ba83c;
    ram_cell[    2806] = 32'h3b57b3ac;
    ram_cell[    2807] = 32'hce365bce;
    ram_cell[    2808] = 32'h798fb700;
    ram_cell[    2809] = 32'hf250ace0;
    ram_cell[    2810] = 32'h255b0583;
    ram_cell[    2811] = 32'hb8fa2ce3;
    ram_cell[    2812] = 32'h2d857d9a;
    ram_cell[    2813] = 32'h82f1aead;
    ram_cell[    2814] = 32'h442aecc7;
    ram_cell[    2815] = 32'h72f050cb;
    ram_cell[    2816] = 32'hab6573ce;
    ram_cell[    2817] = 32'ha763e94c;
    ram_cell[    2818] = 32'hd8eaec6f;
    ram_cell[    2819] = 32'h34b1929c;
    ram_cell[    2820] = 32'h3a409d1d;
    ram_cell[    2821] = 32'ha5bc7666;
    ram_cell[    2822] = 32'h1b7bd948;
    ram_cell[    2823] = 32'he17f7264;
    ram_cell[    2824] = 32'h3e700d68;
    ram_cell[    2825] = 32'h534a2831;
    ram_cell[    2826] = 32'h9c2a5ad4;
    ram_cell[    2827] = 32'h54aae4f9;
    ram_cell[    2828] = 32'h0d3fb56a;
    ram_cell[    2829] = 32'h63bae65c;
    ram_cell[    2830] = 32'h33f0854e;
    ram_cell[    2831] = 32'h0fe7231d;
    ram_cell[    2832] = 32'h0898e36a;
    ram_cell[    2833] = 32'h00bc7fdb;
    ram_cell[    2834] = 32'haca2cd6b;
    ram_cell[    2835] = 32'h996b5d2f;
    ram_cell[    2836] = 32'hb581d324;
    ram_cell[    2837] = 32'hec02b3ff;
    ram_cell[    2838] = 32'h795d4f1b;
    ram_cell[    2839] = 32'h478937c9;
    ram_cell[    2840] = 32'he7694112;
    ram_cell[    2841] = 32'hfe9c2abe;
    ram_cell[    2842] = 32'hd5bb6494;
    ram_cell[    2843] = 32'he70989ef;
    ram_cell[    2844] = 32'h962a578d;
    ram_cell[    2845] = 32'h6e4dfef3;
    ram_cell[    2846] = 32'h488b6899;
    ram_cell[    2847] = 32'hd14f4083;
    ram_cell[    2848] = 32'hbe1d9d03;
    ram_cell[    2849] = 32'ha6d275ea;
    ram_cell[    2850] = 32'h527e29b8;
    ram_cell[    2851] = 32'he4f82248;
    ram_cell[    2852] = 32'hfd1e4d97;
    ram_cell[    2853] = 32'h9677b91c;
    ram_cell[    2854] = 32'ha886b9b4;
    ram_cell[    2855] = 32'hb458db54;
    ram_cell[    2856] = 32'h662c0ac1;
    ram_cell[    2857] = 32'h1b726312;
    ram_cell[    2858] = 32'h7c164b50;
    ram_cell[    2859] = 32'h771781ed;
    ram_cell[    2860] = 32'hcdf8d531;
    ram_cell[    2861] = 32'h49bac06c;
    ram_cell[    2862] = 32'h21726fd3;
    ram_cell[    2863] = 32'h2ea3492f;
    ram_cell[    2864] = 32'h422e6a61;
    ram_cell[    2865] = 32'hdb6eabec;
    ram_cell[    2866] = 32'h92a4d93b;
    ram_cell[    2867] = 32'hb320ee63;
    ram_cell[    2868] = 32'hb1661e36;
    ram_cell[    2869] = 32'h314307b2;
    ram_cell[    2870] = 32'hcb4ddb85;
    ram_cell[    2871] = 32'h321955b4;
    ram_cell[    2872] = 32'h9dd97093;
    ram_cell[    2873] = 32'heb052e07;
    ram_cell[    2874] = 32'hf6c3431a;
    ram_cell[    2875] = 32'hfc0894f9;
    ram_cell[    2876] = 32'h331a1e73;
    ram_cell[    2877] = 32'hb1afcc8e;
    ram_cell[    2878] = 32'ha102a2fe;
    ram_cell[    2879] = 32'hf5a83d7b;
    ram_cell[    2880] = 32'h2cf41d7d;
    ram_cell[    2881] = 32'hb6acf262;
    ram_cell[    2882] = 32'ha1b34061;
    ram_cell[    2883] = 32'h691d2f78;
    ram_cell[    2884] = 32'hed9371f0;
    ram_cell[    2885] = 32'h5077c7cf;
    ram_cell[    2886] = 32'h50efd543;
    ram_cell[    2887] = 32'h1e69e37a;
    ram_cell[    2888] = 32'h1b3c0e89;
    ram_cell[    2889] = 32'h5a793a81;
    ram_cell[    2890] = 32'h9af0f683;
    ram_cell[    2891] = 32'h85166621;
    ram_cell[    2892] = 32'h4b6fb49e;
    ram_cell[    2893] = 32'h28ae61f8;
    ram_cell[    2894] = 32'hc8409bef;
    ram_cell[    2895] = 32'h928e13e4;
    ram_cell[    2896] = 32'h4931b9f0;
    ram_cell[    2897] = 32'h615b361c;
    ram_cell[    2898] = 32'h2af31f66;
    ram_cell[    2899] = 32'h33ad1bbc;
    ram_cell[    2900] = 32'h120b1328;
    ram_cell[    2901] = 32'h69e1b5e1;
    ram_cell[    2902] = 32'hceac2db4;
    ram_cell[    2903] = 32'hcf0abc8e;
    ram_cell[    2904] = 32'he6470d77;
    ram_cell[    2905] = 32'hf46745bf;
    ram_cell[    2906] = 32'hfe57e759;
    ram_cell[    2907] = 32'h3990d85d;
    ram_cell[    2908] = 32'h4bac9fe6;
    ram_cell[    2909] = 32'h114da3b7;
    ram_cell[    2910] = 32'hdc4e0a52;
    ram_cell[    2911] = 32'h27b8e55a;
    ram_cell[    2912] = 32'h478f4d53;
    ram_cell[    2913] = 32'h1711b4bf;
    ram_cell[    2914] = 32'hd85bccf9;
    ram_cell[    2915] = 32'hdb5f1121;
    ram_cell[    2916] = 32'h2cb06960;
    ram_cell[    2917] = 32'h6212cb76;
    ram_cell[    2918] = 32'h7bdb4030;
    ram_cell[    2919] = 32'h258ac099;
    ram_cell[    2920] = 32'h6a55b7b4;
    ram_cell[    2921] = 32'hcc5327a5;
    ram_cell[    2922] = 32'haec2ac8a;
    ram_cell[    2923] = 32'hdc6edabc;
    ram_cell[    2924] = 32'hdc4de14a;
    ram_cell[    2925] = 32'hf8338c2e;
    ram_cell[    2926] = 32'h8466c736;
    ram_cell[    2927] = 32'h6262c33c;
    ram_cell[    2928] = 32'he1588bbd;
    ram_cell[    2929] = 32'h18908122;
    ram_cell[    2930] = 32'hd02426b3;
    ram_cell[    2931] = 32'h3085be75;
    ram_cell[    2932] = 32'h755aabfb;
    ram_cell[    2933] = 32'h924628fc;
    ram_cell[    2934] = 32'h8ec8dfd3;
    ram_cell[    2935] = 32'h1cc8b6eb;
    ram_cell[    2936] = 32'h859234de;
    ram_cell[    2937] = 32'hf3037528;
    ram_cell[    2938] = 32'hc3f97f25;
    ram_cell[    2939] = 32'hd62c57fa;
    ram_cell[    2940] = 32'h1c7cdf5f;
    ram_cell[    2941] = 32'h8a2aa5d4;
    ram_cell[    2942] = 32'hac30e17d;
    ram_cell[    2943] = 32'h331322f7;
    ram_cell[    2944] = 32'hf4a8d6b0;
    ram_cell[    2945] = 32'h105ceb29;
    ram_cell[    2946] = 32'h5cf5030b;
    ram_cell[    2947] = 32'hff457371;
    ram_cell[    2948] = 32'h882764f4;
    ram_cell[    2949] = 32'he9c5d73c;
    ram_cell[    2950] = 32'hfc6ece26;
    ram_cell[    2951] = 32'h0d730a82;
    ram_cell[    2952] = 32'he34a3f48;
    ram_cell[    2953] = 32'hba6f7efd;
    ram_cell[    2954] = 32'h6f5bc988;
    ram_cell[    2955] = 32'h20ac4f5e;
    ram_cell[    2956] = 32'h38a47130;
    ram_cell[    2957] = 32'h60336782;
    ram_cell[    2958] = 32'h92820b84;
    ram_cell[    2959] = 32'ha9cb5af2;
    ram_cell[    2960] = 32'heb910dc7;
    ram_cell[    2961] = 32'h88406e6a;
    ram_cell[    2962] = 32'hd6dd1adf;
    ram_cell[    2963] = 32'h3062295f;
    ram_cell[    2964] = 32'hea802803;
    ram_cell[    2965] = 32'h77116ffc;
    ram_cell[    2966] = 32'ha127c637;
    ram_cell[    2967] = 32'h604f95ae;
    ram_cell[    2968] = 32'h0c272aaa;
    ram_cell[    2969] = 32'hac88e265;
    ram_cell[    2970] = 32'ha9bd3a72;
    ram_cell[    2971] = 32'h5fc67341;
    ram_cell[    2972] = 32'h8aeb512e;
    ram_cell[    2973] = 32'h5c77d446;
    ram_cell[    2974] = 32'hf253ed79;
    ram_cell[    2975] = 32'ha1fc7a57;
    ram_cell[    2976] = 32'ha60481ac;
    ram_cell[    2977] = 32'h448b6065;
    ram_cell[    2978] = 32'h0d55fa97;
    ram_cell[    2979] = 32'h365ed316;
    ram_cell[    2980] = 32'h269a441e;
    ram_cell[    2981] = 32'h359e4e34;
    ram_cell[    2982] = 32'h646285c3;
    ram_cell[    2983] = 32'h150e9234;
    ram_cell[    2984] = 32'h0bd1763e;
    ram_cell[    2985] = 32'h658b867e;
    ram_cell[    2986] = 32'hfae0dbd0;
    ram_cell[    2987] = 32'hfc9535fa;
    ram_cell[    2988] = 32'h2e9b85bf;
    ram_cell[    2989] = 32'h394ed199;
    ram_cell[    2990] = 32'ha0aab6a2;
    ram_cell[    2991] = 32'h5e2ac5ea;
    ram_cell[    2992] = 32'he9bce877;
    ram_cell[    2993] = 32'h1c2ea220;
    ram_cell[    2994] = 32'hcdb1bc9d;
    ram_cell[    2995] = 32'h7b2f5120;
    ram_cell[    2996] = 32'hee0aa163;
    ram_cell[    2997] = 32'h1eae2627;
    ram_cell[    2998] = 32'hbce822f2;
    ram_cell[    2999] = 32'h09e2a975;
    ram_cell[    3000] = 32'h092d45c6;
    ram_cell[    3001] = 32'h726f0e78;
    ram_cell[    3002] = 32'hbebee571;
    ram_cell[    3003] = 32'hef87e000;
    ram_cell[    3004] = 32'h2223007f;
    ram_cell[    3005] = 32'h6301d22b;
    ram_cell[    3006] = 32'h42d2614b;
    ram_cell[    3007] = 32'h40b5039d;
    ram_cell[    3008] = 32'h0fb12ca4;
    ram_cell[    3009] = 32'hd68432ff;
    ram_cell[    3010] = 32'h05af7005;
    ram_cell[    3011] = 32'h77e77dd4;
    ram_cell[    3012] = 32'h146b9278;
    ram_cell[    3013] = 32'h6b565b6c;
    ram_cell[    3014] = 32'hb66ebe43;
    ram_cell[    3015] = 32'h1fbf195f;
    ram_cell[    3016] = 32'hfa79e9d1;
    ram_cell[    3017] = 32'h849d0976;
    ram_cell[    3018] = 32'h744ce655;
    ram_cell[    3019] = 32'hba440075;
    ram_cell[    3020] = 32'h86c253d0;
    ram_cell[    3021] = 32'h60333c8c;
    ram_cell[    3022] = 32'hc7e7d574;
    ram_cell[    3023] = 32'h7eac1200;
    ram_cell[    3024] = 32'h6afda0b6;
    ram_cell[    3025] = 32'h3e030fe1;
    ram_cell[    3026] = 32'hb378da72;
    ram_cell[    3027] = 32'hb22184c0;
    ram_cell[    3028] = 32'he0fc98ac;
    ram_cell[    3029] = 32'hf3d2f127;
    ram_cell[    3030] = 32'h15d286f4;
    ram_cell[    3031] = 32'h07445cc2;
    ram_cell[    3032] = 32'h21062a96;
    ram_cell[    3033] = 32'hbd3a6bda;
    ram_cell[    3034] = 32'h16609c7b;
    ram_cell[    3035] = 32'h2dc67fcf;
    ram_cell[    3036] = 32'hae22b12d;
    ram_cell[    3037] = 32'hdf48447a;
    ram_cell[    3038] = 32'h3fb2f7a7;
    ram_cell[    3039] = 32'hdc3dc370;
    ram_cell[    3040] = 32'h5ac6e4b4;
    ram_cell[    3041] = 32'h7c2bb9bf;
    ram_cell[    3042] = 32'hf456b7ed;
    ram_cell[    3043] = 32'hcf183c28;
    ram_cell[    3044] = 32'h8828c707;
    ram_cell[    3045] = 32'h5490a964;
    ram_cell[    3046] = 32'hd0e30ed2;
    ram_cell[    3047] = 32'ha3a612fa;
    ram_cell[    3048] = 32'h39e61320;
    ram_cell[    3049] = 32'hd6eb3789;
    ram_cell[    3050] = 32'hc3d9e71e;
    ram_cell[    3051] = 32'h2b0c3162;
    ram_cell[    3052] = 32'h9c1e1a32;
    ram_cell[    3053] = 32'h22e59e81;
    ram_cell[    3054] = 32'h70a5cf47;
    ram_cell[    3055] = 32'hfc4282b4;
    ram_cell[    3056] = 32'h75959d48;
    ram_cell[    3057] = 32'h6ddbaec5;
    ram_cell[    3058] = 32'he6502487;
    ram_cell[    3059] = 32'h43cf3442;
    ram_cell[    3060] = 32'he59968e7;
    ram_cell[    3061] = 32'h80ddb3ab;
    ram_cell[    3062] = 32'h35a75384;
    ram_cell[    3063] = 32'h848b2619;
    ram_cell[    3064] = 32'h959c040b;
    ram_cell[    3065] = 32'h43f5219a;
    ram_cell[    3066] = 32'h7986da8c;
    ram_cell[    3067] = 32'hd593aef5;
    ram_cell[    3068] = 32'h45cf0931;
    ram_cell[    3069] = 32'h908d2661;
    ram_cell[    3070] = 32'hf4fafeae;
    ram_cell[    3071] = 32'h27f852c7;
end

endmodule


`timescale 1ns/100ps
//correct read result:
// 00003530 000026eb 000020d5 000033d8 00002082 00000fc1 00003a24 00000f46 00001637 000035da 0000121c 000016d9 00001fc2 00002bac 00001aeb 00002d7d 00001b08 00000251 000029d8 00002b1a 00000e19 00001bee 000008d4 00001274 00002416 00001678 00001ae3 000033e3 00000bf0 00001f8d 000011ae 00000f0a 00001948 00002cb6 000031ff 00000b89 00002b8e 00002797 00002cfe 00003090 00001bef 00003bf8 00002c87 00001328 00003c78 00000f5b 00002c91 000012c4 00000ae1 000019bc 000013f3 00001a35 00000c13 00001d2e 00001525 00000ee1 0000137d 00001caa 00003374 0000130e 00000e8c 0000026e 00002be5 00002e09 00000ebf 00003754 00001680 000020b4 000013a6 000029c8 00002c53 00000b56 00002c2c 000025f9 0000352b 000027a7 000027a8 0000293b 00003652 00001f3e 00001772 0000038b 00003af2 00003e3f 00001ee2 000039e6 00003061 00002026 00001406 0000233d 00000c7a 0000255f 0000261c 000023c8 00002b66 000010e9 000019d9 00000471 00001176 00000281 00002fed 000033cc 00000cb2 0000243b 00001cc4 00001d39 00001f10 00000ab8 000009a6 00001532 0000365b 00003932 00000959 00000706 00002b4a 000039f8 00000cc4 00002b50 00001dcc 000005fa 00002131 0000151e 00000cf7 00002ae7 00001692 0000155b 000029da 00003d50 000032b2 00002978 00003359 00002b52 00000fa7 00003c63 00000386 00002853 000023f3 00003540 00001875 000006af 000004a0 0000273b 00003363 00002fe7 00002155 0000221f 00003691 000000e3 00002101 00002e8e 00002f83 00003efa 0000028b 0000308c 00003307 00002e78 0000327b 0000344c 00002bf2 0000349e 00002d8f 00001485 00001d81 0000013d 0000039d 000007a7 00003b4e 00001e9c 0000289c 000006fd 00003bb9 000029e6 000032be 00003100 00002d04 00000c3f 00001088 00001df4 0000221e 000010cd 00001bde 00001353 00002c4f 0000343a 00002a1f 0000090f 00000e4a 00002bd1 00000102 00003603 00000ce6 000037ad 00001bf5 00000a18 000001e5 000002aa 00002a9d 000013b5 00000ee9 0000252d 00003419 00003341 00001dc4 00000a0a 0000373b 00000a4c 000010d4 00002d5d 0000168d 000014f2 0000342d 00003b29 000023c6 00000933 000007fd 0000068d 0000141e 00000624 000028e9 0000024a 00000855 00000d0c 0000002f 000030fc 00000640 00000188 00001bed 00001d15 00002c89 00002dda 000014a4 000025c9 00002b86 00003e1d 00001fe3 000016e5 00001689 000016fb 00002b45 00003033 00001406 0000396b 0000183c 00001500 0000322e 00000ac8 0000056a 00000b69 00003703 0000259f 0000083a 00001025 00001612 00002a7e 000038a0 000036d9 00000540 00001b94 00000ce5 0000171a 00000b0c 00002e1a 00000d1e 00003cbe 00003f5d 00000b88 00000a48 00002afb 00001ac4 00003378 00000e9b 00003553 000021c4 000023b8 00002dda 00001bc2 00002ce5 00001929 000010b4 00002654 000004d1 0000275d 00000858 0000352f 0000090f 00000ed4 00000eb7 00000752 000008ae 00001f18 00002a6e 00001f64 00003020 00003dd0 00000cbe 000009d6 0000112d 00002a6c 000019bf 000016f8 00002d1e 00003b56 00001da9 00003fe7 000034f8 00000cea 00001a9b 00002191 00003f92 000003c3 00003174 00002e86 00003eaf 00001ca4 00003c39 00002bcd 00001fc8 00002f3b 000010f4 00001e0e 00001ebc 000024d7 0000160b 00000f98 000020fe 000021d0 00003978 00001bdc 00001053 00002109 00003e49 000018dc 00000aee 000006ae 0000223d 00000a7c 0000288e 0000195b 00002366 000021cc 00000dfa 000015ea 00002c7f 00000dac 00002c7a 0000257e 0000059f 00002ec7 000015a0 00000182 00003bf0 0000166a 00001aa8 00000931 00001095 00002000 00000e18 00001911 000033e4 000021eb 00000b8f 00001ec2 000024b7 000032c5 00000c63 00002301 000011d3 00000917 0000365c 0000259d 00000e21 0000311c 000013ca 00001a83 00000203 00002c4b 00003ff8 00001efa 00000e76 00000276 00001bc2 00001026 00001785 00003750 00001c64 0000177d 00003b94 000014bf 00003ff3 00002d4d 0000216f 00003266 00002413 00002588 0000180e 00000470 00000eda 00000211 0000219f 00001deb 00002149 000037fb 00001705 00002a82 00001574 00002fc4 00002977 0000241c 00000d6c 00001673 000024eb 000009af 00000ea1 000025e7 00000735 0000179b 000003f4 00002fbd 00001656 00001041 000036f3 0000242b 00000631 00003257 00000521 0000010a 000009df 00001269 00001add 00000028 0000137c 00000e01 0000280b 00003986 00003e80 000033c8 00003166 00000510 00001f1f 00001946 0000137e 00003895 000030d7 000010a3 00002d73 00002a9e 00000c99 00000487 00000529 00003ef8 00000b82 000008a3 00000fa8 00001846 000007ca 00000b0f 00002a1d 00001d15 000037cd 00002288 00000a54 00002009 00000cf5 0000227d 000028a4 00000291 00003a89 00003734 00001ae0 00002766 00000a7f 000036df 00001c44 00002aed 00001de4 000038bb 00003493 00002c8d 00001597 00003622 00003323 000003a7 00002e30 00002512 00000316 000009d9 00002b52 00003b4c 00002db5 00000567 000017b3 000008f3 000031b1 000016b0 00002439 000010b7 00001834 00002917 000029c8 00002705 000030b4 00003050 00003920 00003b15 000033f7 000025e3 00001e01 00003612 00002de4 00002faf 00002a73 00003599 0000335f 000011b4 00003b58 000032f8 00003596 00002dce 000033a2 00000d6c 000021ae 0000190e 00000c2d 00001d2d 00001842 00000fb5 00002b8d 000008a1 0000298b 00001202 00003f31 000013c5 00002336 00002b99 00001623 000035e0 00003493 000000bb 00002958 00002baf 00002063 0000209c 00000761 00002b28 000022fa 00001100 000029d0 00000d30 00002170 000001bf 00000db1 00000f09 0000204f 0000328d 00003ba5 0000275a 00003126 00000613 000024ab 00000ba9 00001f2f 00001d1f 00003333 00002807 000033f5 000019eb 00002855 0000053f 000032d4 00000a4d 00002d83 000026e6 00000236 00000b50 0000119f 000036ec 000019ed 0000145b 00003527 00003452 00000da9 00003f8b 00002533 000008e2 00002689 000027d1 00003f08 00002a28 00003baa 0000260f 000002f5 00001a5b 0000072c 00003bc2 00001b63 00003bd1 00003415 000024b0 0000077d 00001593 00002b62 000037d5 00003753 00000b08 00003617 00003d64 000007b4 0000260a 0000000d 00002db5 00003c86 0000392a 00003cbc 00003161 00003be1 00002cb9 00000706 000027de 0000319a 000027a1 00002f21 0000070a 00000a3e 00001e6e 00002cd4 00000d1c 00001544 0000218e 00000299 00001eaf 00000b8d 00000264 00000f17 000027ea 00002cfe 000002d9 00000d4e 00002e54 00000ff8 000001fe 0000069a 00001f23 000007b9 00003a32 00000682 00000f0c 000001eb 00001f58 00002d31 00001cee 00003a3c 00002124 000029c7 0000151a 000022b0 000039b4 0000310c 00001694 00000b25 000027eb 000001ed 000032fc 000035c0 000037c7 00001a33 0000122e 00000942 00000645 00001030 000035e1 00001895 00003fb6 00002d1b 0000193c 00000d98 0000031f 000017f6 00000cdd 00001730 000006b2 00003382 00000eca 0000316b 00003e94 00001957 00002561 00003494 00003e4b 00000367 0000292b 00001899 0000189d 000035d4 000025c2 00002c71 0000257e 00001501 0000187d 00001690 0000181c 00001841 00002765 0000094f 00001a39 00002673 00003ebf 000010a1 000030e2 0000316f 0000364c 000010af 00001598 000006c7 00003781 00000bfa 00002a6e 00002c6c 000011fe 00003861 00003868 00002cb3 00002314 00003977 00000a0d 00000ea3 00002c3b 00001aa5 000003dc 000009b0 00000a4f 0000306c 00000097 0000104a 00000e53 000012e3 00003c1c 000011cd 0000169d 00002a5e 000037e4 00001f69 000024ff 00000355 00000e68 0000146c 00002ca7 0000273c 00002ca4 00002b21 00003b85 00002c6d 00002241 000020c2 0000179c 000009f4 00002ec7 000037a1 00002223 000038de 00000c9b 00003b3c 00002c16 00003e5b 00002a1b 00003ed0 00001764 000028e4 0000055e 00003db4 00001540 0000173d 000010b6 00000b46 0000232a 0000117e 00002649 0000035a 00001ae3 0000071c 000014cf 00000c6d 00000795 000014d9 00002956 000013f2 00001bd4 000030e3 000003e9 00003af7 000017cb 0000114e 00002b32 00002daa 00003712 0000279a 00000bc2 0000253b 00001a13 00002a7b 00003b83 00001808 00001acc 00003767 000012d7 00000402 00002880 00003345 0000003a 00003833 0000371b 00001149 000032e5 0000385f 00003c28 0000269a 00001524 0000209b 00002944 00002370 00001bc3 00003677 00003da4 00001f2a 00000f10 000026c4 00003ff8 00001410 00000acd 000031a9 000014a7 0000235b 000004a0 0000232a 00000d96 00000cbc 00000ec1 00003fb3 000004cf 00001d8a 00002e6c 00003cdb 00001fb4 0000344b 000008f8 0000245b 0000234a 00002846 00003cf8 0000389a 0000248d 00002e24 00000a3b 000003e3 000000ab 000035f1 000032e7 0000201e 00001a00 00000971 0000209c 0000109a 00002862 000027e6 00002a6b 000000f1 00003992 00002139 00002ac8 000012a7 00003014 00003995 00002468 000026ec 00002ee8 00002e13 00003b9f 00003b37 000002a5 00001c82 000000b5 00003d3b 000012b1 00000703 00000327 0000323d 00002cad 00003d9c 00003900 000028f9 00003757 00003f5e 000006d2 00000133 0000195f 00002beb 00002bfb 00003733 00000ba1 00001f9f 00002aa8 00000659 00001bd9 00001840 00001d71 00002685 00002c3a 00001217 000021cd 00003c06 00002881 0000111a 00003cca 00001d0a 00001ec5 000034d0 000033ac 0000196d 00003267 00002491 00002a81 000039f4 00002295 00003a7b 0000073a 000028f3 0000354b 00001749 00001d5a 0000348c 00000834 00000cd1 00001f44 00002dec 000019b3 0000301d 000036fc 000022dc 00001783 00002094 00000a6f 00003d9b 0000347b 0000034a 000004c9 000021eb 000010a5 00003706 00000056 00001441 000026ef 00001d6d 00001371 00001dad 000036d5 00003118 000039d2 00002357 0000337f 00000c5b 00003ba5 0000353b 00002dfe 00002f14 00003004 00002483 00002db4 000025c7 00003f9f 00000773 00003a1c 00001ed1 00001149 00003fea 00003f6e 00003686 00000206 00002b95 00000b83 000008cd 00003df5 0000158e 000005d9 0000392b 00000a67 00001260 000017fe 00003a2d 00001c18 00002f0a 000009e9 0000304d 00003a8f 000029ac 00000c42 00000a2e 000032b3 000013fb 00001ff0 00000973 00002b2c 00000d26 0000323a 00002581 00001aaa 00000138 00001134 00000f2a 00001c40 00003ec4 00003584 000037aa 00001db1 00001876 00003f05 00003526 000033e1 00000eb8 000011c3 00002ce5 00003f78 00002b25 000015df 000030ec 00002b40 00000760 00001941 00001fd4 00000165 000013ff 00001b8d 000002be 0000202f 000029cf 00003c9c 0000325c 00003fc6 0000268b 0000282f 000036d1 0000011b 000007db 00001854 00000dcb 00001bc0 000038aa 00003af5 0000203e 0000105d 00003491 0000306f 00001a5c 00002920 00001856 00001989 0000259a 000019da 00003f60 00003b52 00002949 000016d4 00002188 000012fa 0000348f 0000164c 0000381f 00001f95 000032ee 00003e20 00000e69 00001c21 0000006d 00001634 0000166a 00003a8e 00003738 00001946 00002d5f 00001963 000034c7 0000379b 000025bc 00001a5d 00003151 00001f91 00001d19 000027b3 0000362c 0000268e 000021f4 00002480 00003d3c 00001e53 0000242b 00000812 0000068f 0000184b 00000a21 00000cef 0000337e 0000170c 00003001 00003bfd 00002d68 0000109a 000014f6 00003ab9 0000074d 000029e4 00001466 00002ced 000010f5 00001fbf 00001d76 0000311a 000002d1 00003d65 00003e50 00003e03 00003e02 00000dd5 00003b4c 00001f86 000033a9 0000100a 00002986 00001963 00003f5a 00001c03 00003b5a 00000bf5 0000193c 00003755 00001137 0000178b 00002201 0000282d 00002366 000004b9 00001989 00003ee7 0000362b 00002115 00000cd8 00000a00 00001709 000024fe 00000b26 00003ceb 0000379b 00003414 00001599 00001e7d 00000dc5 00002eba 00002305 0000165f 00001a98 00001af0 00001d0e 00003aed 00002135 0000331f 00002d54 00003606 00002e73 00000673 00000f58 00001dc7 000003ae 00001cce 00003ecb 000031bc 0000226f 000006a8 00002ec1 00000a83 00003e5e 00003ba1 00000cdf 00003c30 00001534 0000274e 00002047 00002a8c 000016ea 00001cde 0000108b 000020d5 00001f3c 00002873 000008e7 00002dfb 00003495 00001888 0000150a 0000373d 00003b0c 00000965 000027e0 00001cb7 0000053d 00001a42 00003d36 0000131a 000003c6 0000371b 00002572 00002da5 000020cc 00003cd9 000020ea 000006ae 00000e85 0000114e 00001541 0000313d 00000e48 0000138b 0000131b 0000151a 00000552 00000227 00002daf 00001f7d 000034ee 00003361 0000296b 000010d5 000005a8 000017df 00003f76 000033c2 00003534 00000d16 00003497 00001697 00000aba 00000b0f 000023db 00000d84 000038ab 00003066 0000277b 000031bb 000015b5 00002ac4 00003758 000015bc 00001127 00000b8b 00001581 00003451 000036dc 00003901 000019b9 0000162b 0000346a 00002a61 00001448 00003eb1 00002c47 00001427 000007cd 00002b7c 000037db 00003d21 00000cf6 00001261 00001f03 000022ec 00003954 000034ed 00002683 00003a36 000039db 00001ca0 0000082b 000000a8 00002e56 0000121f 00000598 00002764 00001d8a 00002979 00001e89 00002590 00003ff5 00003fc3 00001a43 00001e7f 00002409 00003a77 00003114 000010ba 000010dc 00000b54 00003e28 000021ba 00001a18 0000164b 00001c5b 000007fa 00000553 000029c9 000012a3 0000144d 000006d9 00000951 000037c2 00002f15 00001be9 0000045b 00001eeb 000023a5 00003d52 00002500 00003561 000011c5 00000a37 00000066 00003abc 00000eb4 00001212 000007de 00001ca3 00001408 0000268e 00003637 00000c9f 00001a18 000030b3 00003cb5 0000099a 00000772 0000034d 000016b1 00003854 000006bc 000003ae 0000175a 00003285 000013df 00003b7f 00002e8d 00002ba3 00003bcf 00001b5c 00002100 00000e4f 00002062 000031c7 00003812 00002a54 00000e09 000039ec 000027c7 00000694 00002c07 00001888 00003c34 00002227 000004ec 0000179d 00002716 00002233 00003a7a 00001f07 00000387 000012f5 000021ba 00003067 0000204c 00003bdb 00001fa6 0000255e 00002679 000036f0 00002240 0000168a 000004c8 00003d06 00001d4c 00003e31 00000175 00003b3d 000008e4 000009c0 00000799 0000015f 00001fcd 0000110a 00003354 0000215b 00001efe 000026c0 0000003d 00003fa2 000019c8 0000157e 00001351 000015e4 00002a30 000004a6 00000607 000011b5 00001f48 0000004a 00003d31 00002e63 00002f24 000031d2 00001015 00000c28 000029d7 00002a06 00000bfe 00003178 0000295b 00002909 000027c3 00001c38 00000550 0000294d 00001130 000004c1 000015a3 000023e8 00003ee5 00002b0e 00000a0d 00001ded 00001822 00003e22 000028be 00000431 00001af7 000002f8 0000028b 00000b47 0000040e 00001f89 00001f6d 00003a6c 000033bc 00001fab 00000292 00003815 00001b12 00003ff7 00001199 00003f90 00002144 00001149 00001bca 00001eba 00003665 00000a5c 00001c1c 00003719 00001299 00003419 0000043f 00000cd4 000004a6 000008b8 000011c6 00001f26 00001e30 0000013d 000003ae 00001c3a 00000695 000030e1 00000cb9 00002f06 000032b9 000012f2 00002abc 00001311 000037b4 00001a53 0000230b 00001789 0000388e 00001cd7 0000295e 00003f06 00002a1a 00000713 000005e4 00003fb3 0000100a 00003d68 00000b72 00003a21 00002449 000031b3 000004fb 00002025 00000e19 00003d32 00001bec 000006f6 00001819 00000886 00003863 000003d0 00000878 0000253c 0000075a 0000253d 000020ce 00001902 0000220d 000033d2 0000168b 00003ae9 000001b0 00003d6e 00001864 000028d4 0000054d 00003f5b 00001cae 00001f48 00002f54 00000988 0000279d 0000399c 00001f8f 00001c31 000013f8 00002da5 00003926 00001cc9 000017eb 0000259c 00003ab1 00003cd4 000002c9 00000c3f 00003e78 00002984 00001b30 00003d0c 000027e2 00002f9a 000021a7 00000b5a 000004b5 0000057c 000022ec 00002d3c 00002cb6 00003f41 00002460 00000edf 0000086d 0000106a 000035e3 00003f18 00002c16 00002a71 00000ca0 000020a8 00003d55 00001d12 0000081c 00002df3 000022d9 0000088d 000009bd 00000a6c 00000442 000006cf 00002b4d 000003c6 000037a9 00000632 000001b9 00002d1e 00000e0f 00002cc7 0000383a 000037a0 000005e7 000012e6 000028e9 000006f2 000020f1 00002ddf 00002721 00001af3 00002104 00000be7 00002fce 00000523 00003967 00000644 00001c67 000031af 00001967 000010b9 00001777 000009a6 00001858 00001ad8 000016d5 0000050c 000009ed 00001ab3 000031b3 000004b6 000007f7 000036aa 00003989 00003867 0000090f 00003165 00003f1f 00002337 00002ba5 0000142b 0000217f 0000352d 000010e2 0000169c 00003b5b 00001813 00001a2f 000036ef 00002d7b 0000049e 00002978 0000175b 00001558 00002ee6 00000c50 00000422 000003cb 00002e79 00003406 00000579 000017d8 00002ad6 00002840 00003615 00000e22 000037fd 000010dd 000030a5 00001b69 00002e60 00001aa0 00000972 0000095f 00003d42 00002226 00002526 000032ce 0000338e 000015f6 00003219 000008b6 00003975 00000667 00003d6b 00000dde 00001d05 00003f11 00002d1d 0000201e 000002f1 000017a3 00003100 00001724 000034f1 00000cc1 00003407 000028fc 00002bff 00003d9d 000027d3 00000df1 00001408 0000289b 00002a29 000033be 00000236 00003aaa 00001254 00001591 0000078f 000003c1 0000038d 00001e53 000033ef 000000c0 00001bf7 00002bbd 0000397f 00000b97 00003fe1 00000129 00000680 00001db5 00002d72 00002990 000000ff 00002b22 00000de4 000020d0 000034d5 00003276 00000189 0000232e 00003ec4 0000385b 0000323f 00000edd 0000093f 00000a70 000034a8 00001cd6 00002e7d 00003570 00003b51 00000067 00000992 00001a02 000007e0 00000009 00000f17 0000324d 00000025 00000a5e 00000241 00002e68 00002110 0000064e 00003534 00001d06 000029d5 000037b6 000001af 0000041b 000023f8 00003632 000006e0 000028a3 00003ab2 00000db8 00002f99 00003cb0 000003a8 0000347e 00000724 000002ac 000007f9 00000d8e 0000080b 0000264e 00002e88 00003527 000004b2 00002731 0000211f 00002802 00000547 00003249 00003fa6 00003476 00000bb1 000002a1 00002598 000025b4 0000118b 00001318 00003007 00001fbf 000036f0 00002f0a 000015de 000002ec 0000365a 0000121a 00000625 000027a9 00002fc2 00003e94 00002ada 000036a9 0000308c 00002e75 00000def 00003aed 0000063e 00000e26 00002ea1 00000f83 00000e59 000039c3 00002385 00003f65 00000f00 00002bcb 00002e80 000015e1 000034bb 00000ee1 00003a13 00002cf4 00001dcc 00003afd 00001638 00003556 00003ca1 0000367c 00002b44 00002c70 00001f73 00000dda 00001088 00000441 00002d9d 000003be 00000b6c 00000b79 000015f7 00001d23 00001a8b 00001d46 00002684 00003882 000036af 00001dd1 00001131 0000213b 00001baf 00000b54 00001243 00001ca9 00001b41 00001536 00001638 00000a5a 00003b26 00002244 00000f8c 00003544 00001572 00001c4c 00003a79 00003859 000001f9 00000f49 000007bb 0000163b 00002e64 000020a9 00002616 00003678 00002df1 00000942 00001abd 000029e7 00001b85 00000ff4 000018f6 00002ee6 00000fcb 00002912 00003388 000009c4 00002ba9 0000347e 0000364c 000010d3 00000eb7 00001b9c 00003883 0000139c 00003eae 00002251 000020b8 000022bc 00001219 00003cc8 000032d0 00001677 000021fd 0000253d 000012b0 00001957 00000932 00003c9f 00000fc9 00001121 00000234 00000824 000036c9 00001f0c 0000349b 00003aab 00003ba6 00002ff9 00001314 00003b4c 00001340 00003028 00000cd7 00000acd 00001ca4 00001b0d 00000881 000026c3 00003a19 00003329 0000385f 00001523 00002963 00000ee0 00000791 00003ebf 00000bef 00000436 00003a7f 00001b27 000018fc 00003369 0000092d 0000315a 00000d37 00001a85 000036c2 00001ab8 00001157 00003157 00003f8e 000017fe 00003d25 00001dad 000021ef 00002c66 00003882 00000453 00003075 00000d3f 00001d4e 00001f55 00000ec0 00002535 000037d8 00003cb0 0000094a 0000283b 00001d4d 00000170 00001848 00003c6f 00003804 00003b64 000019ea 000019da 000006e7 00000eec 00001995 000032ab 000022ea 000016c9 00001e48 0000346d 000021d8 00001b44 000038ae 00002d6a 000030ef 0000032f 000002d5 00002cb3 000036fb 000009fb 000006ff 00000c26 0000212c 000035d2 0000000d 00003d02 000007b6 00003fdd 00001de6 00000faa 00002cb2 00002b28 0000232d 0000372a 0000127f 00002aa0 00000631 00003296 000035cb 00001734 00003f74 000034dc 00003060 00002d1d 0000330d 00001236 00003ef9 00001dde 000017f0 00003961 00002923 00003e6b 000030a0 0000087f 000033a9 00000789 00000441 00001d9d 00002511 00002b77 000023e1 00002757 000010d5 00000595 00003295 0000025d 0000037f 00002bab 000036a5 00001411 00001cdc 000038be 000030d9 00002a4f 000000f9 000028bc 000009df 00000f05 00000746 00002b23 00003442 0000307e 0000011b 00003e62 00001981 000004dc 00001858 000015a4 00002d00 00003afc 000030e3 0000207b 00001337 000024f9 00000fde 00003e84 0000202c 00002494 00001e2b 00003a9a 000002c1 00000f98 00001b62 00003b15 00001c35 000031f8 00002a0f 00000708 00000623 00000488 0000192e 00002dd6 00000209 00003b59 00001857 0000100e 00003eff 00000e11 000017f7 00000e58 00000649 00002c33 000029b4 00003b2c 000031e6 00002851 000038d5 000038e1 00001254 0000261b 00002c28 00000233 00000067 00001927 00000874 00003969 00000688 0000156c 00002993 00002c53 00000ec1 00000602 00000dce 0000305f 00003a3d 00003aea 00000fe5 0000130f 00001c6b 00002d8a 00001d8b 00001616 0000397b 00002b05 000023ca 0000366f 00001c91 000019ac 0000014f 00001478 00002d62 000027cd 00003d37 00002e7c 00001322 00001399 00002560 00000377 00002da8 00001adc 000013a5 000023b0 00000271 00001d75 00003777 0000325d 00002c20 000017b9 000022b7 000004a6 0000039d 00001e01 00002f44 00001ce0 000002e3 000014d0 000021b2 00003320 000013e7 00003ec6 00001f35 00001685 000017e7 00003595 00000f8b 000031ad 00003d3a 00002d20 0000231d 00003b22 0000291d 00001d6c 0000276a 000008ae 00000c37 00000bee 0000130c 00001552 00000584 0000193e 0000108e 000013f8 00001f6f 000032fb 000000b2 00000827 00000a98 00002bfe 0000037a 00000fb5 000035e0 00002878 00003a6f 00002acb 00000b3a 0000048d 000039b9 00001f5e 000015e4 000019de 000012ad 000025a5 00002797 00003a48 00003883 00000159 00003acb 00003cab 0000349e 00001647 0000335d 00001859 00000163 00001b38 0000224b 0000091e 000019a8 00003ec5 00003897 00000d24 00000bd9 00000a36 00001e16 00003d55 000017b1 0000221d 000000b0 00003fd4 000037f7 00003c4e 00002943 000021ec 00003571 000020ac 00002e80 00000ec4 0000065c 00001fcf 00000032 0000309d 00003f46 00002495 00000c8f 000027b2 0000238f 00000597 00000f54 00000e85 00003bbc 0000116f 00002bf9 000001dd 00003333 00003440 000016e9 00001251 000000f7 00003642 000018a1 00003604 000011d9 000031a3 00001dda 000037b1 00000d48 0000381b 00003689 00003059 000000a9 00001c5f 0000327a 0000064f 00003574 000021f5 0000372d 00003cf9 00000464 0000190c 00000235 0000260d 00001254 00000991 0000268d 000029b9 000034aa 000030f7 000000a3 0000030d 00003a99 00003156 000015e9 00003b4f 00002626 000020a5 000036be 00003266 00003145 0000241a 00000c06 000030da 00003b0e 00003f8e 00001fa5 00001133 00003d93 00003bcb 00002047 00001115 00001e57 00002d32 00001fd7 00001228 00000d16 0000282c 000009c4 0000277a 00003ee2 000003fe 00002991 0000129f 00003bc2 000011de 00000a05 00000638 000035d3 000034cc 00001cee 00000dc8 000035b5 0000144a 0000157a 00003e98 000031ba 0000229c 00002420 00002051 000005bf 00001a7c 00002a55 0000399b 00000976 00001417 00001b83 0000365d 00000083 00002b0b 0000216b 00002e2f 00000796 000029ad 00003ddf 00002b71 0000217e 00003d9e 000032f4 00000a9d 000016e9 00002bc8 00000188 00000714 000039f8 00000ec0 0000371b 0000050e 00000557 000009c8 00003a1e 000026a5 00002605 000020d6 0000066d 000027b0 0000110d 000005fc 00002968 000038c6 00001a91 000016f7 00000d42 00000625 00000686 00001454 000017eb 00001693 00003b9e 00003b20 00001e56 00001461 00002046 00000aa8 0000167f 00003fd8 00001c82 00003d73 000023d2 000010c7 000003d9 000021e4 00003594 00001969 00003188 00003a2e 00003272 00002223 00000563 000036c6 00000a9b 00000aa9 00000d02 0000348e 00000217 00003971 00001b32 0000349d 00003d5a 00001187 00001538 00001bd0 00000e11 00001604 00001be7 00002357 000011e4 00001bea 00002400 00003c0c 0000202e 00000dd0 00003381 00000418 000035f7 00002b6b 000020c8 00002db8 00002316 00001888 0000324f 000036e8 00002fed 000036c3 0000354b 00001e6f 00003742 00003fb7 000038f3 000003b7 00003b22 00001a07 0000115a 000033a8 000022e5 00003b13 00002142 000009d5 000006ff 000036b4 000010f9 00000484 000038f8 00002358 00001863 0000341d 00003200 00002a5a 0000057a 00001b9b 0000047c 000012e3 000015f3 00001587 00002b6a 00000a4b 00001ebd 00000f91 000038b7 000001be 0000318d 0000330f 000002cf 000012d5 00001c95 00003096 00001ee6 0000217a 0000018b 00000629 0000239f 00000a01 00000edc 00001832 000006dc 000023ff 000037e9 00003bba 0000114d 000014b6 000010d4 00002560 00003fc1 00000990 0000098c 000037fd 00000615 000036aa 0000107f 00000317 00000b02 00000167 00001c6f 000019cb 0000318a 00000005 0000382a 00001a73 000036e6 00002e6c 00003610 00001f6b 00002b1a 000021ca 00003a70 00002933 000012ea 000016eb 00001c82 00003808 000022ee 00001f2d 000008b3 00003231 000023de 000034d6 00003928 000039fe 0000053a 000021c7 0000186c 000022d0 00003816 0000191d 00001483 000037d9 00000a4d 00000cfa 0000260e 00003b8c 000032d2 000000f8 00003f5a 0000154a 00001e35 000017cf 0000073f 00001756 000007ff 00001302 00003eff 000029e1 00003416 00001bf2 000020c6 00002967 000014f1 000038cf 00003cb2 00003fec 00003c8b 0000109b 00001727 000013e9 0000052b 00001811 00001097 00001503 000011f0 000008b0 0000310f 0000166e 00002fbc 00002172 00000ce1 00000e55 00002b34 000000b6 00001056 00000133 00000e2f 00001792 00003546 00003a8d 000018e0 00003b86 00002f94 00003333 0000163c 000010d6 00002781 000039a5 0000337f 000027a3 000008f2 00003a8c 000025af 00001d76 000023d8 0000215b 00001a12 000036f9 00000ea0 00001e18 000029bb 00003ca3 00001f70 000006de 0000349d 000009fd 00003401 000024f0 00003f47 00003b76 000018fe 00003d9b 000038b7 000015a2 00001216 000033a0 00001ed0 000019e4 0000262c 000036c9 00003e86 00002c8e 00003277 000036b2 00002da6 000025ec 0000276f 00002f91 000008b6 00001cbf 00002381 000029cf 00000f9d 00003ab7 00001a8a 00003770 000029b3 00000a3e 00003250 0000362f 00000d7c 00003dee 000009b8 000022c3 00002bcd 000007f2 00000a8a 00000454 0000310e 00001a87 00000e61 000033de 00003fd2 00001cff 00003bf0 0000384f 00003997 000005a3 00002ffb 0000317c 00002771 00002343 000016bd 00001c89 00003b94 00003806 00001ea6 00001b7c 00000998 0000317d 00002b0a 00003b68 00003389 00001c79 000033f8 00002fef 000030fc 000028cb 0000024a 00002a48 00003fac 00002dad 00001077 000039bd 00002f47 00003ba5 00000c09 00003802 000031c2 000010e8 00001812 000002c9 00002aab 00000d65 00002ac6 000020f7 00001c57 000024bb 000015d3 0000286f 0000209b 00000698 00000a75 00001832 000000ff 000023ff 00002ea0 000018eb 0000013b 00003a50 000030cb 00001bd2 000001ae 00001673 000039bb 00001aeb 000030e5 0000383b 00002a0c 00003791 00000a9e 000033af 00003a41 000007ad 00003638 00002188 0000220d 000039a4 00001b14 00002636 0000107f 000032e8 0000181d 00003bb6 000024ad 0000182a 0000245f 0000022e 0000101b 00002974 00002d51 00002d76 00001ab8 000022a4 00000c2b 00000c36 00002bb8 000012e5 0000345f 00002447 0000364d 00000cca 00003e8e 00001e55 000023d9 00003ce1 00000bda 00002b71 00002595 00001037 000018ef 000014b0 00001565 00003b27 00002cf5 000011f0 00002b29 00000d72 000002c6 00001d75 00001cf0 00001114 0000366f 000031c3 000005c1 000007d4 00001238 000004a2 00001ad0 000023b6 00000bec 00002401 00002f6b 00002eab 0000243f 00001dbc 00002d0c 00002580 000001e0 000021a5 000034a3 00001383 0000219c 000032d4 00003b16 00002667 0000365c 00001745 00003ef1 00002095 00002c62 0000343c 00001fe6 00003778 00000704 0000187e 000002f6 000025e9 000018db 00002fd3 00003baa 00001a90 00001a3f 00003044 00002f31 0000223b 00000a55 00002040 0000312f 00001b31 00003532 000024f4 00003d65 00001a96 00003c9f 00001b82 0000008e 00002334 00000a6a 00000dd9 00002df3 0000315d 0000078b 00000b00 00000bba 000023fb 000035bf 00003ac4 000011b6 000014a3 000025f9 00003ef7 000016c0 000020f2 0000074b 0000231d 00000196 00003acf 00003d56 0000234b 0000002e 00002f8f 00000ae0 00001d20 0000395f 000025f2 00000aa1 00002eaf 00003a74 00000526 00001d15 000010d3 000025fe 00001da6 000010aa 00002b9c 0000040d 000011ca 000006a4 000015e1 00001939 00001a34 0000034f 000024c8 000026d7 0000120b 0000080e 00000ab9 0000363f 00001a55 00000c8b 000020e8 00000d3b 00001f10 000039f0 000022da 000014bf 00000215 0000025d 00000c9e 000020ee 00002593 0000212c 000013f4 00001193 00001f44 00003484 000014ba 00000894 00000be8 00003d18 0000288b 00003bc3 000039a3 0000021e 00003265 00003066 0000351f 000024ee 00002f3c 00003a2e 00000a06 00001914 000018f4 000011e9 00003c88 00000cb7 00001a74 00001f57 000024c4 0000358b 000024c3 00002618 00002bc6 0000204b 00002e40 00001587 000025d5 000008cb 00003451 00002b35 0000329c 00001a11 00003c5e 00001860 00001966 00001842 000035d7 00001902 0000399c 0000207b 000029ae 00000064 00003d6d 00002bc6 00001710 00003ad8 000001bb 000001a7 0000222d 000031cb 0000255a 0000324f 00002f30 0000098d 00003213 00001e27 00002883 00003dd2 00003546 00001513 000035c8 00001be3 00002f50 000015d9 00001a1b 00003762 000009db 00001604 000011b2 000000fc 00003559 00002815 00000e09 00001a1d 00003248 000038ea 00002c2d 00003f72 0000059b 00003157 00003d30 000015ff 00003fa9 000002b2 0000178b 000006b8 000001af 00000475 000010db 00002874 00001b76 000012ac 00002bde 000017fc 00001573 00002219 000009ce 00000452 0000040b 00002b0a 00002cbf 00001a13 000013cf 00000674 0000227a 00001a25 00000a00 00001a3c 000000e3 00003d1a 00000ef0 00003800 000020d7 00003c39 0000016e 00003662 00000e76 00002a17 00000271 00000386 00002a08 000017b9 000007a0 000006f9 000006ac 00002c38 00003531 000022e3 00002a8d 0000377c 00000003 00002645 00002941 00002b68 00000823 00000cc9 00002fac 00001e2c 00001191 00003716 00001707 0000145a 00003d3b 000027e7 00001658 000012d4 000013e0 000017cf 00003ca3 000026de 00002064 00001648 0000171d 000001b2 00001069 00000f19 00000d76 00000c92 0000070a 00000c09 00001b88 00001844 0000221e 00000fa5 00003d48 000000d9 00003fe9 0000072f 000029f6 00000eec 000011ff 000006f9 000006a6 000017a9 00001f7e 00003e71 00000d01 000015dc 00002ff4 000013be 00003465 00001349 00003d3c 00003cb5 00000ea0 0000226d 00002a50 000038a7 00001070 000020d8 00000525 0000124d 00002247 000009c4 000037d4 0000275b 00000611 00000303 000026df 00003ea0 00002cdf 0000000f 00000fa8 00002ab6 00001ae8 0000071f 000019a0 00002df6 000028c1 000009d0 00000b27 0000362d 000017c7 000006a3 00002bd7 00003481 00001702 000015fe 00001db5 00003ea2 0000103d 000017ad 00001cd2 00001f4b 00000eed 000031eb 0000287e 00000d4e 000015ee 000006cc 00002b5d 00000783 000013f5 0000162b 000013f6 00000daf 00001fa5 000017ca 00001e4f 000015a7 00001a57 000012fe 0000117b 00003aae 00000e3f 00000a83 00001622 000013d7 000018a5 00000a56 000028e8 00003e2a 000004e2 00002996 00002306 00003476 00002c62 000029ca 00002008 000006f2 00000a4b 00003ee7 00001a3d 00001997 00002e9f 00001370 000026ff 000012e3 000017ef 000012c8 000035ef 00003a61 00002550 00003271 000023d2 000039c8 000038f3 000012bd 000016b8 000005a5 000021e3 00003c8e 00003151 0000214d 00001c9d 00003f31 0000345e 000027c7 00003883 000009a6 00001d3d 00000f6e 00000c9e 00000e0d 00002c0e 0000279f 00002232 0000296c 00001dd8 00001c78 00003b66 00001a87 00003a00 00000f23 00000776 00000d6a 00000775 00000431 00001046 00003bd7 00003c1e 00002be9 00000203 00003a03 00002c53 00000cba 0000146a 00003d8d 00001091 00003302 00003941 00002818 00001aa2 000001ec 00000e08 00003c8f 00001dbd 0000275f 00003b0f 00000889 000035d6 00002484 00000370 0000266f 00003596 0000114b 000005e8 000027fa 00002178 0000174a 000020bd 00003cde 00000f2d 000013d0 00000202 00002f9f 00002040 00001ebe 00000f19 00002a1f 0000209d 000003a5 00003832 0000336a 000035ed 0000352e 000034aa 000017d7 00000bba 000000fd 00001fe7 00002abb 0000397c 00003177 0000165d 00001a05 00000ddd 00002fca 00002dd5 00002026 000009fc 000002bc 00000e58 00000768 00001f9b 000013aa 000012ba 000001cd 00002caf 00003707 000037de 000026ba 000036a8 00002b04 00002e70 000017f1 0000389a 00001303 000030b2 00002488 0000256e 00002a60 00003ccd 000037b9 000032a0 00000788 000023b5 00001b01 0000258c 00002d94 00003d68 00001f1a 000034f9 000023c2 00001914 000028d4 00000f6d 00000081 00001d04 00000cb1 000013ff 000005e1 00002b8b 00002acc 000003d9 00000fb7 000003f7 00000f6e 00000af5 00003ea5 000020bd 00003fbc 00002f5a 0000094c 00000b32 00002195 0000359c 00002a00 0000092d 00002df8 000007d9 00003342 00002e55 00000919 00000b7d 0000253f 00001010 00003ef9 00003421 0000290e 0000355d 00002cde 000027c2 00002f21 00002c61 00001cd9 000030b6 000026bb 00001199 0000037a 00001abf 000001ed 00003660 00003639 00002c4e 00001f15 0000149f 000006cd 00000245 00002a0c 000037be 0000134b 00000a60 00002590 000027da 0000111e 000017f2 00001bab 00000cb4 00001db8 00003937 00003323 00003b9c 00001dab 00003a8d 00001182 00001b0e 000032f1 00002e25 00000529 00002f5a 00000c0a 00002bf3 00001216 000026c5 00003320 00001dec 00002a4c 00003868 0000274c 0000158d 00003025 00003557 00003740 000033f0 00000b6a 000004c6 000027d5 000005ff 00001fb8 00001510 00003800 00002f57 00003be2 0000303f 00003bc2 000000fb 00000cb7 00000bd6 00002fe8 00003133 000013d1 00000e89 000023ae 00000f99 000032d4 0000239c 00002e69 00001704 00003732 00002128 00003752 00002100 00001e3a 00000d1a 00000662 0000185c 00000103 00001211 00000bb4 00000cdc 000023d9 00003cf3 000003f5 000022b4 00001147 00001789 00002428 00001bb0 0000236d 00000aa5 00000788 00002f94 00000597 00001891 00002611 0000118e 00002e6f 0000075c 0000052b 00002ad8 00003311 00002a67 00001b4f 0000372f 00001c5e 00001c7c 00002625 00000121 00001ca5 000015cd 00001266 0000024f 00003941 00002f1c 00000a48 000036e8 00002f45 00001a83 0000002b 00003677 00000ff5 0000121e 000017b9 00000fbd 000017de 00002eec 00000274 0000369f 00003be0 00003019 0000071d 00001d03 00000a3b 00001980 0000031c 00002b54 00003f9d 000002c1 00003db3 00002b51 00000ce3 00001200 00000515 00003448 00003510 0000011b 00002dd6 000010de 00002382 00003044 000005a2 00002985 00002916 000032a3 0000194b 000008ef 000026c4 00001fb3 000018d5 00003ebc 000001f3 00002f19 00000f1b 0000080f 00002cdc 000023df 00000cc6 00003b45 00000dcb 000005d7 00003406 00000218 00000928 00001e7f 000036fb 00003e16 00003af4 0000132e 00000c77 00003772 0000095b 00002b56 0000378a 0000395b 00000aad 0000305c 00000670 00001136 00002073 00000372 0000246a 00001509 00000f22 00000362 00003841 0000227f 00002b00 00003bab 0000328a 00002dd8 00002c10 000015c7 000013b9 00000393 00003b9d 00002702 00001276 000029b5 0000265b 000021c4 000021b8 00003a2a 00003baf 00000f4c 00002832 000015b5 00000637 00000f4c 00002d5d 00001663 0000252b 00001762 00002de4 00001cd4 00001a13 00002c45 00001c06 000039db 0000102c 00001f5d 0000334f 000036e0 00002a17 00000ef3 0000043b 00002b36 000021ba 000005ec 000016e0 00002b4b 000008c2 000007f3 0000154b 000029ae 000034ab 00001e32 000025cf 00000120 0000025d 00000706 00002218 00002404 00001951 0000206c 000010d2 00002ddd 00002040 00001786 000006e2 00000ae2 000006e6 00000b7c 00000ecc 0000045a 0000253e 0000011d 0000232d 0000150e 0000370f 00001290 000018ac 00003397 00001365 00000237 00002769 00000f45 000035dd 0000202e 0000003a 0000291b 00000a41 00001aad 00002373 00000e93 00000e3e 000004ff 00000ad9 0000246c 000037d3 00002d00 00001ac4 000017e2 00002428 00000656 00000df7 0000021f 00000106 00001cd0 000005e2 00000434 00003f5f 00002142 00001183 00003ed2 000003fa 00003c09 0000176a 00003717 000034f6 0000342a 00000358 00001c38 00003e55 000005fe 0000199f 0000057c 0000103b 000021c7 00003c6f 000028c0 0000066d 000003c6 00003b2d 00003fdd 00003d51 00001c09 000028bb 0000000c 00001381 00003f17 00003528 00000be2 00003d4f 00002b03 00002ab6 00001e4c 00000621 00003ac3 00001e05 0000161a 000004b7 00000e67 0000130a 00003a8d 00000d73 00000653 00002813 00003e9c 00001ec0 00002d97 000025ae 00000054 00002fe3 00003974 00001c9b 000003da 000019fa 0000226b 00002f27 000007f7 00000b91 000012ff 000031d0 00001f6a 00003270 000008b5 00002714 00002480 00002ed9 000014b9 00003283 00002eb7 0000260d 00000394 00001d0c 00002913 00001323 00000c25 00001552 00003dd8 00001ec5 00000948 000030e4 00003636 00003294 000032e7 000033d8 00000b77 00002a67 00003185 00001394 00000d62 000007dc 000022bb 00000845 0000261a 00003846 00001a06 0000341a 00000f3d 00001ebb 00001b14 00002dd0 00002c1b 00003054 00001b85 000020df 00002b10 000016d3 00002035 00002196 00000963 000016aa 00000640 00003425 00001c38 00002b8e 00001452 00001686 00000a71 00003dec 00003870 00000029 000000c1 00002675 00000666 00001eba 0000127c 00001f23 00000af1 000001b0 0000040a 00002fce 00003ee3 00000dcb 00000079 00000cd0 00002a18 00001ca5 00001875 000005fc 000007a6 00002ae5 0000232a 00001e12 0000166f 000023f5 00000928 0000165d 00003302 00000a58 00001368 000012ff 00003213 000023f4 00002556 00001582 00003eb2 00002a33 00003c86 00000d55 00003489 00002af2 0000065a 00001935 00003536 00003512 00001f35 000030b1 00001e82 000022c6 00002218 00000f3b 00003b5f 00002107 00003fb6 000031f2 00000c49 00000737 00002ffc 00001d65 00003fd9 00003ca1 00002918 00001be8 00000bd2 00000c75 00002967 00001c3a 0000090a 00000684 000034a1 0000012a 00003ddf 000000fa 00001b6e 000022bf 00002912 000023aa 00000061 00002a28 000014c0 00001177 00002580 00002d9b 00003f13 00002108 00000a19 0000094f 00000ec7 00001404 00001914 00001389 000003aa 00000117 0000113d 000016ba 00000893 000038c0 0000050c 000037ad 0000061c 0000076a 000009e7 00003491 00000fda 00003316 00002426 00003e01 0000176f 00003b6d 00003a09 00003908 00000a25 000006b9 00002d7f 0000351c 00000d70 00000625 00003f3b 000002dd 000020e1 00000694 000000cc 00000ed9 0000322d 0000123c 00000e06 000033dc 000039a2 00002ae9 00000fb6 00000a34 00000ba7 00002805 00002623 000020fd 000028cd 000014d9 000007d1 000025e5 00002b97 000038dd 00001999 00000273 000031c2 000027ad 000010cf 00000323 00001d52 00002947 000033fc 00002f12 000011b4 000027de 00002b5f 00003550 00002126 00002024 00000263 000025be 00003995 00000f7e 00000d3c 0000244e 000010ba 000030c2 00002928 000036c1 0000388a 00000bbc 0000138e 00000136 0000228a 000008f4 00001ae6 0000354c 00003bf1 0000147c 000025fc 00001bd3 00003c1c 00001f7b 00003ac2 00003e83 00000d1c 00003b99 00000318 000024c7 0000268d 0000059e 00000a5c 00000a9c 00001790 0000021b 0000263d 00001ae1 000015ff 0000272f 0000375e 00000e77 0000347d 00002784 000015a5 00003731 00000fb9 00002008 000003c5 00003f29 00001dfc 000011c4 00003717 00001e1b 0000248e 00000e46 000029e4 000037b1 0000340d 00002f27 0000155c 000039f2 00000bcc 0000318d 00003c88 0000376b 00000cb5 00003eba 00000238 00002353 00003fb5 00001030 00001798 00001d39 00001d12 00001b27 00001b38 000023de 000020e2 00002c60 000034d6 000015a2 00000596 000037ab 000011ef 00002f24 00003e87 00001eb0 00002651 00000f1e 00003008 00000166 00002344 00003af6 000037e0 00001b71 00002e6e 00000863 00003022 00002e31 00003cf7 00001762 0000220a 00003ef7 000015a4 0000070e 0000292a 00003d4b 00002eba 0000127e 00000f03 00002c7b 000014c8 00000cb0 0000321e 0000075c 00000f16 000027fe 00003dd5 000031b4 0000140d 00000932 000038b5 00003cfb 00000a82 0000146d 00003965 000016cf 000000fc 00000211 00002583 00003dee 00001192 0000162b 00002696 00002e4d 00000685 00002cbd 00001065 00002f3f 00003798 000034d5 00001350 00002461 00002593 00003ac3 00001362 000036c3 00001e4f 000034d3 00001cc8 00001884 00000d20 0000105d 00000ee7 0000070b 000035a5 000009ce 00003e0e 00001f7f 00000d7b 00001a1f 000033ed

module cache_tb();

`define DATA_COUNT (4096)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 4096 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000144;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h000026eb;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h00000478;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h000026ec;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h00001206;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h00002b82;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h0000143c;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h000024ef;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h00001637;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h00001b28;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h0000121c;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h000016d9;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h000030d7;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h000013be;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h00000895;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h000012ca;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h00001b08;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h00000251;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h0000297f;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h000016f1;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h00002001;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h00001cc5;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h000008d4;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h00002e0b;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h00002416;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h00001678;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h00000077;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h00000838;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h000003a2;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h000037f4;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h0000373c;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h00003961;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h0000229f;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h00001d6f;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h00000bbe;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h00000b89;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h0000187d;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h0000326b;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h00002cfe;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h00003090;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h00001bef;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h0000063a;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h00000266;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h00001328;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h00003ca1;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h00002f09;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h000034df;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h00002255;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h00002751;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h000019bc;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h0000174b;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h00002da2;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h00000bfb;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h000012fa;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h00001525;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h000026ef;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h0000137d;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h00003687;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h00003374;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h000026f2;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h00000529;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h00001abe;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h0000359b;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h00002ee2;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h00000d6c;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h00003754;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h0000165e;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h000020b4;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h00001d48;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h00001c0b;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h000039e7;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h00000b56;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h00002c2c;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h00001aa1;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h0000352b;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h00003580;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h000027a8;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h0000293b;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h00000cfe;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h00001b6f;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h00001772;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h000007b1;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h00003af2;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h00003e8c;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h00001ee2;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h00001795;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h000006ee;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h000002f9;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h000020d1;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h00001f59;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h00003b21;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h0000255f;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h00003319;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h0000339f;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h00002b66;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h0000148d;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h00000aaf;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h00001a30;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h00003145;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h00002c21;
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h00000190;  wr_data_rom[  100]='h00002fed;
    rd_cycle[  101] = 1'b0;  wr_cycle[  101] = 1'b1;  addr_rom[  101]='h00000194;  wr_data_rom[  101]='h00003c58;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h00000198;  wr_data_rom[  102]='h00003679;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h0000019c;  wr_data_rom[  103]='h0000082e;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000001a0;  wr_data_rom[  104]='h000022ff;
    rd_cycle[  105] = 1'b0;  wr_cycle[  105] = 1'b1;  addr_rom[  105]='h000001a4;  wr_data_rom[  105]='h00001d39;
    rd_cycle[  106] = 1'b0;  wr_cycle[  106] = 1'b1;  addr_rom[  106]='h000001a8;  wr_data_rom[  106]='h000007be;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h000001ac;  wr_data_rom[  107]='h00002a2e;
    rd_cycle[  108] = 1'b0;  wr_cycle[  108] = 1'b1;  addr_rom[  108]='h000001b0;  wr_data_rom[  108]='h00000411;
    rd_cycle[  109] = 1'b0;  wr_cycle[  109] = 1'b1;  addr_rom[  109]='h000001b4;  wr_data_rom[  109]='h00001532;
    rd_cycle[  110] = 1'b0;  wr_cycle[  110] = 1'b1;  addr_rom[  110]='h000001b8;  wr_data_rom[  110]='h00000e32;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h000001bc;  wr_data_rom[  111]='h00003932;
    rd_cycle[  112] = 1'b0;  wr_cycle[  112] = 1'b1;  addr_rom[  112]='h000001c0;  wr_data_rom[  112]='h00000959;
    rd_cycle[  113] = 1'b0;  wr_cycle[  113] = 1'b1;  addr_rom[  113]='h000001c4;  wr_data_rom[  113]='h00003d82;
    rd_cycle[  114] = 1'b0;  wr_cycle[  114] = 1'b1;  addr_rom[  114]='h000001c8;  wr_data_rom[  114]='h00002b4a;
    rd_cycle[  115] = 1'b0;  wr_cycle[  115] = 1'b1;  addr_rom[  115]='h000001cc;  wr_data_rom[  115]='h00003ee8;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h000001d0;  wr_data_rom[  116]='h00002041;
    rd_cycle[  117] = 1'b0;  wr_cycle[  117] = 1'b1;  addr_rom[  117]='h000001d4;  wr_data_rom[  117]='h00002b50;
    rd_cycle[  118] = 1'b0;  wr_cycle[  118] = 1'b1;  addr_rom[  118]='h000001d8;  wr_data_rom[  118]='h00001451;
    rd_cycle[  119] = 1'b0;  wr_cycle[  119] = 1'b1;  addr_rom[  119]='h000001dc;  wr_data_rom[  119]='h000005fa;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h000001e0;  wr_data_rom[  120]='h00002131;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h000001e4;  wr_data_rom[  121]='h0000350a;
    rd_cycle[  122] = 1'b0;  wr_cycle[  122] = 1'b1;  addr_rom[  122]='h000001e8;  wr_data_rom[  122]='h000032d5;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h000001ec;  wr_data_rom[  123]='h00002cee;
    rd_cycle[  124] = 1'b0;  wr_cycle[  124] = 1'b1;  addr_rom[  124]='h000001f0;  wr_data_rom[  124]='h000021bf;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000001f4;  wr_data_rom[  125]='h00003be9;
    rd_cycle[  126] = 1'b0;  wr_cycle[  126] = 1'b1;  addr_rom[  126]='h000001f8;  wr_data_rom[  126]='h000003b2;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h000001fc;  wr_data_rom[  127]='h000006be;
    rd_cycle[  128] = 1'b0;  wr_cycle[  128] = 1'b1;  addr_rom[  128]='h00000200;  wr_data_rom[  128]='h00000eb9;
    rd_cycle[  129] = 1'b0;  wr_cycle[  129] = 1'b1;  addr_rom[  129]='h00000204;  wr_data_rom[  129]='h00001d7f;
    rd_cycle[  130] = 1'b0;  wr_cycle[  130] = 1'b1;  addr_rom[  130]='h00000208;  wr_data_rom[  130]='h0000077f;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h0000020c;  wr_data_rom[  131]='h00002b52;
    rd_cycle[  132] = 1'b0;  wr_cycle[  132] = 1'b1;  addr_rom[  132]='h00000210;  wr_data_rom[  132]='h00000193;
    rd_cycle[  133] = 1'b0;  wr_cycle[  133] = 1'b1;  addr_rom[  133]='h00000214;  wr_data_rom[  133]='h00002a5c;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h00000218;  wr_data_rom[  134]='h00000386;
    rd_cycle[  135] = 1'b0;  wr_cycle[  135] = 1'b1;  addr_rom[  135]='h0000021c;  wr_data_rom[  135]='h00002853;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h00000220;  wr_data_rom[  136]='h000039ed;
    rd_cycle[  137] = 1'b0;  wr_cycle[  137] = 1'b1;  addr_rom[  137]='h00000224;  wr_data_rom[  137]='h00003540;
    rd_cycle[  138] = 1'b0;  wr_cycle[  138] = 1'b1;  addr_rom[  138]='h00000228;  wr_data_rom[  138]='h00002fad;
    rd_cycle[  139] = 1'b0;  wr_cycle[  139] = 1'b1;  addr_rom[  139]='h0000022c;  wr_data_rom[  139]='h00001e08;
    rd_cycle[  140] = 1'b0;  wr_cycle[  140] = 1'b1;  addr_rom[  140]='h00000230;  wr_data_rom[  140]='h00002a61;
    rd_cycle[  141] = 1'b0;  wr_cycle[  141] = 1'b1;  addr_rom[  141]='h00000234;  wr_data_rom[  141]='h000030df;
    rd_cycle[  142] = 1'b0;  wr_cycle[  142] = 1'b1;  addr_rom[  142]='h00000238;  wr_data_rom[  142]='h00001c38;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h0000023c;  wr_data_rom[  143]='h00002fe7;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h00000240;  wr_data_rom[  144]='h00002155;
    rd_cycle[  145] = 1'b0;  wr_cycle[  145] = 1'b1;  addr_rom[  145]='h00000244;  wr_data_rom[  145]='h00003b9d;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h00000248;  wr_data_rom[  146]='h00000c04;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h0000024c;  wr_data_rom[  147]='h000007b7;
    rd_cycle[  148] = 1'b0;  wr_cycle[  148] = 1'b1;  addr_rom[  148]='h00000250;  wr_data_rom[  148]='h000034b5;
    rd_cycle[  149] = 1'b0;  wr_cycle[  149] = 1'b1;  addr_rom[  149]='h00000254;  wr_data_rom[  149]='h00000c25;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000258;  wr_data_rom[  150]='h00002cf2;
    rd_cycle[  151] = 1'b0;  wr_cycle[  151] = 1'b1;  addr_rom[  151]='h0000025c;  wr_data_rom[  151]='h00002517;
    rd_cycle[  152] = 1'b0;  wr_cycle[  152] = 1'b1;  addr_rom[  152]='h00000260;  wr_data_rom[  152]='h0000188a;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h00000264;  wr_data_rom[  153]='h00000faa;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000268;  wr_data_rom[  154]='h00003307;
    rd_cycle[  155] = 1'b0;  wr_cycle[  155] = 1'b1;  addr_rom[  155]='h0000026c;  wr_data_rom[  155]='h000029ea;
    rd_cycle[  156] = 1'b0;  wr_cycle[  156] = 1'b1;  addr_rom[  156]='h00000270;  wr_data_rom[  156]='h0000342f;
    rd_cycle[  157] = 1'b0;  wr_cycle[  157] = 1'b1;  addr_rom[  157]='h00000274;  wr_data_rom[  157]='h00002e91;
    rd_cycle[  158] = 1'b0;  wr_cycle[  158] = 1'b1;  addr_rom[  158]='h00000278;  wr_data_rom[  158]='h00003c56;
    rd_cycle[  159] = 1'b0;  wr_cycle[  159] = 1'b1;  addr_rom[  159]='h0000027c;  wr_data_rom[  159]='h0000349e;
    rd_cycle[  160] = 1'b0;  wr_cycle[  160] = 1'b1;  addr_rom[  160]='h00000280;  wr_data_rom[  160]='h0000195b;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h00000284;  wr_data_rom[  161]='h0000142d;
    rd_cycle[  162] = 1'b0;  wr_cycle[  162] = 1'b1;  addr_rom[  162]='h00000288;  wr_data_rom[  162]='h00003399;
    rd_cycle[  163] = 1'b0;  wr_cycle[  163] = 1'b1;  addr_rom[  163]='h0000028c;  wr_data_rom[  163]='h00001c3a;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000290;  wr_data_rom[  164]='h0000039d;
    rd_cycle[  165] = 1'b0;  wr_cycle[  165] = 1'b1;  addr_rom[  165]='h00000294;  wr_data_rom[  165]='h0000381e;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h00000298;  wr_data_rom[  166]='h00000507;
    rd_cycle[  167] = 1'b0;  wr_cycle[  167] = 1'b1;  addr_rom[  167]='h0000029c;  wr_data_rom[  167]='h00001e9c;
    rd_cycle[  168] = 1'b0;  wr_cycle[  168] = 1'b1;  addr_rom[  168]='h000002a0;  wr_data_rom[  168]='h00003bbe;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h000002a4;  wr_data_rom[  169]='h00000fa6;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h000002a8;  wr_data_rom[  170]='h00003bb9;
    rd_cycle[  171] = 1'b0;  wr_cycle[  171] = 1'b1;  addr_rom[  171]='h000002ac;  wr_data_rom[  171]='h000029e6;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000002b0;  wr_data_rom[  172]='h000008f5;
    rd_cycle[  173] = 1'b0;  wr_cycle[  173] = 1'b1;  addr_rom[  173]='h000002b4;  wr_data_rom[  173]='h00003100;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h000002b8;  wr_data_rom[  174]='h00001340;
    rd_cycle[  175] = 1'b0;  wr_cycle[  175] = 1'b1;  addr_rom[  175]='h000002bc;  wr_data_rom[  175]='h00002e81;
    rd_cycle[  176] = 1'b0;  wr_cycle[  176] = 1'b1;  addr_rom[  176]='h000002c0;  wr_data_rom[  176]='h00000022;
    rd_cycle[  177] = 1'b0;  wr_cycle[  177] = 1'b1;  addr_rom[  177]='h000002c4;  wr_data_rom[  177]='h00001398;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h000002c8;  wr_data_rom[  178]='h00001ef8;
    rd_cycle[  179] = 1'b0;  wr_cycle[  179] = 1'b1;  addr_rom[  179]='h000002cc;  wr_data_rom[  179]='h00000598;
    rd_cycle[  180] = 1'b0;  wr_cycle[  180] = 1'b1;  addr_rom[  180]='h000002d0;  wr_data_rom[  180]='h00001904;
    rd_cycle[  181] = 1'b0;  wr_cycle[  181] = 1'b1;  addr_rom[  181]='h000002d4;  wr_data_rom[  181]='h00001353;
    rd_cycle[  182] = 1'b0;  wr_cycle[  182] = 1'b1;  addr_rom[  182]='h000002d8;  wr_data_rom[  182]='h00002c4f;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h000002dc;  wr_data_rom[  183]='h000018e8;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000002e0;  wr_data_rom[  184]='h00003cf8;
    rd_cycle[  185] = 1'b0;  wr_cycle[  185] = 1'b1;  addr_rom[  185]='h000002e4;  wr_data_rom[  185]='h000039e6;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h000002e8;  wr_data_rom[  186]='h00000e4a;
    rd_cycle[  187] = 1'b0;  wr_cycle[  187] = 1'b1;  addr_rom[  187]='h000002ec;  wr_data_rom[  187]='h0000269e;
    rd_cycle[  188] = 1'b0;  wr_cycle[  188] = 1'b1;  addr_rom[  188]='h000002f0;  wr_data_rom[  188]='h00003fe3;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000002f4;  wr_data_rom[  189]='h000013aa;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000002f8;  wr_data_rom[  190]='h00002e0c;
    rd_cycle[  191] = 1'b0;  wr_cycle[  191] = 1'b1;  addr_rom[  191]='h000002fc;  wr_data_rom[  191]='h00002bbe;
    rd_cycle[  192] = 1'b0;  wr_cycle[  192] = 1'b1;  addr_rom[  192]='h00000300;  wr_data_rom[  192]='h000024ec;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000304;  wr_data_rom[  193]='h00002188;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000308;  wr_data_rom[  194]='h00000051;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h0000030c;  wr_data_rom[  195]='h0000112f;
    rd_cycle[  196] = 1'b0;  wr_cycle[  196] = 1'b1;  addr_rom[  196]='h00000310;  wr_data_rom[  196]='h0000325d;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h00000314;  wr_data_rom[  197]='h00002c55;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h00000318;  wr_data_rom[  198]='h00000ee9;
    rd_cycle[  199] = 1'b0;  wr_cycle[  199] = 1'b1;  addr_rom[  199]='h0000031c;  wr_data_rom[  199]='h00000c7e;
    rd_cycle[  200] = 1'b0;  wr_cycle[  200] = 1'b1;  addr_rom[  200]='h00000320;  wr_data_rom[  200]='h00003419;
    rd_cycle[  201] = 1'b0;  wr_cycle[  201] = 1'b1;  addr_rom[  201]='h00000324;  wr_data_rom[  201]='h00003341;
    rd_cycle[  202] = 1'b0;  wr_cycle[  202] = 1'b1;  addr_rom[  202]='h00000328;  wr_data_rom[  202]='h00000956;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h0000032c;  wr_data_rom[  203]='h0000011b;
    rd_cycle[  204] = 1'b0;  wr_cycle[  204] = 1'b1;  addr_rom[  204]='h00000330;  wr_data_rom[  204]='h0000392c;
    rd_cycle[  205] = 1'b0;  wr_cycle[  205] = 1'b1;  addr_rom[  205]='h00000334;  wr_data_rom[  205]='h00000a4c;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000338;  wr_data_rom[  206]='h000029c7;
    rd_cycle[  207] = 1'b0;  wr_cycle[  207] = 1'b1;  addr_rom[  207]='h0000033c;  wr_data_rom[  207]='h000012ea;
    rd_cycle[  208] = 1'b0;  wr_cycle[  208] = 1'b1;  addr_rom[  208]='h00000340;  wr_data_rom[  208]='h00001b55;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000344;  wr_data_rom[  209]='h00000126;
    rd_cycle[  210] = 1'b0;  wr_cycle[  210] = 1'b1;  addr_rom[  210]='h00000348;  wr_data_rom[  210]='h0000371d;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h0000034c;  wr_data_rom[  211]='h00003b53;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000350;  wr_data_rom[  212]='h00001e4e;
    rd_cycle[  213] = 1'b0;  wr_cycle[  213] = 1'b1;  addr_rom[  213]='h00000354;  wr_data_rom[  213]='h00003615;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000358;  wr_data_rom[  214]='h00002fab;
    rd_cycle[  215] = 1'b0;  wr_cycle[  215] = 1'b1;  addr_rom[  215]='h0000035c;  wr_data_rom[  215]='h0000068d;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h00000360;  wr_data_rom[  216]='h00000000;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h00000364;  wr_data_rom[  217]='h00000624;
    rd_cycle[  218] = 1'b0;  wr_cycle[  218] = 1'b1;  addr_rom[  218]='h00000368;  wr_data_rom[  218]='h000028e9;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h0000036c;  wr_data_rom[  219]='h0000381e;
    rd_cycle[  220] = 1'b0;  wr_cycle[  220] = 1'b1;  addr_rom[  220]='h00000370;  wr_data_rom[  220]='h0000255c;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h00000374;  wr_data_rom[  221]='h00001b9f;
    rd_cycle[  222] = 1'b0;  wr_cycle[  222] = 1'b1;  addr_rom[  222]='h00000378;  wr_data_rom[  222]='h0000002f;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h0000037c;  wr_data_rom[  223]='h000031e1;
    rd_cycle[  224] = 1'b0;  wr_cycle[  224] = 1'b1;  addr_rom[  224]='h00000380;  wr_data_rom[  224]='h000025d1;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000384;  wr_data_rom[  225]='h00000188;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000388;  wr_data_rom[  226]='h00003e9c;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h0000038c;  wr_data_rom[  227]='h00001d15;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000390;  wr_data_rom[  228]='h000029d0;
    rd_cycle[  229] = 1'b0;  wr_cycle[  229] = 1'b1;  addr_rom[  229]='h00000394;  wr_data_rom[  229]='h000011a0;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h00000398;  wr_data_rom[  230]='h000015e6;
    rd_cycle[  231] = 1'b0;  wr_cycle[  231] = 1'b1;  addr_rom[  231]='h0000039c;  wr_data_rom[  231]='h000025c9;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h000003a0;  wr_data_rom[  232]='h00002607;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h000003a4;  wr_data_rom[  233]='h00003e1d;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h000003a8;  wr_data_rom[  234]='h00000e06;
    rd_cycle[  235] = 1'b0;  wr_cycle[  235] = 1'b1;  addr_rom[  235]='h000003ac;  wr_data_rom[  235]='h00003a2a;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000003b0;  wr_data_rom[  236]='h00002447;
    rd_cycle[  237] = 1'b0;  wr_cycle[  237] = 1'b1;  addr_rom[  237]='h000003b4;  wr_data_rom[  237]='h00003349;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h000003b8;  wr_data_rom[  238]='h000015e6;
    rd_cycle[  239] = 1'b0;  wr_cycle[  239] = 1'b1;  addr_rom[  239]='h000003bc;  wr_data_rom[  239]='h00003cb8;
    rd_cycle[  240] = 1'b0;  wr_cycle[  240] = 1'b1;  addr_rom[  240]='h000003c0;  wr_data_rom[  240]='h00001406;
    rd_cycle[  241] = 1'b0;  wr_cycle[  241] = 1'b1;  addr_rom[  241]='h000003c4;  wr_data_rom[  241]='h0000230b;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h000003c8;  wr_data_rom[  242]='h00002b3a;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h000003cc;  wr_data_rom[  243]='h000030f3;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h000003d0;  wr_data_rom[  244]='h0000322e;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h000003d4;  wr_data_rom[  245]='h00000ac8;
    rd_cycle[  246] = 1'b0;  wr_cycle[  246] = 1'b1;  addr_rom[  246]='h000003d8;  wr_data_rom[  246]='h000029ad;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h000003dc;  wr_data_rom[  247]='h00003691;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000003e0;  wr_data_rom[  248]='h00001c05;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h000003e4;  wr_data_rom[  249]='h000010a4;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h000003e8;  wr_data_rom[  250]='h00003d6e;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h000003ec;  wr_data_rom[  251]='h000012e3;
    rd_cycle[  252] = 1'b0;  wr_cycle[  252] = 1'b1;  addr_rom[  252]='h000003f0;  wr_data_rom[  252]='h00001612;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h000003f4;  wr_data_rom[  253]='h00001ac5;
    rd_cycle[  254] = 1'b0;  wr_cycle[  254] = 1'b1;  addr_rom[  254]='h000003f8;  wr_data_rom[  254]='h000038a0;
    rd_cycle[  255] = 1'b0;  wr_cycle[  255] = 1'b1;  addr_rom[  255]='h000003fc;  wr_data_rom[  255]='h000036d9;
    rd_cycle[  256] = 1'b0;  wr_cycle[  256] = 1'b1;  addr_rom[  256]='h00000400;  wr_data_rom[  256]='h000035d6;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h00000404;  wr_data_rom[  257]='h0000139a;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000408;  wr_data_rom[  258]='h000000fa;
    rd_cycle[  259] = 1'b0;  wr_cycle[  259] = 1'b1;  addr_rom[  259]='h0000040c;  wr_data_rom[  259]='h00002436;
    rd_cycle[  260] = 1'b0;  wr_cycle[  260] = 1'b1;  addr_rom[  260]='h00000410;  wr_data_rom[  260]='h00000776;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000414;  wr_data_rom[  261]='h00002e1a;
    rd_cycle[  262] = 1'b0;  wr_cycle[  262] = 1'b1;  addr_rom[  262]='h00000418;  wr_data_rom[  262]='h00000d1e;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h0000041c;  wr_data_rom[  263]='h00003a7a;
    rd_cycle[  264] = 1'b0;  wr_cycle[  264] = 1'b1;  addr_rom[  264]='h00000420;  wr_data_rom[  264]='h00000d85;
    rd_cycle[  265] = 1'b0;  wr_cycle[  265] = 1'b1;  addr_rom[  265]='h00000424;  wr_data_rom[  265]='h000021f5;
    rd_cycle[  266] = 1'b0;  wr_cycle[  266] = 1'b1;  addr_rom[  266]='h00000428;  wr_data_rom[  266]='h00000b10;
    rd_cycle[  267] = 1'b0;  wr_cycle[  267] = 1'b1;  addr_rom[  267]='h0000042c;  wr_data_rom[  267]='h00003341;
    rd_cycle[  268] = 1'b0;  wr_cycle[  268] = 1'b1;  addr_rom[  268]='h00000430;  wr_data_rom[  268]='h00000492;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h00000434;  wr_data_rom[  269]='h00000a4d;
    rd_cycle[  270] = 1'b0;  wr_cycle[  270] = 1'b1;  addr_rom[  270]='h00000438;  wr_data_rom[  270]='h00001097;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h0000043c;  wr_data_rom[  271]='h00003ee3;
    rd_cycle[  272] = 1'b0;  wr_cycle[  272] = 1'b1;  addr_rom[  272]='h00000440;  wr_data_rom[  272]='h000014fa;
    rd_cycle[  273] = 1'b0;  wr_cycle[  273] = 1'b1;  addr_rom[  273]='h00000444;  wr_data_rom[  273]='h00002bc2;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000448;  wr_data_rom[  274]='h00002dda;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h0000044c;  wr_data_rom[  275]='h00000cb4;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h00000450;  wr_data_rom[  276]='h00003a32;
    rd_cycle[  277] = 1'b0;  wr_cycle[  277] = 1'b1;  addr_rom[  277]='h00000454;  wr_data_rom[  277]='h00001929;
    rd_cycle[  278] = 1'b0;  wr_cycle[  278] = 1'b1;  addr_rom[  278]='h00000458;  wr_data_rom[  278]='h000000d3;
    rd_cycle[  279] = 1'b0;  wr_cycle[  279] = 1'b1;  addr_rom[  279]='h0000045c;  wr_data_rom[  279]='h00002ee7;
    rd_cycle[  280] = 1'b0;  wr_cycle[  280] = 1'b1;  addr_rom[  280]='h00000460;  wr_data_rom[  280]='h00003724;
    rd_cycle[  281] = 1'b0;  wr_cycle[  281] = 1'b1;  addr_rom[  281]='h00000464;  wr_data_rom[  281]='h00003466;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h00000468;  wr_data_rom[  282]='h0000240b;
    rd_cycle[  283] = 1'b0;  wr_cycle[  283] = 1'b1;  addr_rom[  283]='h0000046c;  wr_data_rom[  283]='h0000395b;
    rd_cycle[  284] = 1'b0;  wr_cycle[  284] = 1'b1;  addr_rom[  284]='h00000470;  wr_data_rom[  284]='h00002394;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h00000474;  wr_data_rom[  285]='h000015e3;
    rd_cycle[  286] = 1'b0;  wr_cycle[  286] = 1'b1;  addr_rom[  286]='h00000478;  wr_data_rom[  286]='h000017f1;
    rd_cycle[  287] = 1'b0;  wr_cycle[  287] = 1'b1;  addr_rom[  287]='h0000047c;  wr_data_rom[  287]='h000005ee;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h00000480;  wr_data_rom[  288]='h000009d7;
    rd_cycle[  289] = 1'b0;  wr_cycle[  289] = 1'b1;  addr_rom[  289]='h00000484;  wr_data_rom[  289]='h000003b4;
    rd_cycle[  290] = 1'b0;  wr_cycle[  290] = 1'b1;  addr_rom[  290]='h00000488;  wr_data_rom[  290]='h00001ca1;
    rd_cycle[  291] = 1'b0;  wr_cycle[  291] = 1'b1;  addr_rom[  291]='h0000048c;  wr_data_rom[  291]='h0000021e;
    rd_cycle[  292] = 1'b0;  wr_cycle[  292] = 1'b1;  addr_rom[  292]='h00000490;  wr_data_rom[  292]='h00003ecc;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h00000494;  wr_data_rom[  293]='h00001af5;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h00000498;  wr_data_rom[  294]='h00000320;
    rd_cycle[  295] = 1'b0;  wr_cycle[  295] = 1'b1;  addr_rom[  295]='h0000049c;  wr_data_rom[  295]='h00003e13;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h000004a0;  wr_data_rom[  296]='h00002d96;
    rd_cycle[  297] = 1'b0;  wr_cycle[  297] = 1'b1;  addr_rom[  297]='h000004a4;  wr_data_rom[  297]='h00002a6c;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h000004a8;  wr_data_rom[  298]='h00002999;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h000004ac;  wr_data_rom[  299]='h00003c08;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h000004b0;  wr_data_rom[  300]='h00000574;
    rd_cycle[  301] = 1'b0;  wr_cycle[  301] = 1'b1;  addr_rom[  301]='h000004b4;  wr_data_rom[  301]='h00003ff8;
    rd_cycle[  302] = 1'b0;  wr_cycle[  302] = 1'b1;  addr_rom[  302]='h000004b8;  wr_data_rom[  302]='h000036d3;
    rd_cycle[  303] = 1'b0;  wr_cycle[  303] = 1'b1;  addr_rom[  303]='h000004bc;  wr_data_rom[  303]='h00003fe7;
    rd_cycle[  304] = 1'b0;  wr_cycle[  304] = 1'b1;  addr_rom[  304]='h000004c0;  wr_data_rom[  304]='h000034f8;
    rd_cycle[  305] = 1'b0;  wr_cycle[  305] = 1'b1;  addr_rom[  305]='h000004c4;  wr_data_rom[  305]='h00001d9b;
    rd_cycle[  306] = 1'b0;  wr_cycle[  306] = 1'b1;  addr_rom[  306]='h000004c8;  wr_data_rom[  306]='h00000e9d;
    rd_cycle[  307] = 1'b0;  wr_cycle[  307] = 1'b1;  addr_rom[  307]='h000004cc;  wr_data_rom[  307]='h00003aa7;
    rd_cycle[  308] = 1'b0;  wr_cycle[  308] = 1'b1;  addr_rom[  308]='h000004d0;  wr_data_rom[  308]='h0000193b;
    rd_cycle[  309] = 1'b0;  wr_cycle[  309] = 1'b1;  addr_rom[  309]='h000004d4;  wr_data_rom[  309]='h000010dc;
    rd_cycle[  310] = 1'b0;  wr_cycle[  310] = 1'b1;  addr_rom[  310]='h000004d8;  wr_data_rom[  310]='h00003174;
    rd_cycle[  311] = 1'b0;  wr_cycle[  311] = 1'b1;  addr_rom[  311]='h000004dc;  wr_data_rom[  311]='h00003351;
    rd_cycle[  312] = 1'b0;  wr_cycle[  312] = 1'b1;  addr_rom[  312]='h000004e0;  wr_data_rom[  312]='h00000db4;
    rd_cycle[  313] = 1'b0;  wr_cycle[  313] = 1'b1;  addr_rom[  313]='h000004e4;  wr_data_rom[  313]='h00002dde;
    rd_cycle[  314] = 1'b0;  wr_cycle[  314] = 1'b1;  addr_rom[  314]='h000004e8;  wr_data_rom[  314]='h00000dd4;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h000004ec;  wr_data_rom[  315]='h00002bcd;
    rd_cycle[  316] = 1'b0;  wr_cycle[  316] = 1'b1;  addr_rom[  316]='h000004f0;  wr_data_rom[  316]='h00000e27;
    rd_cycle[  317] = 1'b0;  wr_cycle[  317] = 1'b1;  addr_rom[  317]='h000004f4;  wr_data_rom[  317]='h00002f3b;
    rd_cycle[  318] = 1'b0;  wr_cycle[  318] = 1'b1;  addr_rom[  318]='h000004f8;  wr_data_rom[  318]='h000003c1;
    rd_cycle[  319] = 1'b0;  wr_cycle[  319] = 1'b1;  addr_rom[  319]='h000004fc;  wr_data_rom[  319]='h0000063e;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000500;  wr_data_rom[  320]='h0000347b;
    rd_cycle[  321] = 1'b0;  wr_cycle[  321] = 1'b1;  addr_rom[  321]='h00000504;  wr_data_rom[  321]='h00003e26;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h00000508;  wr_data_rom[  322]='h0000202f;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h0000050c;  wr_data_rom[  323]='h0000138a;
    rd_cycle[  324] = 1'b0;  wr_cycle[  324] = 1'b1;  addr_rom[  324]='h00000510;  wr_data_rom[  324]='h000006c4;
    rd_cycle[  325] = 1'b0;  wr_cycle[  325] = 1'b1;  addr_rom[  325]='h00000514;  wr_data_rom[  325]='h00003445;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000518;  wr_data_rom[  326]='h00001522;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h0000051c;  wr_data_rom[  327]='h00001a56;
    rd_cycle[  328] = 1'b0;  wr_cycle[  328] = 1'b1;  addr_rom[  328]='h00000520;  wr_data_rom[  328]='h00000d43;
    rd_cycle[  329] = 1'b0;  wr_cycle[  329] = 1'b1;  addr_rom[  329]='h00000524;  wr_data_rom[  329]='h00002109;
    rd_cycle[  330] = 1'b0;  wr_cycle[  330] = 1'b1;  addr_rom[  330]='h00000528;  wr_data_rom[  330]='h0000371c;
    rd_cycle[  331] = 1'b0;  wr_cycle[  331] = 1'b1;  addr_rom[  331]='h0000052c;  wr_data_rom[  331]='h00003166;
    rd_cycle[  332] = 1'b0;  wr_cycle[  332] = 1'b1;  addr_rom[  332]='h00000530;  wr_data_rom[  332]='h000030df;
    rd_cycle[  333] = 1'b0;  wr_cycle[  333] = 1'b1;  addr_rom[  333]='h00000534;  wr_data_rom[  333]='h000023da;
    rd_cycle[  334] = 1'b0;  wr_cycle[  334] = 1'b1;  addr_rom[  334]='h00000538;  wr_data_rom[  334]='h000034f7;
    rd_cycle[  335] = 1'b0;  wr_cycle[  335] = 1'b1;  addr_rom[  335]='h0000053c;  wr_data_rom[  335]='h00003ecd;
    rd_cycle[  336] = 1'b0;  wr_cycle[  336] = 1'b1;  addr_rom[  336]='h00000540;  wr_data_rom[  336]='h00000ac8;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h00000544;  wr_data_rom[  337]='h00000050;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000548;  wr_data_rom[  338]='h00001b5e;
    rd_cycle[  339] = 1'b0;  wr_cycle[  339] = 1'b1;  addr_rom[  339]='h0000054c;  wr_data_rom[  339]='h0000009e;
    rd_cycle[  340] = 1'b0;  wr_cycle[  340] = 1'b1;  addr_rom[  340]='h00000550;  wr_data_rom[  340]='h000036cb;
    rd_cycle[  341] = 1'b0;  wr_cycle[  341] = 1'b1;  addr_rom[  341]='h00000554;  wr_data_rom[  341]='h000015ea;
    rd_cycle[  342] = 1'b0;  wr_cycle[  342] = 1'b1;  addr_rom[  342]='h00000558;  wr_data_rom[  342]='h00000030;
    rd_cycle[  343] = 1'b0;  wr_cycle[  343] = 1'b1;  addr_rom[  343]='h0000055c;  wr_data_rom[  343]='h00001933;
    rd_cycle[  344] = 1'b0;  wr_cycle[  344] = 1'b1;  addr_rom[  344]='h00000560;  wr_data_rom[  344]='h00002412;
    rd_cycle[  345] = 1'b0;  wr_cycle[  345] = 1'b1;  addr_rom[  345]='h00000564;  wr_data_rom[  345]='h00000eff;
    rd_cycle[  346] = 1'b0;  wr_cycle[  346] = 1'b1;  addr_rom[  346]='h00000568;  wr_data_rom[  346]='h0000059f;
    rd_cycle[  347] = 1'b0;  wr_cycle[  347] = 1'b1;  addr_rom[  347]='h0000056c;  wr_data_rom[  347]='h0000015a;
    rd_cycle[  348] = 1'b0;  wr_cycle[  348] = 1'b1;  addr_rom[  348]='h00000570;  wr_data_rom[  348]='h00001e80;
    rd_cycle[  349] = 1'b0;  wr_cycle[  349] = 1'b1;  addr_rom[  349]='h00000574;  wr_data_rom[  349]='h00000182;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h00000578;  wr_data_rom[  350]='h00001fa3;
    rd_cycle[  351] = 1'b0;  wr_cycle[  351] = 1'b1;  addr_rom[  351]='h0000057c;  wr_data_rom[  351]='h0000166a;
    rd_cycle[  352] = 1'b0;  wr_cycle[  352] = 1'b1;  addr_rom[  352]='h00000580;  wr_data_rom[  352]='h00001c60;
    rd_cycle[  353] = 1'b0;  wr_cycle[  353] = 1'b1;  addr_rom[  353]='h00000584;  wr_data_rom[  353]='h00003533;
    rd_cycle[  354] = 1'b0;  wr_cycle[  354] = 1'b1;  addr_rom[  354]='h00000588;  wr_data_rom[  354]='h000007e8;
    rd_cycle[  355] = 1'b0;  wr_cycle[  355] = 1'b1;  addr_rom[  355]='h0000058c;  wr_data_rom[  355]='h00002e16;
    rd_cycle[  356] = 1'b0;  wr_cycle[  356] = 1'b1;  addr_rom[  356]='h00000590;  wr_data_rom[  356]='h00000e18;
    rd_cycle[  357] = 1'b0;  wr_cycle[  357] = 1'b1;  addr_rom[  357]='h00000594;  wr_data_rom[  357]='h00002735;
    rd_cycle[  358] = 1'b0;  wr_cycle[  358] = 1'b1;  addr_rom[  358]='h00000598;  wr_data_rom[  358]='h00001b81;
    rd_cycle[  359] = 1'b0;  wr_cycle[  359] = 1'b1;  addr_rom[  359]='h0000059c;  wr_data_rom[  359]='h00000dda;
    rd_cycle[  360] = 1'b0;  wr_cycle[  360] = 1'b1;  addr_rom[  360]='h000005a0;  wr_data_rom[  360]='h00002676;
    rd_cycle[  361] = 1'b0;  wr_cycle[  361] = 1'b1;  addr_rom[  361]='h000005a4;  wr_data_rom[  361]='h00001ec2;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h000005a8;  wr_data_rom[  362]='h00003b37;
    rd_cycle[  363] = 1'b0;  wr_cycle[  363] = 1'b1;  addr_rom[  363]='h000005ac;  wr_data_rom[  363]='h000032c5;
    rd_cycle[  364] = 1'b0;  wr_cycle[  364] = 1'b1;  addr_rom[  364]='h000005b0;  wr_data_rom[  364]='h00002c0b;
    rd_cycle[  365] = 1'b0;  wr_cycle[  365] = 1'b1;  addr_rom[  365]='h000005b4;  wr_data_rom[  365]='h00000065;
    rd_cycle[  366] = 1'b0;  wr_cycle[  366] = 1'b1;  addr_rom[  366]='h000005b8;  wr_data_rom[  366]='h00001689;
    rd_cycle[  367] = 1'b0;  wr_cycle[  367] = 1'b1;  addr_rom[  367]='h000005bc;  wr_data_rom[  367]='h00000667;
    rd_cycle[  368] = 1'b0;  wr_cycle[  368] = 1'b1;  addr_rom[  368]='h000005c0;  wr_data_rom[  368]='h00002e41;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h000005c4;  wr_data_rom[  369]='h00003e97;
    rd_cycle[  370] = 1'b0;  wr_cycle[  370] = 1'b1;  addr_rom[  370]='h000005c8;  wr_data_rom[  370]='h00000e21;
    rd_cycle[  371] = 1'b0;  wr_cycle[  371] = 1'b1;  addr_rom[  371]='h000005cc;  wr_data_rom[  371]='h0000311c;
    rd_cycle[  372] = 1'b0;  wr_cycle[  372] = 1'b1;  addr_rom[  372]='h000005d0;  wr_data_rom[  372]='h000013ac;
    rd_cycle[  373] = 1'b0;  wr_cycle[  373] = 1'b1;  addr_rom[  373]='h000005d4;  wr_data_rom[  373]='h000001d2;
    rd_cycle[  374] = 1'b0;  wr_cycle[  374] = 1'b1;  addr_rom[  374]='h000005d8;  wr_data_rom[  374]='h00000efd;
    rd_cycle[  375] = 1'b0;  wr_cycle[  375] = 1'b1;  addr_rom[  375]='h000005dc;  wr_data_rom[  375]='h0000287a;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h000005e0;  wr_data_rom[  376]='h00003ff8;
    rd_cycle[  377] = 1'b0;  wr_cycle[  377] = 1'b1;  addr_rom[  377]='h000005e4;  wr_data_rom[  377]='h00003887;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h000005e8;  wr_data_rom[  378]='h0000255b;
    rd_cycle[  379] = 1'b0;  wr_cycle[  379] = 1'b1;  addr_rom[  379]='h000005ec;  wr_data_rom[  379]='h0000068a;
    rd_cycle[  380] = 1'b0;  wr_cycle[  380] = 1'b1;  addr_rom[  380]='h000005f0;  wr_data_rom[  380]='h00003ee2;
    rd_cycle[  381] = 1'b0;  wr_cycle[  381] = 1'b1;  addr_rom[  381]='h000005f4;  wr_data_rom[  381]='h00000530;
    rd_cycle[  382] = 1'b0;  wr_cycle[  382] = 1'b1;  addr_rom[  382]='h000005f8;  wr_data_rom[  382]='h000003ad;
    rd_cycle[  383] = 1'b0;  wr_cycle[  383] = 1'b1;  addr_rom[  383]='h000005fc;  wr_data_rom[  383]='h00002041;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h00000600;  wr_data_rom[  384]='h00001c64;
    rd_cycle[  385] = 1'b0;  wr_cycle[  385] = 1'b1;  addr_rom[  385]='h00000604;  wr_data_rom[  385]='h00000ef2;
    rd_cycle[  386] = 1'b0;  wr_cycle[  386] = 1'b1;  addr_rom[  386]='h00000608;  wr_data_rom[  386]='h00003b94;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h0000060c;  wr_data_rom[  387]='h00001b16;
    rd_cycle[  388] = 1'b0;  wr_cycle[  388] = 1'b1;  addr_rom[  388]='h00000610;  wr_data_rom[  388]='h000005c7;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h00000614;  wr_data_rom[  389]='h00002194;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h00000618;  wr_data_rom[  390]='h0000228d;
    rd_cycle[  391] = 1'b0;  wr_cycle[  391] = 1'b1;  addr_rom[  391]='h0000061c;  wr_data_rom[  391]='h00000716;
    rd_cycle[  392] = 1'b0;  wr_cycle[  392] = 1'b1;  addr_rom[  392]='h00000620;  wr_data_rom[  392]='h00002413;
    rd_cycle[  393] = 1'b0;  wr_cycle[  393] = 1'b1;  addr_rom[  393]='h00000624;  wr_data_rom[  393]='h00002588;
    rd_cycle[  394] = 1'b0;  wr_cycle[  394] = 1'b1;  addr_rom[  394]='h00000628;  wr_data_rom[  394]='h0000180e;
    rd_cycle[  395] = 1'b0;  wr_cycle[  395] = 1'b1;  addr_rom[  395]='h0000062c;  wr_data_rom[  395]='h00000470;
    rd_cycle[  396] = 1'b0;  wr_cycle[  396] = 1'b1;  addr_rom[  396]='h00000630;  wr_data_rom[  396]='h00000e38;
    rd_cycle[  397] = 1'b0;  wr_cycle[  397] = 1'b1;  addr_rom[  397]='h00000634;  wr_data_rom[  397]='h00001831;
    rd_cycle[  398] = 1'b0;  wr_cycle[  398] = 1'b1;  addr_rom[  398]='h00000638;  wr_data_rom[  398]='h00000c07;
    rd_cycle[  399] = 1'b0;  wr_cycle[  399] = 1'b1;  addr_rom[  399]='h0000063c;  wr_data_rom[  399]='h0000198e;
    rd_cycle[  400] = 1'b0;  wr_cycle[  400] = 1'b1;  addr_rom[  400]='h00000640;  wr_data_rom[  400]='h000020ea;
    rd_cycle[  401] = 1'b0;  wr_cycle[  401] = 1'b1;  addr_rom[  401]='h00000644;  wr_data_rom[  401]='h00003798;
    rd_cycle[  402] = 1'b0;  wr_cycle[  402] = 1'b1;  addr_rom[  402]='h00000648;  wr_data_rom[  402]='h00003aa2;
    rd_cycle[  403] = 1'b0;  wr_cycle[  403] = 1'b1;  addr_rom[  403]='h0000064c;  wr_data_rom[  403]='h0000357f;
    rd_cycle[  404] = 1'b0;  wr_cycle[  404] = 1'b1;  addr_rom[  404]='h00000650;  wr_data_rom[  404]='h00003b3d;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b1;  addr_rom[  405]='h00000654;  wr_data_rom[  405]='h00002fc4;
    rd_cycle[  406] = 1'b0;  wr_cycle[  406] = 1'b1;  addr_rom[  406]='h00000658;  wr_data_rom[  406]='h00001f7c;
    rd_cycle[  407] = 1'b0;  wr_cycle[  407] = 1'b1;  addr_rom[  407]='h0000065c;  wr_data_rom[  407]='h00001f7e;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b1;  addr_rom[  408]='h00000660;  wr_data_rom[  408]='h00000d6c;
    rd_cycle[  409] = 1'b0;  wr_cycle[  409] = 1'b1;  addr_rom[  409]='h00000664;  wr_data_rom[  409]='h000032df;
    rd_cycle[  410] = 1'b0;  wr_cycle[  410] = 1'b1;  addr_rom[  410]='h00000668;  wr_data_rom[  410]='h000010f5;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b1;  addr_rom[  411]='h0000066c;  wr_data_rom[  411]='h000009af;
    rd_cycle[  412] = 1'b0;  wr_cycle[  412] = 1'b1;  addr_rom[  412]='h00000670;  wr_data_rom[  412]='h00000a3b;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b1;  addr_rom[  413]='h00000674;  wr_data_rom[  413]='h00003a3a;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b1;  addr_rom[  414]='h00000678;  wr_data_rom[  414]='h000016b5;
    rd_cycle[  415] = 1'b0;  wr_cycle[  415] = 1'b1;  addr_rom[  415]='h0000067c;  wr_data_rom[  415]='h0000179b;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b1;  addr_rom[  416]='h00000680;  wr_data_rom[  416]='h00000480;
    rd_cycle[  417] = 1'b0;  wr_cycle[  417] = 1'b1;  addr_rom[  417]='h00000684;  wr_data_rom[  417]='h00002b21;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b1;  addr_rom[  418]='h00000688;  wr_data_rom[  418]='h000037b2;
    rd_cycle[  419] = 1'b0;  wr_cycle[  419] = 1'b1;  addr_rom[  419]='h0000068c;  wr_data_rom[  419]='h00003156;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b1;  addr_rom[  420]='h00000690;  wr_data_rom[  420]='h000036f3;
    rd_cycle[  421] = 1'b0;  wr_cycle[  421] = 1'b1;  addr_rom[  421]='h00000694;  wr_data_rom[  421]='h0000242b;
    rd_cycle[  422] = 1'b0;  wr_cycle[  422] = 1'b1;  addr_rom[  422]='h00000698;  wr_data_rom[  422]='h00003160;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b1;  addr_rom[  423]='h0000069c;  wr_data_rom[  423]='h00002bc3;
    rd_cycle[  424] = 1'b0;  wr_cycle[  424] = 1'b1;  addr_rom[  424]='h000006a0;  wr_data_rom[  424]='h00000521;
    rd_cycle[  425] = 1'b0;  wr_cycle[  425] = 1'b1;  addr_rom[  425]='h000006a4;  wr_data_rom[  425]='h00000ee6;
    rd_cycle[  426] = 1'b0;  wr_cycle[  426] = 1'b1;  addr_rom[  426]='h000006a8;  wr_data_rom[  426]='h00001c52;
    rd_cycle[  427] = 1'b0;  wr_cycle[  427] = 1'b1;  addr_rom[  427]='h000006ac;  wr_data_rom[  427]='h0000160a;
    rd_cycle[  428] = 1'b0;  wr_cycle[  428] = 1'b1;  addr_rom[  428]='h000006b0;  wr_data_rom[  428]='h00001f40;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b1;  addr_rom[  429]='h000006b4;  wr_data_rom[  429]='h00000da7;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b1;  addr_rom[  430]='h000006b8;  wr_data_rom[  430]='h0000137c;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b1;  addr_rom[  431]='h000006bc;  wr_data_rom[  431]='h00003767;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b1;  addr_rom[  432]='h000006c0;  wr_data_rom[  432]='h0000280b;
    rd_cycle[  433] = 1'b0;  wr_cycle[  433] = 1'b1;  addr_rom[  433]='h000006c4;  wr_data_rom[  433]='h00001e4e;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b1;  addr_rom[  434]='h000006c8;  wr_data_rom[  434]='h00003510;
    rd_cycle[  435] = 1'b0;  wr_cycle[  435] = 1'b1;  addr_rom[  435]='h000006cc;  wr_data_rom[  435]='h000033c8;
    rd_cycle[  436] = 1'b0;  wr_cycle[  436] = 1'b1;  addr_rom[  436]='h000006d0;  wr_data_rom[  436]='h00000f70;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b1;  addr_rom[  437]='h000006d4;  wr_data_rom[  437]='h000036b8;
    rd_cycle[  438] = 1'b0;  wr_cycle[  438] = 1'b1;  addr_rom[  438]='h000006d8;  wr_data_rom[  438]='h00003a5a;
    rd_cycle[  439] = 1'b0;  wr_cycle[  439] = 1'b1;  addr_rom[  439]='h000006dc;  wr_data_rom[  439]='h00001a1e;
    rd_cycle[  440] = 1'b0;  wr_cycle[  440] = 1'b1;  addr_rom[  440]='h000006e0;  wr_data_rom[  440]='h00002cfa;
    rd_cycle[  441] = 1'b0;  wr_cycle[  441] = 1'b1;  addr_rom[  441]='h000006e4;  wr_data_rom[  441]='h00003be4;
    rd_cycle[  442] = 1'b0;  wr_cycle[  442] = 1'b1;  addr_rom[  442]='h000006e8;  wr_data_rom[  442]='h000018d6;
    rd_cycle[  443] = 1'b0;  wr_cycle[  443] = 1'b1;  addr_rom[  443]='h000006ec;  wr_data_rom[  443]='h00003fb5;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b1;  addr_rom[  444]='h000006f0;  wr_data_rom[  444]='h00001fcc;
    rd_cycle[  445] = 1'b0;  wr_cycle[  445] = 1'b1;  addr_rom[  445]='h000006f4;  wr_data_rom[  445]='h00003dc1;
    rd_cycle[  446] = 1'b0;  wr_cycle[  446] = 1'b1;  addr_rom[  446]='h000006f8;  wr_data_rom[  446]='h00003291;
    rd_cycle[  447] = 1'b0;  wr_cycle[  447] = 1'b1;  addr_rom[  447]='h000006fc;  wr_data_rom[  447]='h00002671;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b1;  addr_rom[  448]='h00000700;  wr_data_rom[  448]='h00003278;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b1;  addr_rom[  449]='h00000704;  wr_data_rom[  449]='h00002a09;
    rd_cycle[  450] = 1'b0;  wr_cycle[  450] = 1'b1;  addr_rom[  450]='h00000708;  wr_data_rom[  450]='h000000c1;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b1;  addr_rom[  451]='h0000070c;  wr_data_rom[  451]='h00001cd6;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b1;  addr_rom[  452]='h00000710;  wr_data_rom[  452]='h000028e0;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b1;  addr_rom[  453]='h00000714;  wr_data_rom[  453]='h00000521;
    rd_cycle[  454] = 1'b0;  wr_cycle[  454] = 1'b1;  addr_rom[  454]='h00000718;  wr_data_rom[  454]='h000007ca;
    rd_cycle[  455] = 1'b0;  wr_cycle[  455] = 1'b1;  addr_rom[  455]='h0000071c;  wr_data_rom[  455]='h00000b0f;
    rd_cycle[  456] = 1'b0;  wr_cycle[  456] = 1'b1;  addr_rom[  456]='h00000720;  wr_data_rom[  456]='h00001bc4;
    rd_cycle[  457] = 1'b0;  wr_cycle[  457] = 1'b1;  addr_rom[  457]='h00000724;  wr_data_rom[  457]='h00000eb3;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b1;  addr_rom[  458]='h00000728;  wr_data_rom[  458]='h000037cd;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b1;  addr_rom[  459]='h0000072c;  wr_data_rom[  459]='h00002288;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b1;  addr_rom[  460]='h00000730;  wr_data_rom[  460]='h000028c2;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b1;  addr_rom[  461]='h00000734;  wr_data_rom[  461]='h00003c99;
    rd_cycle[  462] = 1'b0;  wr_cycle[  462] = 1'b1;  addr_rom[  462]='h00000738;  wr_data_rom[  462]='h00000c8c;
    rd_cycle[  463] = 1'b0;  wr_cycle[  463] = 1'b1;  addr_rom[  463]='h0000073c;  wr_data_rom[  463]='h00000b36;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b1;  addr_rom[  464]='h00000740;  wr_data_rom[  464]='h0000003c;
    rd_cycle[  465] = 1'b0;  wr_cycle[  465] = 1'b1;  addr_rom[  465]='h00000744;  wr_data_rom[  465]='h000017b5;
    rd_cycle[  466] = 1'b0;  wr_cycle[  466] = 1'b1;  addr_rom[  466]='h00000748;  wr_data_rom[  466]='h00002699;
    rd_cycle[  467] = 1'b0;  wr_cycle[  467] = 1'b1;  addr_rom[  467]='h0000074c;  wr_data_rom[  467]='h00003734;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b1;  addr_rom[  468]='h00000750;  wr_data_rom[  468]='h00000c34;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b1;  addr_rom[  469]='h00000754;  wr_data_rom[  469]='h000002e9;
    rd_cycle[  470] = 1'b0;  wr_cycle[  470] = 1'b1;  addr_rom[  470]='h00000758;  wr_data_rom[  470]='h00003901;
    rd_cycle[  471] = 1'b0;  wr_cycle[  471] = 1'b1;  addr_rom[  471]='h0000075c;  wr_data_rom[  471]='h000036df;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b1;  addr_rom[  472]='h00000760;  wr_data_rom[  472]='h00002c9f;
    rd_cycle[  473] = 1'b0;  wr_cycle[  473] = 1'b1;  addr_rom[  473]='h00000764;  wr_data_rom[  473]='h0000089a;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b1;  addr_rom[  474]='h00000768;  wr_data_rom[  474]='h000017ba;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b1;  addr_rom[  475]='h0000076c;  wr_data_rom[  475]='h00003889;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b1;  addr_rom[  476]='h00000770;  wr_data_rom[  476]='h00000465;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b1;  addr_rom[  477]='h00000774;  wr_data_rom[  477]='h00002ffa;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b1;  addr_rom[  478]='h00000778;  wr_data_rom[  478]='h00001e66;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b1;  addr_rom[  479]='h0000077c;  wr_data_rom[  479]='h00003622;
    rd_cycle[  480] = 1'b0;  wr_cycle[  480] = 1'b1;  addr_rom[  480]='h00000780;  wr_data_rom[  480]='h00003323;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b1;  addr_rom[  481]='h00000784;  wr_data_rom[  481]='h000003a7;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b1;  addr_rom[  482]='h00000788;  wr_data_rom[  482]='h00001af4;
    rd_cycle[  483] = 1'b0;  wr_cycle[  483] = 1'b1;  addr_rom[  483]='h0000078c;  wr_data_rom[  483]='h00002512;
    rd_cycle[  484] = 1'b0;  wr_cycle[  484] = 1'b1;  addr_rom[  484]='h00000790;  wr_data_rom[  484]='h0000358d;
    rd_cycle[  485] = 1'b0;  wr_cycle[  485] = 1'b1;  addr_rom[  485]='h00000794;  wr_data_rom[  485]='h000009ea;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b1;  addr_rom[  486]='h00000798;  wr_data_rom[  486]='h00000e0e;
    rd_cycle[  487] = 1'b0;  wr_cycle[  487] = 1'b1;  addr_rom[  487]='h0000079c;  wr_data_rom[  487]='h000038a0;
    rd_cycle[  488] = 1'b0;  wr_cycle[  488] = 1'b1;  addr_rom[  488]='h000007a0;  wr_data_rom[  488]='h00001939;
    rd_cycle[  489] = 1'b0;  wr_cycle[  489] = 1'b1;  addr_rom[  489]='h000007a4;  wr_data_rom[  489]='h00003820;
    rd_cycle[  490] = 1'b0;  wr_cycle[  490] = 1'b1;  addr_rom[  490]='h000007a8;  wr_data_rom[  490]='h000004d6;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b1;  addr_rom[  491]='h000007ac;  wr_data_rom[  491]='h00001a69;
    rd_cycle[  492] = 1'b0;  wr_cycle[  492] = 1'b1;  addr_rom[  492]='h000007b0;  wr_data_rom[  492]='h00000603;
    rd_cycle[  493] = 1'b0;  wr_cycle[  493] = 1'b1;  addr_rom[  493]='h000007b4;  wr_data_rom[  493]='h000016b0;
    rd_cycle[  494] = 1'b0;  wr_cycle[  494] = 1'b1;  addr_rom[  494]='h000007b8;  wr_data_rom[  494]='h000012fe;
    rd_cycle[  495] = 1'b0;  wr_cycle[  495] = 1'b1;  addr_rom[  495]='h000007bc;  wr_data_rom[  495]='h00002b95;
    rd_cycle[  496] = 1'b0;  wr_cycle[  496] = 1'b1;  addr_rom[  496]='h000007c0;  wr_data_rom[  496]='h000005af;
    rd_cycle[  497] = 1'b0;  wr_cycle[  497] = 1'b1;  addr_rom[  497]='h000007c4;  wr_data_rom[  497]='h00002917;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b1;  addr_rom[  498]='h000007c8;  wr_data_rom[  498]='h000029c8;
    rd_cycle[  499] = 1'b0;  wr_cycle[  499] = 1'b1;  addr_rom[  499]='h000007cc;  wr_data_rom[  499]='h00002d67;
    rd_cycle[  500] = 1'b0;  wr_cycle[  500] = 1'b1;  addr_rom[  500]='h000007d0;  wr_data_rom[  500]='h00001f58;
    rd_cycle[  501] = 1'b0;  wr_cycle[  501] = 1'b1;  addr_rom[  501]='h000007d4;  wr_data_rom[  501]='h00001b37;
    rd_cycle[  502] = 1'b0;  wr_cycle[  502] = 1'b1;  addr_rom[  502]='h000007d8;  wr_data_rom[  502]='h0000062b;
    rd_cycle[  503] = 1'b0;  wr_cycle[  503] = 1'b1;  addr_rom[  503]='h000007dc;  wr_data_rom[  503]='h00002185;
    rd_cycle[  504] = 1'b0;  wr_cycle[  504] = 1'b1;  addr_rom[  504]='h000007e0;  wr_data_rom[  504]='h00001f96;
    rd_cycle[  505] = 1'b0;  wr_cycle[  505] = 1'b1;  addr_rom[  505]='h000007e4;  wr_data_rom[  505]='h00002f4b;
    rd_cycle[  506] = 1'b0;  wr_cycle[  506] = 1'b1;  addr_rom[  506]='h000007e8;  wr_data_rom[  506]='h00001e01;
    rd_cycle[  507] = 1'b0;  wr_cycle[  507] = 1'b1;  addr_rom[  507]='h000007ec;  wr_data_rom[  507]='h00000f12;
    rd_cycle[  508] = 1'b0;  wr_cycle[  508] = 1'b1;  addr_rom[  508]='h000007f0;  wr_data_rom[  508]='h000020b8;
    rd_cycle[  509] = 1'b0;  wr_cycle[  509] = 1'b1;  addr_rom[  509]='h000007f4;  wr_data_rom[  509]='h00002faf;
    rd_cycle[  510] = 1'b0;  wr_cycle[  510] = 1'b1;  addr_rom[  510]='h000007f8;  wr_data_rom[  510]='h00003891;
    rd_cycle[  511] = 1'b0;  wr_cycle[  511] = 1'b1;  addr_rom[  511]='h000007fc;  wr_data_rom[  511]='h0000360c;
    rd_cycle[  512] = 1'b0;  wr_cycle[  512] = 1'b1;  addr_rom[  512]='h00000800;  wr_data_rom[  512]='h00002b1e;
    rd_cycle[  513] = 1'b0;  wr_cycle[  513] = 1'b1;  addr_rom[  513]='h00000804;  wr_data_rom[  513]='h00001dca;
    rd_cycle[  514] = 1'b0;  wr_cycle[  514] = 1'b1;  addr_rom[  514]='h00000808;  wr_data_rom[  514]='h00003b58;
    rd_cycle[  515] = 1'b0;  wr_cycle[  515] = 1'b1;  addr_rom[  515]='h0000080c;  wr_data_rom[  515]='h000033cf;
    rd_cycle[  516] = 1'b0;  wr_cycle[  516] = 1'b1;  addr_rom[  516]='h00000810;  wr_data_rom[  516]='h00000fc6;
    rd_cycle[  517] = 1'b0;  wr_cycle[  517] = 1'b1;  addr_rom[  517]='h00000814;  wr_data_rom[  517]='h00002dce;
    rd_cycle[  518] = 1'b0;  wr_cycle[  518] = 1'b1;  addr_rom[  518]='h00000818;  wr_data_rom[  518]='h00002470;
    rd_cycle[  519] = 1'b0;  wr_cycle[  519] = 1'b1;  addr_rom[  519]='h0000081c;  wr_data_rom[  519]='h000001a8;
    rd_cycle[  520] = 1'b0;  wr_cycle[  520] = 1'b1;  addr_rom[  520]='h00000820;  wr_data_rom[  520]='h00001900;
    rd_cycle[  521] = 1'b0;  wr_cycle[  521] = 1'b1;  addr_rom[  521]='h00000824;  wr_data_rom[  521]='h00002d68;
    rd_cycle[  522] = 1'b0;  wr_cycle[  522] = 1'b1;  addr_rom[  522]='h00000828;  wr_data_rom[  522]='h00000c2d;
    rd_cycle[  523] = 1'b0;  wr_cycle[  523] = 1'b1;  addr_rom[  523]='h0000082c;  wr_data_rom[  523]='h000029fe;
    rd_cycle[  524] = 1'b0;  wr_cycle[  524] = 1'b1;  addr_rom[  524]='h00000830;  wr_data_rom[  524]='h000013ac;
    rd_cycle[  525] = 1'b0;  wr_cycle[  525] = 1'b1;  addr_rom[  525]='h00000834;  wr_data_rom[  525]='h00003a04;
    rd_cycle[  526] = 1'b0;  wr_cycle[  526] = 1'b1;  addr_rom[  526]='h00000838;  wr_data_rom[  526]='h00000e83;
    rd_cycle[  527] = 1'b0;  wr_cycle[  527] = 1'b1;  addr_rom[  527]='h0000083c;  wr_data_rom[  527]='h00002001;
    rd_cycle[  528] = 1'b0;  wr_cycle[  528] = 1'b1;  addr_rom[  528]='h00000840;  wr_data_rom[  528]='h00003631;
    rd_cycle[  529] = 1'b0;  wr_cycle[  529] = 1'b1;  addr_rom[  529]='h00000844;  wr_data_rom[  529]='h00001930;
    rd_cycle[  530] = 1'b0;  wr_cycle[  530] = 1'b1;  addr_rom[  530]='h00000848;  wr_data_rom[  530]='h00001701;
    rd_cycle[  531] = 1'b0;  wr_cycle[  531] = 1'b1;  addr_rom[  531]='h0000084c;  wr_data_rom[  531]='h00001e31;
    rd_cycle[  532] = 1'b0;  wr_cycle[  532] = 1'b1;  addr_rom[  532]='h00000850;  wr_data_rom[  532]='h000020f3;
    rd_cycle[  533] = 1'b0;  wr_cycle[  533] = 1'b1;  addr_rom[  533]='h00000854;  wr_data_rom[  533]='h0000320b;
    rd_cycle[  534] = 1'b0;  wr_cycle[  534] = 1'b1;  addr_rom[  534]='h00000858;  wr_data_rom[  534]='h00001623;
    rd_cycle[  535] = 1'b0;  wr_cycle[  535] = 1'b1;  addr_rom[  535]='h0000085c;  wr_data_rom[  535]='h00000f48;
    rd_cycle[  536] = 1'b0;  wr_cycle[  536] = 1'b1;  addr_rom[  536]='h00000860;  wr_data_rom[  536]='h00000291;
    rd_cycle[  537] = 1'b0;  wr_cycle[  537] = 1'b1;  addr_rom[  537]='h00000864;  wr_data_rom[  537]='h00001a9e;
    rd_cycle[  538] = 1'b0;  wr_cycle[  538] = 1'b1;  addr_rom[  538]='h00000868;  wr_data_rom[  538]='h0000165b;
    rd_cycle[  539] = 1'b0;  wr_cycle[  539] = 1'b1;  addr_rom[  539]='h0000086c;  wr_data_rom[  539]='h00002baf;
    rd_cycle[  540] = 1'b0;  wr_cycle[  540] = 1'b1;  addr_rom[  540]='h00000870;  wr_data_rom[  540]='h00000e87;
    rd_cycle[  541] = 1'b0;  wr_cycle[  541] = 1'b1;  addr_rom[  541]='h00000874;  wr_data_rom[  541]='h0000224e;
    rd_cycle[  542] = 1'b0;  wr_cycle[  542] = 1'b1;  addr_rom[  542]='h00000878;  wr_data_rom[  542]='h00000761;
    rd_cycle[  543] = 1'b0;  wr_cycle[  543] = 1'b1;  addr_rom[  543]='h0000087c;  wr_data_rom[  543]='h0000273c;
    rd_cycle[  544] = 1'b0;  wr_cycle[  544] = 1'b1;  addr_rom[  544]='h00000880;  wr_data_rom[  544]='h0000182e;
    rd_cycle[  545] = 1'b0;  wr_cycle[  545] = 1'b1;  addr_rom[  545]='h00000884;  wr_data_rom[  545]='h000030e7;
    rd_cycle[  546] = 1'b0;  wr_cycle[  546] = 1'b1;  addr_rom[  546]='h00000888;  wr_data_rom[  546]='h00000132;
    rd_cycle[  547] = 1'b0;  wr_cycle[  547] = 1'b1;  addr_rom[  547]='h0000088c;  wr_data_rom[  547]='h0000233f;
    rd_cycle[  548] = 1'b0;  wr_cycle[  548] = 1'b1;  addr_rom[  548]='h00000890;  wr_data_rom[  548]='h00002170;
    rd_cycle[  549] = 1'b0;  wr_cycle[  549] = 1'b1;  addr_rom[  549]='h00000894;  wr_data_rom[  549]='h000014fa;
    rd_cycle[  550] = 1'b0;  wr_cycle[  550] = 1'b1;  addr_rom[  550]='h00000898;  wr_data_rom[  550]='h000037fc;
    rd_cycle[  551] = 1'b0;  wr_cycle[  551] = 1'b1;  addr_rom[  551]='h0000089c;  wr_data_rom[  551]='h00000ed8;
    rd_cycle[  552] = 1'b0;  wr_cycle[  552] = 1'b1;  addr_rom[  552]='h000008a0;  wr_data_rom[  552]='h000009c6;
    rd_cycle[  553] = 1'b0;  wr_cycle[  553] = 1'b1;  addr_rom[  553]='h000008a4;  wr_data_rom[  553]='h0000328d;
    rd_cycle[  554] = 1'b0;  wr_cycle[  554] = 1'b1;  addr_rom[  554]='h000008a8;  wr_data_rom[  554]='h00003ba5;
    rd_cycle[  555] = 1'b0;  wr_cycle[  555] = 1'b1;  addr_rom[  555]='h000008ac;  wr_data_rom[  555]='h00003174;
    rd_cycle[  556] = 1'b0;  wr_cycle[  556] = 1'b1;  addr_rom[  556]='h000008b0;  wr_data_rom[  556]='h00003126;
    rd_cycle[  557] = 1'b0;  wr_cycle[  557] = 1'b1;  addr_rom[  557]='h000008b4;  wr_data_rom[  557]='h000024fa;
    rd_cycle[  558] = 1'b0;  wr_cycle[  558] = 1'b1;  addr_rom[  558]='h000008b8;  wr_data_rom[  558]='h000018d8;
    rd_cycle[  559] = 1'b0;  wr_cycle[  559] = 1'b1;  addr_rom[  559]='h000008bc;  wr_data_rom[  559]='h000027cd;
    rd_cycle[  560] = 1'b0;  wr_cycle[  560] = 1'b1;  addr_rom[  560]='h000008c0;  wr_data_rom[  560]='h00003b9f;
    rd_cycle[  561] = 1'b0;  wr_cycle[  561] = 1'b1;  addr_rom[  561]='h000008c4;  wr_data_rom[  561]='h000031e7;
    rd_cycle[  562] = 1'b0;  wr_cycle[  562] = 1'b1;  addr_rom[  562]='h000008c8;  wr_data_rom[  562]='h00000fe6;
    rd_cycle[  563] = 1'b0;  wr_cycle[  563] = 1'b1;  addr_rom[  563]='h000008cc;  wr_data_rom[  563]='h00001ca9;
    rd_cycle[  564] = 1'b0;  wr_cycle[  564] = 1'b1;  addr_rom[  564]='h000008d0;  wr_data_rom[  564]='h00002a15;
    rd_cycle[  565] = 1'b0;  wr_cycle[  565] = 1'b1;  addr_rom[  565]='h000008d4;  wr_data_rom[  565]='h0000184e;
    rd_cycle[  566] = 1'b0;  wr_cycle[  566] = 1'b1;  addr_rom[  566]='h000008d8;  wr_data_rom[  566]='h00002c67;
    rd_cycle[  567] = 1'b0;  wr_cycle[  567] = 1'b1;  addr_rom[  567]='h000008dc;  wr_data_rom[  567]='h00001963;
    rd_cycle[  568] = 1'b0;  wr_cycle[  568] = 1'b1;  addr_rom[  568]='h000008e0;  wr_data_rom[  568]='h00001605;
    rd_cycle[  569] = 1'b0;  wr_cycle[  569] = 1'b1;  addr_rom[  569]='h000008e4;  wr_data_rom[  569]='h00000a4d;
    rd_cycle[  570] = 1'b0;  wr_cycle[  570] = 1'b1;  addr_rom[  570]='h000008e8;  wr_data_rom[  570]='h00001c73;
    rd_cycle[  571] = 1'b0;  wr_cycle[  571] = 1'b1;  addr_rom[  571]='h000008ec;  wr_data_rom[  571]='h00001a96;
    rd_cycle[  572] = 1'b0;  wr_cycle[  572] = 1'b1;  addr_rom[  572]='h000008f0;  wr_data_rom[  572]='h00002f38;
    rd_cycle[  573] = 1'b0;  wr_cycle[  573] = 1'b1;  addr_rom[  573]='h000008f4;  wr_data_rom[  573]='h00000f49;
    rd_cycle[  574] = 1'b0;  wr_cycle[  574] = 1'b1;  addr_rom[  574]='h000008f8;  wr_data_rom[  574]='h00000185;
    rd_cycle[  575] = 1'b0;  wr_cycle[  575] = 1'b1;  addr_rom[  575]='h000008fc;  wr_data_rom[  575]='h0000002c;
    rd_cycle[  576] = 1'b0;  wr_cycle[  576] = 1'b1;  addr_rom[  576]='h00000900;  wr_data_rom[  576]='h00001fb9;
    rd_cycle[  577] = 1'b0;  wr_cycle[  577] = 1'b1;  addr_rom[  577]='h00000904;  wr_data_rom[  577]='h0000145b;
    rd_cycle[  578] = 1'b0;  wr_cycle[  578] = 1'b1;  addr_rom[  578]='h00000908;  wr_data_rom[  578]='h00003527;
    rd_cycle[  579] = 1'b0;  wr_cycle[  579] = 1'b1;  addr_rom[  579]='h0000090c;  wr_data_rom[  579]='h00001ab7;
    rd_cycle[  580] = 1'b0;  wr_cycle[  580] = 1'b1;  addr_rom[  580]='h00000910;  wr_data_rom[  580]='h000008ee;
    rd_cycle[  581] = 1'b0;  wr_cycle[  581] = 1'b1;  addr_rom[  581]='h00000914;  wr_data_rom[  581]='h00000564;
    rd_cycle[  582] = 1'b0;  wr_cycle[  582] = 1'b1;  addr_rom[  582]='h00000918;  wr_data_rom[  582]='h0000055d;
    rd_cycle[  583] = 1'b0;  wr_cycle[  583] = 1'b1;  addr_rom[  583]='h0000091c;  wr_data_rom[  583]='h00002467;
    rd_cycle[  584] = 1'b0;  wr_cycle[  584] = 1'b1;  addr_rom[  584]='h00000920;  wr_data_rom[  584]='h00002689;
    rd_cycle[  585] = 1'b0;  wr_cycle[  585] = 1'b1;  addr_rom[  585]='h00000924;  wr_data_rom[  585]='h000027d1;
    rd_cycle[  586] = 1'b0;  wr_cycle[  586] = 1'b1;  addr_rom[  586]='h00000928;  wr_data_rom[  586]='h00003115;
    rd_cycle[  587] = 1'b0;  wr_cycle[  587] = 1'b1;  addr_rom[  587]='h0000092c;  wr_data_rom[  587]='h00002a28;
    rd_cycle[  588] = 1'b0;  wr_cycle[  588] = 1'b1;  addr_rom[  588]='h00000930;  wr_data_rom[  588]='h000000d0;
    rd_cycle[  589] = 1'b0;  wr_cycle[  589] = 1'b1;  addr_rom[  589]='h00000934;  wr_data_rom[  589]='h00000a7f;
    rd_cycle[  590] = 1'b0;  wr_cycle[  590] = 1'b1;  addr_rom[  590]='h00000938;  wr_data_rom[  590]='h000002f5;
    rd_cycle[  591] = 1'b0;  wr_cycle[  591] = 1'b1;  addr_rom[  591]='h0000093c;  wr_data_rom[  591]='h000037cb;
    rd_cycle[  592] = 1'b0;  wr_cycle[  592] = 1'b1;  addr_rom[  592]='h00000940;  wr_data_rom[  592]='h000021be;
    rd_cycle[  593] = 1'b0;  wr_cycle[  593] = 1'b1;  addr_rom[  593]='h00000944;  wr_data_rom[  593]='h0000017e;
    rd_cycle[  594] = 1'b0;  wr_cycle[  594] = 1'b1;  addr_rom[  594]='h00000948;  wr_data_rom[  594]='h00003fb4;
    rd_cycle[  595] = 1'b0;  wr_cycle[  595] = 1'b1;  addr_rom[  595]='h0000094c;  wr_data_rom[  595]='h000036e2;
    rd_cycle[  596] = 1'b0;  wr_cycle[  596] = 1'b1;  addr_rom[  596]='h00000950;  wr_data_rom[  596]='h00003415;
    rd_cycle[  597] = 1'b0;  wr_cycle[  597] = 1'b1;  addr_rom[  597]='h00000954;  wr_data_rom[  597]='h000037c5;
    rd_cycle[  598] = 1'b0;  wr_cycle[  598] = 1'b1;  addr_rom[  598]='h00000958;  wr_data_rom[  598]='h0000077d;
    rd_cycle[  599] = 1'b0;  wr_cycle[  599] = 1'b1;  addr_rom[  599]='h0000095c;  wr_data_rom[  599]='h00001593;
    rd_cycle[  600] = 1'b0;  wr_cycle[  600] = 1'b1;  addr_rom[  600]='h00000960;  wr_data_rom[  600]='h00002b62;
    rd_cycle[  601] = 1'b0;  wr_cycle[  601] = 1'b1;  addr_rom[  601]='h00000964;  wr_data_rom[  601]='h00002726;
    rd_cycle[  602] = 1'b0;  wr_cycle[  602] = 1'b1;  addr_rom[  602]='h00000968;  wr_data_rom[  602]='h00001711;
    rd_cycle[  603] = 1'b0;  wr_cycle[  603] = 1'b1;  addr_rom[  603]='h0000096c;  wr_data_rom[  603]='h00000b08;
    rd_cycle[  604] = 1'b0;  wr_cycle[  604] = 1'b1;  addr_rom[  604]='h00000970;  wr_data_rom[  604]='h0000011b;
    rd_cycle[  605] = 1'b0;  wr_cycle[  605] = 1'b1;  addr_rom[  605]='h00000974;  wr_data_rom[  605]='h00003817;
    rd_cycle[  606] = 1'b0;  wr_cycle[  606] = 1'b1;  addr_rom[  606]='h00000978;  wr_data_rom[  606]='h00002e91;
    rd_cycle[  607] = 1'b0;  wr_cycle[  607] = 1'b1;  addr_rom[  607]='h0000097c;  wr_data_rom[  607]='h00001219;
    rd_cycle[  608] = 1'b0;  wr_cycle[  608] = 1'b1;  addr_rom[  608]='h00000980;  wr_data_rom[  608]='h000005ce;
    rd_cycle[  609] = 1'b0;  wr_cycle[  609] = 1'b1;  addr_rom[  609]='h00000984;  wr_data_rom[  609]='h000006da;
    rd_cycle[  610] = 1'b0;  wr_cycle[  610] = 1'b1;  addr_rom[  610]='h00000988;  wr_data_rom[  610]='h00001f38;
    rd_cycle[  611] = 1'b0;  wr_cycle[  611] = 1'b1;  addr_rom[  611]='h0000098c;  wr_data_rom[  611]='h00002ccb;
    rd_cycle[  612] = 1'b0;  wr_cycle[  612] = 1'b1;  addr_rom[  612]='h00000990;  wr_data_rom[  612]='h0000103b;
    rd_cycle[  613] = 1'b0;  wr_cycle[  613] = 1'b1;  addr_rom[  613]='h00000994;  wr_data_rom[  613]='h00003123;
    rd_cycle[  614] = 1'b0;  wr_cycle[  614] = 1'b1;  addr_rom[  614]='h00000998;  wr_data_rom[  614]='h000024e7;
    rd_cycle[  615] = 1'b0;  wr_cycle[  615] = 1'b1;  addr_rom[  615]='h0000099c;  wr_data_rom[  615]='h00000e6b;
    rd_cycle[  616] = 1'b0;  wr_cycle[  616] = 1'b1;  addr_rom[  616]='h000009a0;  wr_data_rom[  616]='h00001d4e;
    rd_cycle[  617] = 1'b0;  wr_cycle[  617] = 1'b1;  addr_rom[  617]='h000009a4;  wr_data_rom[  617]='h000027de;
    rd_cycle[  618] = 1'b0;  wr_cycle[  618] = 1'b1;  addr_rom[  618]='h000009a8;  wr_data_rom[  618]='h00003fce;
    rd_cycle[  619] = 1'b0;  wr_cycle[  619] = 1'b1;  addr_rom[  619]='h000009ac;  wr_data_rom[  619]='h000028bc;
    rd_cycle[  620] = 1'b0;  wr_cycle[  620] = 1'b1;  addr_rom[  620]='h000009b0;  wr_data_rom[  620]='h0000356a;
    rd_cycle[  621] = 1'b0;  wr_cycle[  621] = 1'b1;  addr_rom[  621]='h000009b4;  wr_data_rom[  621]='h000026de;
    rd_cycle[  622] = 1'b0;  wr_cycle[  622] = 1'b1;  addr_rom[  622]='h000009b8;  wr_data_rom[  622]='h0000178e;
    rd_cycle[  623] = 1'b0;  wr_cycle[  623] = 1'b1;  addr_rom[  623]='h000009bc;  wr_data_rom[  623]='h0000106d;
    rd_cycle[  624] = 1'b0;  wr_cycle[  624] = 1'b1;  addr_rom[  624]='h000009c0;  wr_data_rom[  624]='h00002cd4;
    rd_cycle[  625] = 1'b0;  wr_cycle[  625] = 1'b1;  addr_rom[  625]='h000009c4;  wr_data_rom[  625]='h00000d1c;
    rd_cycle[  626] = 1'b0;  wr_cycle[  626] = 1'b1;  addr_rom[  626]='h000009c8;  wr_data_rom[  626]='h00003b4b;
    rd_cycle[  627] = 1'b0;  wr_cycle[  627] = 1'b1;  addr_rom[  627]='h000009cc;  wr_data_rom[  627]='h000006e2;
    rd_cycle[  628] = 1'b0;  wr_cycle[  628] = 1'b1;  addr_rom[  628]='h000009d0;  wr_data_rom[  628]='h00003260;
    rd_cycle[  629] = 1'b0;  wr_cycle[  629] = 1'b1;  addr_rom[  629]='h000009d4;  wr_data_rom[  629]='h0000314a;
    rd_cycle[  630] = 1'b0;  wr_cycle[  630] = 1'b1;  addr_rom[  630]='h000009d8;  wr_data_rom[  630]='h0000300c;
    rd_cycle[  631] = 1'b0;  wr_cycle[  631] = 1'b1;  addr_rom[  631]='h000009dc;  wr_data_rom[  631]='h00000264;
    rd_cycle[  632] = 1'b0;  wr_cycle[  632] = 1'b1;  addr_rom[  632]='h000009e0;  wr_data_rom[  632]='h00000022;
    rd_cycle[  633] = 1'b0;  wr_cycle[  633] = 1'b1;  addr_rom[  633]='h000009e4;  wr_data_rom[  633]='h00001905;
    rd_cycle[  634] = 1'b0;  wr_cycle[  634] = 1'b1;  addr_rom[  634]='h000009e8;  wr_data_rom[  634]='h00001c69;
    rd_cycle[  635] = 1'b0;  wr_cycle[  635] = 1'b1;  addr_rom[  635]='h000009ec;  wr_data_rom[  635]='h00003173;
    rd_cycle[  636] = 1'b0;  wr_cycle[  636] = 1'b1;  addr_rom[  636]='h000009f0;  wr_data_rom[  636]='h0000346e;
    rd_cycle[  637] = 1'b0;  wr_cycle[  637] = 1'b1;  addr_rom[  637]='h000009f4;  wr_data_rom[  637]='h000008a9;
    rd_cycle[  638] = 1'b0;  wr_cycle[  638] = 1'b1;  addr_rom[  638]='h000009f8;  wr_data_rom[  638]='h00000ff8;
    rd_cycle[  639] = 1'b0;  wr_cycle[  639] = 1'b1;  addr_rom[  639]='h000009fc;  wr_data_rom[  639]='h00003309;
    rd_cycle[  640] = 1'b0;  wr_cycle[  640] = 1'b1;  addr_rom[  640]='h00000a00;  wr_data_rom[  640]='h000020a9;
    rd_cycle[  641] = 1'b0;  wr_cycle[  641] = 1'b1;  addr_rom[  641]='h00000a04;  wr_data_rom[  641]='h00001d18;
    rd_cycle[  642] = 1'b0;  wr_cycle[  642] = 1'b1;  addr_rom[  642]='h00000a08;  wr_data_rom[  642]='h00001a5a;
    rd_cycle[  643] = 1'b0;  wr_cycle[  643] = 1'b1;  addr_rom[  643]='h00000a0c;  wr_data_rom[  643]='h00003a32;
    rd_cycle[  644] = 1'b0;  wr_cycle[  644] = 1'b1;  addr_rom[  644]='h00000a10;  wr_data_rom[  644]='h00001a2d;
    rd_cycle[  645] = 1'b0;  wr_cycle[  645] = 1'b1;  addr_rom[  645]='h00000a14;  wr_data_rom[  645]='h000018f3;
    rd_cycle[  646] = 1'b0;  wr_cycle[  646] = 1'b1;  addr_rom[  646]='h00000a18;  wr_data_rom[  646]='h000001eb;
    rd_cycle[  647] = 1'b0;  wr_cycle[  647] = 1'b1;  addr_rom[  647]='h00000a1c;  wr_data_rom[  647]='h00001ff7;
    rd_cycle[  648] = 1'b0;  wr_cycle[  648] = 1'b1;  addr_rom[  648]='h00000a20;  wr_data_rom[  648]='h0000319e;
    rd_cycle[  649] = 1'b0;  wr_cycle[  649] = 1'b1;  addr_rom[  649]='h00000a24;  wr_data_rom[  649]='h000003f4;
    rd_cycle[  650] = 1'b0;  wr_cycle[  650] = 1'b1;  addr_rom[  650]='h00000a28;  wr_data_rom[  650]='h00001e7f;
    rd_cycle[  651] = 1'b0;  wr_cycle[  651] = 1'b1;  addr_rom[  651]='h00000a2c;  wr_data_rom[  651]='h00002a34;
    rd_cycle[  652] = 1'b0;  wr_cycle[  652] = 1'b1;  addr_rom[  652]='h00000a30;  wr_data_rom[  652]='h00001eb2;
    rd_cycle[  653] = 1'b0;  wr_cycle[  653] = 1'b1;  addr_rom[  653]='h00000a34;  wr_data_rom[  653]='h0000007c;
    rd_cycle[  654] = 1'b0;  wr_cycle[  654] = 1'b1;  addr_rom[  654]='h00000a38;  wr_data_rom[  654]='h000022b0;
    rd_cycle[  655] = 1'b0;  wr_cycle[  655] = 1'b1;  addr_rom[  655]='h00000a3c;  wr_data_rom[  655]='h00000bba;
    rd_cycle[  656] = 1'b0;  wr_cycle[  656] = 1'b1;  addr_rom[  656]='h00000a40;  wr_data_rom[  656]='h00000f65;
    rd_cycle[  657] = 1'b0;  wr_cycle[  657] = 1'b1;  addr_rom[  657]='h00000a44;  wr_data_rom[  657]='h00001694;
    rd_cycle[  658] = 1'b0;  wr_cycle[  658] = 1'b1;  addr_rom[  658]='h00000a48;  wr_data_rom[  658]='h00000b25;
    rd_cycle[  659] = 1'b0;  wr_cycle[  659] = 1'b1;  addr_rom[  659]='h00000a4c;  wr_data_rom[  659]='h00002175;
    rd_cycle[  660] = 1'b0;  wr_cycle[  660] = 1'b1;  addr_rom[  660]='h00000a50;  wr_data_rom[  660]='h00000991;
    rd_cycle[  661] = 1'b0;  wr_cycle[  661] = 1'b1;  addr_rom[  661]='h00000a54;  wr_data_rom[  661]='h00000ecc;
    rd_cycle[  662] = 1'b0;  wr_cycle[  662] = 1'b1;  addr_rom[  662]='h00000a58;  wr_data_rom[  662]='h000035c0;
    rd_cycle[  663] = 1'b0;  wr_cycle[  663] = 1'b1;  addr_rom[  663]='h00000a5c;  wr_data_rom[  663]='h00003738;
    rd_cycle[  664] = 1'b0;  wr_cycle[  664] = 1'b1;  addr_rom[  664]='h00000a60;  wr_data_rom[  664]='h00001a33;
    rd_cycle[  665] = 1'b0;  wr_cycle[  665] = 1'b1;  addr_rom[  665]='h00000a64;  wr_data_rom[  665]='h00002958;
    rd_cycle[  666] = 1'b0;  wr_cycle[  666] = 1'b1;  addr_rom[  666]='h00000a68;  wr_data_rom[  666]='h00002c84;
    rd_cycle[  667] = 1'b0;  wr_cycle[  667] = 1'b1;  addr_rom[  667]='h00000a6c;  wr_data_rom[  667]='h00000645;
    rd_cycle[  668] = 1'b0;  wr_cycle[  668] = 1'b1;  addr_rom[  668]='h00000a70;  wr_data_rom[  668]='h00002927;
    rd_cycle[  669] = 1'b0;  wr_cycle[  669] = 1'b1;  addr_rom[  669]='h00000a74;  wr_data_rom[  669]='h00001087;
    rd_cycle[  670] = 1'b0;  wr_cycle[  670] = 1'b1;  addr_rom[  670]='h00000a78;  wr_data_rom[  670]='h00000ab1;
    rd_cycle[  671] = 1'b0;  wr_cycle[  671] = 1'b1;  addr_rom[  671]='h00000a7c;  wr_data_rom[  671]='h000020de;
    rd_cycle[  672] = 1'b0;  wr_cycle[  672] = 1'b1;  addr_rom[  672]='h00000a80;  wr_data_rom[  672]='h00002e28;
    rd_cycle[  673] = 1'b0;  wr_cycle[  673] = 1'b1;  addr_rom[  673]='h00000a84;  wr_data_rom[  673]='h00001b0e;
    rd_cycle[  674] = 1'b0;  wr_cycle[  674] = 1'b1;  addr_rom[  674]='h00000a88;  wr_data_rom[  674]='h00002859;
    rd_cycle[  675] = 1'b0;  wr_cycle[  675] = 1'b1;  addr_rom[  675]='h00000a8c;  wr_data_rom[  675]='h0000031f;
    rd_cycle[  676] = 1'b0;  wr_cycle[  676] = 1'b1;  addr_rom[  676]='h00000a90;  wr_data_rom[  676]='h000017f6;
    rd_cycle[  677] = 1'b0;  wr_cycle[  677] = 1'b1;  addr_rom[  677]='h00000a94;  wr_data_rom[  677]='h00000cdd;
    rd_cycle[  678] = 1'b0;  wr_cycle[  678] = 1'b1;  addr_rom[  678]='h00000a98;  wr_data_rom[  678]='h000023b8;
    rd_cycle[  679] = 1'b0;  wr_cycle[  679] = 1'b1;  addr_rom[  679]='h00000a9c;  wr_data_rom[  679]='h00001173;
    rd_cycle[  680] = 1'b0;  wr_cycle[  680] = 1'b1;  addr_rom[  680]='h00000aa0;  wr_data_rom[  680]='h00002d2b;
    rd_cycle[  681] = 1'b0;  wr_cycle[  681] = 1'b1;  addr_rom[  681]='h00000aa4;  wr_data_rom[  681]='h00000eca;
    rd_cycle[  682] = 1'b0;  wr_cycle[  682] = 1'b1;  addr_rom[  682]='h00000aa8;  wr_data_rom[  682]='h00001391;
    rd_cycle[  683] = 1'b0;  wr_cycle[  683] = 1'b1;  addr_rom[  683]='h00000aac;  wr_data_rom[  683]='h00002af3;
    rd_cycle[  684] = 1'b0;  wr_cycle[  684] = 1'b1;  addr_rom[  684]='h00000ab0;  wr_data_rom[  684]='h00001957;
    rd_cycle[  685] = 1'b0;  wr_cycle[  685] = 1'b1;  addr_rom[  685]='h00000ab4;  wr_data_rom[  685]='h000038c6;
    rd_cycle[  686] = 1'b0;  wr_cycle[  686] = 1'b1;  addr_rom[  686]='h00000ab8;  wr_data_rom[  686]='h00001e0c;
    rd_cycle[  687] = 1'b0;  wr_cycle[  687] = 1'b1;  addr_rom[  687]='h00000abc;  wr_data_rom[  687]='h00003960;
    rd_cycle[  688] = 1'b0;  wr_cycle[  688] = 1'b1;  addr_rom[  688]='h00000ac0;  wr_data_rom[  688]='h00002d9c;
    rd_cycle[  689] = 1'b0;  wr_cycle[  689] = 1'b1;  addr_rom[  689]='h00000ac4;  wr_data_rom[  689]='h0000244d;
    rd_cycle[  690] = 1'b0;  wr_cycle[  690] = 1'b1;  addr_rom[  690]='h00000ac8;  wr_data_rom[  690]='h00001899;
    rd_cycle[  691] = 1'b0;  wr_cycle[  691] = 1'b1;  addr_rom[  691]='h00000acc;  wr_data_rom[  691]='h00000787;
    rd_cycle[  692] = 1'b0;  wr_cycle[  692] = 1'b1;  addr_rom[  692]='h00000ad0;  wr_data_rom[  692]='h00001aa9;
    rd_cycle[  693] = 1'b0;  wr_cycle[  693] = 1'b1;  addr_rom[  693]='h00000ad4;  wr_data_rom[  693]='h0000043a;
    rd_cycle[  694] = 1'b0;  wr_cycle[  694] = 1'b1;  addr_rom[  694]='h00000ad8;  wr_data_rom[  694]='h00002c71;
    rd_cycle[  695] = 1'b0;  wr_cycle[  695] = 1'b1;  addr_rom[  695]='h00000adc;  wr_data_rom[  695]='h00001ffc;
    rd_cycle[  696] = 1'b0;  wr_cycle[  696] = 1'b1;  addr_rom[  696]='h00000ae0;  wr_data_rom[  696]='h00000fbf;
    rd_cycle[  697] = 1'b0;  wr_cycle[  697] = 1'b1;  addr_rom[  697]='h00000ae4;  wr_data_rom[  697]='h00001952;
    rd_cycle[  698] = 1'b0;  wr_cycle[  698] = 1'b1;  addr_rom[  698]='h00000ae8;  wr_data_rom[  698]='h00003594;
    rd_cycle[  699] = 1'b0;  wr_cycle[  699] = 1'b1;  addr_rom[  699]='h00000aec;  wr_data_rom[  699]='h000034ad;
    rd_cycle[  700] = 1'b0;  wr_cycle[  700] = 1'b1;  addr_rom[  700]='h00000af0;  wr_data_rom[  700]='h00001841;
    rd_cycle[  701] = 1'b0;  wr_cycle[  701] = 1'b1;  addr_rom[  701]='h00000af4;  wr_data_rom[  701]='h00003537;
    rd_cycle[  702] = 1'b0;  wr_cycle[  702] = 1'b1;  addr_rom[  702]='h00000af8;  wr_data_rom[  702]='h00000076;
    rd_cycle[  703] = 1'b0;  wr_cycle[  703] = 1'b1;  addr_rom[  703]='h00000afc;  wr_data_rom[  703]='h00000df3;
    rd_cycle[  704] = 1'b0;  wr_cycle[  704] = 1'b1;  addr_rom[  704]='h00000b00;  wr_data_rom[  704]='h000023b2;
    rd_cycle[  705] = 1'b0;  wr_cycle[  705] = 1'b1;  addr_rom[  705]='h00000b04;  wr_data_rom[  705]='h000013f7;
    rd_cycle[  706] = 1'b0;  wr_cycle[  706] = 1'b1;  addr_rom[  706]='h00000b08;  wr_data_rom[  706]='h00000d60;
    rd_cycle[  707] = 1'b0;  wr_cycle[  707] = 1'b1;  addr_rom[  707]='h00000b0c;  wr_data_rom[  707]='h00002a76;
    rd_cycle[  708] = 1'b0;  wr_cycle[  708] = 1'b1;  addr_rom[  708]='h00000b10;  wr_data_rom[  708]='h0000035b;
    rd_cycle[  709] = 1'b0;  wr_cycle[  709] = 1'b1;  addr_rom[  709]='h00000b14;  wr_data_rom[  709]='h00000bf5;
    rd_cycle[  710] = 1'b0;  wr_cycle[  710] = 1'b1;  addr_rom[  710]='h00000b18;  wr_data_rom[  710]='h00003974;
    rd_cycle[  711] = 1'b0;  wr_cycle[  711] = 1'b1;  addr_rom[  711]='h00000b1c;  wr_data_rom[  711]='h00000a9b;
    rd_cycle[  712] = 1'b0;  wr_cycle[  712] = 1'b1;  addr_rom[  712]='h00000b20;  wr_data_rom[  712]='h0000250f;
    rd_cycle[  713] = 1'b0;  wr_cycle[  713] = 1'b1;  addr_rom[  713]='h00000b24;  wr_data_rom[  713]='h00001b01;
    rd_cycle[  714] = 1'b0;  wr_cycle[  714] = 1'b1;  addr_rom[  714]='h00000b28;  wr_data_rom[  714]='h00000df5;
    rd_cycle[  715] = 1'b0;  wr_cycle[  715] = 1'b1;  addr_rom[  715]='h00000b2c;  wr_data_rom[  715]='h00002a6e;
    rd_cycle[  716] = 1'b0;  wr_cycle[  716] = 1'b1;  addr_rom[  716]='h00000b30;  wr_data_rom[  716]='h0000255a;
    rd_cycle[  717] = 1'b0;  wr_cycle[  717] = 1'b1;  addr_rom[  717]='h00000b34;  wr_data_rom[  717]='h000016f1;
    rd_cycle[  718] = 1'b0;  wr_cycle[  718] = 1'b1;  addr_rom[  718]='h00000b38;  wr_data_rom[  718]='h00000f59;
    rd_cycle[  719] = 1'b0;  wr_cycle[  719] = 1'b1;  addr_rom[  719]='h00000b3c;  wr_data_rom[  719]='h000009d0;
    rd_cycle[  720] = 1'b0;  wr_cycle[  720] = 1'b1;  addr_rom[  720]='h00000b40;  wr_data_rom[  720]='h00000f71;
    rd_cycle[  721] = 1'b0;  wr_cycle[  721] = 1'b1;  addr_rom[  721]='h00000b44;  wr_data_rom[  721]='h00000376;
    rd_cycle[  722] = 1'b0;  wr_cycle[  722] = 1'b1;  addr_rom[  722]='h00000b48;  wr_data_rom[  722]='h00003977;
    rd_cycle[  723] = 1'b0;  wr_cycle[  723] = 1'b1;  addr_rom[  723]='h00000b4c;  wr_data_rom[  723]='h000006b5;
    rd_cycle[  724] = 1'b0;  wr_cycle[  724] = 1'b1;  addr_rom[  724]='h00000b50;  wr_data_rom[  724]='h00001ae7;
    rd_cycle[  725] = 1'b0;  wr_cycle[  725] = 1'b1;  addr_rom[  725]='h00000b54;  wr_data_rom[  725]='h00001b3a;
    rd_cycle[  726] = 1'b0;  wr_cycle[  726] = 1'b1;  addr_rom[  726]='h00000b58;  wr_data_rom[  726]='h00001aa5;
    rd_cycle[  727] = 1'b0;  wr_cycle[  727] = 1'b1;  addr_rom[  727]='h00000b5c;  wr_data_rom[  727]='h00001fd0;
    rd_cycle[  728] = 1'b0;  wr_cycle[  728] = 1'b1;  addr_rom[  728]='h00000b60;  wr_data_rom[  728]='h000009b0;
    rd_cycle[  729] = 1'b0;  wr_cycle[  729] = 1'b1;  addr_rom[  729]='h00000b64;  wr_data_rom[  729]='h00000a4f;
    rd_cycle[  730] = 1'b0;  wr_cycle[  730] = 1'b1;  addr_rom[  730]='h00000b68;  wr_data_rom[  730]='h0000163f;
    rd_cycle[  731] = 1'b0;  wr_cycle[  731] = 1'b1;  addr_rom[  731]='h00000b6c;  wr_data_rom[  731]='h00000097;
    rd_cycle[  732] = 1'b0;  wr_cycle[  732] = 1'b1;  addr_rom[  732]='h00000b70;  wr_data_rom[  732]='h00000121;
    rd_cycle[  733] = 1'b0;  wr_cycle[  733] = 1'b1;  addr_rom[  733]='h00000b74;  wr_data_rom[  733]='h00002704;
    rd_cycle[  734] = 1'b0;  wr_cycle[  734] = 1'b1;  addr_rom[  734]='h00000b78;  wr_data_rom[  734]='h000012e3;
    rd_cycle[  735] = 1'b0;  wr_cycle[  735] = 1'b1;  addr_rom[  735]='h00000b7c;  wr_data_rom[  735]='h000000f4;
    rd_cycle[  736] = 1'b0;  wr_cycle[  736] = 1'b1;  addr_rom[  736]='h00000b80;  wr_data_rom[  736]='h00000195;
    rd_cycle[  737] = 1'b0;  wr_cycle[  737] = 1'b1;  addr_rom[  737]='h00000b84;  wr_data_rom[  737]='h00002ae3;
    rd_cycle[  738] = 1'b0;  wr_cycle[  738] = 1'b1;  addr_rom[  738]='h00000b88;  wr_data_rom[  738]='h00003cfe;
    rd_cycle[  739] = 1'b0;  wr_cycle[  739] = 1'b1;  addr_rom[  739]='h00000b8c;  wr_data_rom[  739]='h000039df;
    rd_cycle[  740] = 1'b0;  wr_cycle[  740] = 1'b1;  addr_rom[  740]='h00000b90;  wr_data_rom[  740]='h0000068e;
    rd_cycle[  741] = 1'b0;  wr_cycle[  741] = 1'b1;  addr_rom[  741]='h00000b94;  wr_data_rom[  741]='h000023f9;
    rd_cycle[  742] = 1'b0;  wr_cycle[  742] = 1'b1;  addr_rom[  742]='h00000b98;  wr_data_rom[  742]='h000019cc;
    rd_cycle[  743] = 1'b0;  wr_cycle[  743] = 1'b1;  addr_rom[  743]='h00000b9c;  wr_data_rom[  743]='h00003a77;
    rd_cycle[  744] = 1'b0;  wr_cycle[  744] = 1'b1;  addr_rom[  744]='h00000ba0;  wr_data_rom[  744]='h00003fdf;
    rd_cycle[  745] = 1'b0;  wr_cycle[  745] = 1'b1;  addr_rom[  745]='h00000ba4;  wr_data_rom[  745]='h00002ca7;
    rd_cycle[  746] = 1'b0;  wr_cycle[  746] = 1'b1;  addr_rom[  746]='h00000ba8;  wr_data_rom[  746]='h00000ee3;
    rd_cycle[  747] = 1'b0;  wr_cycle[  747] = 1'b1;  addr_rom[  747]='h00000bac;  wr_data_rom[  747]='h00001cc5;
    rd_cycle[  748] = 1'b0;  wr_cycle[  748] = 1'b1;  addr_rom[  748]='h00000bb0;  wr_data_rom[  748]='h00000b33;
    rd_cycle[  749] = 1'b0;  wr_cycle[  749] = 1'b1;  addr_rom[  749]='h00000bb4;  wr_data_rom[  749]='h00002196;
    rd_cycle[  750] = 1'b0;  wr_cycle[  750] = 1'b1;  addr_rom[  750]='h00000bb8;  wr_data_rom[  750]='h0000054d;
    rd_cycle[  751] = 1'b0;  wr_cycle[  751] = 1'b1;  addr_rom[  751]='h00000bbc;  wr_data_rom[  751]='h00002241;
    rd_cycle[  752] = 1'b0;  wr_cycle[  752] = 1'b1;  addr_rom[  752]='h00000bc0;  wr_data_rom[  752]='h00001c0e;
    rd_cycle[  753] = 1'b0;  wr_cycle[  753] = 1'b1;  addr_rom[  753]='h00000bc4;  wr_data_rom[  753]='h000023bf;
    rd_cycle[  754] = 1'b0;  wr_cycle[  754] = 1'b1;  addr_rom[  754]='h00000bc8;  wr_data_rom[  754]='h00000e11;
    rd_cycle[  755] = 1'b0;  wr_cycle[  755] = 1'b1;  addr_rom[  755]='h00000bcc;  wr_data_rom[  755]='h00002ec7;
    rd_cycle[  756] = 1'b0;  wr_cycle[  756] = 1'b1;  addr_rom[  756]='h00000bd0;  wr_data_rom[  756]='h000037a1;
    rd_cycle[  757] = 1'b0;  wr_cycle[  757] = 1'b1;  addr_rom[  757]='h00000bd4;  wr_data_rom[  757]='h000029e3;
    rd_cycle[  758] = 1'b0;  wr_cycle[  758] = 1'b1;  addr_rom[  758]='h00000bd8;  wr_data_rom[  758]='h00003d61;
    rd_cycle[  759] = 1'b0;  wr_cycle[  759] = 1'b1;  addr_rom[  759]='h00000bdc;  wr_data_rom[  759]='h00003004;
    rd_cycle[  760] = 1'b0;  wr_cycle[  760] = 1'b1;  addr_rom[  760]='h00000be0;  wr_data_rom[  760]='h00001a0e;
    rd_cycle[  761] = 1'b0;  wr_cycle[  761] = 1'b1;  addr_rom[  761]='h00000be4;  wr_data_rom[  761]='h000013b0;
    rd_cycle[  762] = 1'b0;  wr_cycle[  762] = 1'b1;  addr_rom[  762]='h00000be8;  wr_data_rom[  762]='h00003e5b;
    rd_cycle[  763] = 1'b0;  wr_cycle[  763] = 1'b1;  addr_rom[  763]='h00000bec;  wr_data_rom[  763]='h000018a9;
    rd_cycle[  764] = 1'b0;  wr_cycle[  764] = 1'b1;  addr_rom[  764]='h00000bf0;  wr_data_rom[  764]='h00001b09;
    rd_cycle[  765] = 1'b0;  wr_cycle[  765] = 1'b1;  addr_rom[  765]='h00000bf4;  wr_data_rom[  765]='h00001764;
    rd_cycle[  766] = 1'b0;  wr_cycle[  766] = 1'b1;  addr_rom[  766]='h00000bf8;  wr_data_rom[  766]='h00003f75;
    rd_cycle[  767] = 1'b0;  wr_cycle[  767] = 1'b1;  addr_rom[  767]='h00000bfc;  wr_data_rom[  767]='h00001d44;
    rd_cycle[  768] = 1'b0;  wr_cycle[  768] = 1'b1;  addr_rom[  768]='h00000c00;  wr_data_rom[  768]='h000029b1;
    rd_cycle[  769] = 1'b0;  wr_cycle[  769] = 1'b1;  addr_rom[  769]='h00000c04;  wr_data_rom[  769]='h00002206;
    rd_cycle[  770] = 1'b0;  wr_cycle[  770] = 1'b1;  addr_rom[  770]='h00000c08;  wr_data_rom[  770]='h00003a70;
    rd_cycle[  771] = 1'b0;  wr_cycle[  771] = 1'b1;  addr_rom[  771]='h00000c0c;  wr_data_rom[  771]='h000029d6;
    rd_cycle[  772] = 1'b0;  wr_cycle[  772] = 1'b1;  addr_rom[  772]='h00000c10;  wr_data_rom[  772]='h00001a26;
    rd_cycle[  773] = 1'b0;  wr_cycle[  773] = 1'b1;  addr_rom[  773]='h00000c14;  wr_data_rom[  773]='h0000232a;
    rd_cycle[  774] = 1'b0;  wr_cycle[  774] = 1'b1;  addr_rom[  774]='h00000c18;  wr_data_rom[  774]='h00001876;
    rd_cycle[  775] = 1'b0;  wr_cycle[  775] = 1'b1;  addr_rom[  775]='h00000c1c;  wr_data_rom[  775]='h00002403;
    rd_cycle[  776] = 1'b0;  wr_cycle[  776] = 1'b1;  addr_rom[  776]='h00000c20;  wr_data_rom[  776]='h00003eff;
    rd_cycle[  777] = 1'b0;  wr_cycle[  777] = 1'b1;  addr_rom[  777]='h00000c24;  wr_data_rom[  777]='h00001ae3;
    rd_cycle[  778] = 1'b0;  wr_cycle[  778] = 1'b1;  addr_rom[  778]='h00000c28;  wr_data_rom[  778]='h000023a2;
    rd_cycle[  779] = 1'b0;  wr_cycle[  779] = 1'b1;  addr_rom[  779]='h00000c2c;  wr_data_rom[  779]='h00000e08;
    rd_cycle[  780] = 1'b0;  wr_cycle[  780] = 1'b1;  addr_rom[  780]='h00000c30;  wr_data_rom[  780]='h0000279a;
    rd_cycle[  781] = 1'b0;  wr_cycle[  781] = 1'b1;  addr_rom[  781]='h00000c34;  wr_data_rom[  781]='h00001b47;
    rd_cycle[  782] = 1'b0;  wr_cycle[  782] = 1'b1;  addr_rom[  782]='h00000c38;  wr_data_rom[  782]='h0000392f;
    rd_cycle[  783] = 1'b0;  wr_cycle[  783] = 1'b1;  addr_rom[  783]='h00000c3c;  wr_data_rom[  783]='h00002956;
    rd_cycle[  784] = 1'b0;  wr_cycle[  784] = 1'b1;  addr_rom[  784]='h00000c40;  wr_data_rom[  784]='h00001a81;
    rd_cycle[  785] = 1'b0;  wr_cycle[  785] = 1'b1;  addr_rom[  785]='h00000c44;  wr_data_rom[  785]='h000017bd;
    rd_cycle[  786] = 1'b0;  wr_cycle[  786] = 1'b1;  addr_rom[  786]='h00000c48;  wr_data_rom[  786]='h0000038f;
    rd_cycle[  787] = 1'b0;  wr_cycle[  787] = 1'b1;  addr_rom[  787]='h00000c4c;  wr_data_rom[  787]='h000005f4;
    rd_cycle[  788] = 1'b0;  wr_cycle[  788] = 1'b1;  addr_rom[  788]='h00000c50;  wr_data_rom[  788]='h0000299e;
    rd_cycle[  789] = 1'b0;  wr_cycle[  789] = 1'b1;  addr_rom[  789]='h00000c54;  wr_data_rom[  789]='h00001728;
    rd_cycle[  790] = 1'b0;  wr_cycle[  790] = 1'b1;  addr_rom[  790]='h00000c58;  wr_data_rom[  790]='h0000072f;
    rd_cycle[  791] = 1'b0;  wr_cycle[  791] = 1'b1;  addr_rom[  791]='h00000c5c;  wr_data_rom[  791]='h00002324;
    rd_cycle[  792] = 1'b0;  wr_cycle[  792] = 1'b1;  addr_rom[  792]='h00000c60;  wr_data_rom[  792]='h00000c28;
    rd_cycle[  793] = 1'b0;  wr_cycle[  793] = 1'b1;  addr_rom[  793]='h00000c64;  wr_data_rom[  793]='h00000627;
    rd_cycle[  794] = 1'b0;  wr_cycle[  794] = 1'b1;  addr_rom[  794]='h00000c68;  wr_data_rom[  794]='h0000279a;
    rd_cycle[  795] = 1'b0;  wr_cycle[  795] = 1'b1;  addr_rom[  795]='h00000c6c;  wr_data_rom[  795]='h00002d14;
    rd_cycle[  796] = 1'b0;  wr_cycle[  796] = 1'b1;  addr_rom[  796]='h00000c70;  wr_data_rom[  796]='h0000261d;
    rd_cycle[  797] = 1'b0;  wr_cycle[  797] = 1'b1;  addr_rom[  797]='h00000c74;  wr_data_rom[  797]='h00000279;
    rd_cycle[  798] = 1'b0;  wr_cycle[  798] = 1'b1;  addr_rom[  798]='h00000c78;  wr_data_rom[  798]='h00001c96;
    rd_cycle[  799] = 1'b0;  wr_cycle[  799] = 1'b1;  addr_rom[  799]='h00000c7c;  wr_data_rom[  799]='h00003b83;
    rd_cycle[  800] = 1'b0;  wr_cycle[  800] = 1'b1;  addr_rom[  800]='h00000c80;  wr_data_rom[  800]='h0000177e;
    rd_cycle[  801] = 1'b0;  wr_cycle[  801] = 1'b1;  addr_rom[  801]='h00000c84;  wr_data_rom[  801]='h00001acc;
    rd_cycle[  802] = 1'b0;  wr_cycle[  802] = 1'b1;  addr_rom[  802]='h00000c88;  wr_data_rom[  802]='h000007fa;
    rd_cycle[  803] = 1'b0;  wr_cycle[  803] = 1'b1;  addr_rom[  803]='h00000c8c;  wr_data_rom[  803]='h000012d7;
    rd_cycle[  804] = 1'b0;  wr_cycle[  804] = 1'b1;  addr_rom[  804]='h00000c90;  wr_data_rom[  804]='h0000112e;
    rd_cycle[  805] = 1'b0;  wr_cycle[  805] = 1'b1;  addr_rom[  805]='h00000c94;  wr_data_rom[  805]='h0000030a;
    rd_cycle[  806] = 1'b0;  wr_cycle[  806] = 1'b1;  addr_rom[  806]='h00000c98;  wr_data_rom[  806]='h00003d25;
    rd_cycle[  807] = 1'b0;  wr_cycle[  807] = 1'b1;  addr_rom[  807]='h00000c9c;  wr_data_rom[  807]='h00001b28;
    rd_cycle[  808] = 1'b0;  wr_cycle[  808] = 1'b1;  addr_rom[  808]='h00000ca0;  wr_data_rom[  808]='h0000005e;
    rd_cycle[  809] = 1'b0;  wr_cycle[  809] = 1'b1;  addr_rom[  809]='h00000ca4;  wr_data_rom[  809]='h0000371b;
    rd_cycle[  810] = 1'b0;  wr_cycle[  810] = 1'b1;  addr_rom[  810]='h00000ca8;  wr_data_rom[  810]='h0000180a;
    rd_cycle[  811] = 1'b0;  wr_cycle[  811] = 1'b1;  addr_rom[  811]='h00000cac;  wr_data_rom[  811]='h00000b02;
    rd_cycle[  812] = 1'b0;  wr_cycle[  812] = 1'b1;  addr_rom[  812]='h00000cb0;  wr_data_rom[  812]='h00001be2;
    rd_cycle[  813] = 1'b0;  wr_cycle[  813] = 1'b1;  addr_rom[  813]='h00000cb4;  wr_data_rom[  813]='h000018d9;
    rd_cycle[  814] = 1'b0;  wr_cycle[  814] = 1'b1;  addr_rom[  814]='h00000cb8;  wr_data_rom[  814]='h0000269a;
    rd_cycle[  815] = 1'b0;  wr_cycle[  815] = 1'b1;  addr_rom[  815]='h00000cbc;  wr_data_rom[  815]='h000019fd;
    rd_cycle[  816] = 1'b0;  wr_cycle[  816] = 1'b1;  addr_rom[  816]='h00000cc0;  wr_data_rom[  816]='h0000337f;
    rd_cycle[  817] = 1'b0;  wr_cycle[  817] = 1'b1;  addr_rom[  817]='h00000cc4;  wr_data_rom[  817]='h00002944;
    rd_cycle[  818] = 1'b0;  wr_cycle[  818] = 1'b1;  addr_rom[  818]='h00000cc8;  wr_data_rom[  818]='h00002802;
    rd_cycle[  819] = 1'b0;  wr_cycle[  819] = 1'b1;  addr_rom[  819]='h00000ccc;  wr_data_rom[  819]='h00001bc3;
    rd_cycle[  820] = 1'b0;  wr_cycle[  820] = 1'b1;  addr_rom[  820]='h00000cd0;  wr_data_rom[  820]='h000023fa;
    rd_cycle[  821] = 1'b0;  wr_cycle[  821] = 1'b1;  addr_rom[  821]='h00000cd4;  wr_data_rom[  821]='h000038a7;
    rd_cycle[  822] = 1'b0;  wr_cycle[  822] = 1'b1;  addr_rom[  822]='h00000cd8;  wr_data_rom[  822]='h00001f2a;
    rd_cycle[  823] = 1'b0;  wr_cycle[  823] = 1'b1;  addr_rom[  823]='h00000cdc;  wr_data_rom[  823]='h00002ab3;
    rd_cycle[  824] = 1'b0;  wr_cycle[  824] = 1'b1;  addr_rom[  824]='h00000ce0;  wr_data_rom[  824]='h000030cc;
    rd_cycle[  825] = 1'b0;  wr_cycle[  825] = 1'b1;  addr_rom[  825]='h00000ce4;  wr_data_rom[  825]='h00003429;
    rd_cycle[  826] = 1'b0;  wr_cycle[  826] = 1'b1;  addr_rom[  826]='h00000ce8;  wr_data_rom[  826]='h00002bf8;
    rd_cycle[  827] = 1'b0;  wr_cycle[  827] = 1'b1;  addr_rom[  827]='h00000cec;  wr_data_rom[  827]='h0000050a;
    rd_cycle[  828] = 1'b0;  wr_cycle[  828] = 1'b1;  addr_rom[  828]='h00000cf0;  wr_data_rom[  828]='h00002181;
    rd_cycle[  829] = 1'b0;  wr_cycle[  829] = 1'b1;  addr_rom[  829]='h00000cf4;  wr_data_rom[  829]='h000014a7;
    rd_cycle[  830] = 1'b0;  wr_cycle[  830] = 1'b1;  addr_rom[  830]='h00000cf8;  wr_data_rom[  830]='h00003d91;
    rd_cycle[  831] = 1'b0;  wr_cycle[  831] = 1'b1;  addr_rom[  831]='h00000cfc;  wr_data_rom[  831]='h00001d0a;
    rd_cycle[  832] = 1'b0;  wr_cycle[  832] = 1'b1;  addr_rom[  832]='h00000d00;  wr_data_rom[  832]='h000004e4;
    rd_cycle[  833] = 1'b0;  wr_cycle[  833] = 1'b1;  addr_rom[  833]='h00000d04;  wr_data_rom[  833]='h00000d96;
    rd_cycle[  834] = 1'b0;  wr_cycle[  834] = 1'b1;  addr_rom[  834]='h00000d08;  wr_data_rom[  834]='h00000b57;
    rd_cycle[  835] = 1'b0;  wr_cycle[  835] = 1'b1;  addr_rom[  835]='h00000d0c;  wr_data_rom[  835]='h00002410;
    rd_cycle[  836] = 1'b0;  wr_cycle[  836] = 1'b1;  addr_rom[  836]='h00000d10;  wr_data_rom[  836]='h00003de8;
    rd_cycle[  837] = 1'b0;  wr_cycle[  837] = 1'b1;  addr_rom[  837]='h00000d14;  wr_data_rom[  837]='h000004cf;
    rd_cycle[  838] = 1'b0;  wr_cycle[  838] = 1'b1;  addr_rom[  838]='h00000d18;  wr_data_rom[  838]='h000027be;
    rd_cycle[  839] = 1'b0;  wr_cycle[  839] = 1'b1;  addr_rom[  839]='h00000d1c;  wr_data_rom[  839]='h00000515;
    rd_cycle[  840] = 1'b0;  wr_cycle[  840] = 1'b1;  addr_rom[  840]='h00000d20;  wr_data_rom[  840]='h00002f77;
    rd_cycle[  841] = 1'b0;  wr_cycle[  841] = 1'b1;  addr_rom[  841]='h00000d24;  wr_data_rom[  841]='h00003f9f;
    rd_cycle[  842] = 1'b0;  wr_cycle[  842] = 1'b1;  addr_rom[  842]='h00000d28;  wr_data_rom[  842]='h00000d6d;
    rd_cycle[  843] = 1'b0;  wr_cycle[  843] = 1'b1;  addr_rom[  843]='h00000d2c;  wr_data_rom[  843]='h0000174e;
    rd_cycle[  844] = 1'b0;  wr_cycle[  844] = 1'b1;  addr_rom[  844]='h00000d30;  wr_data_rom[  844]='h000003e9;
    rd_cycle[  845] = 1'b0;  wr_cycle[  845] = 1'b1;  addr_rom[  845]='h00000d34;  wr_data_rom[  845]='h000015c8;
    rd_cycle[  846] = 1'b0;  wr_cycle[  846] = 1'b1;  addr_rom[  846]='h00000d38;  wr_data_rom[  846]='h00000baa;
    rd_cycle[  847] = 1'b0;  wr_cycle[  847] = 1'b1;  addr_rom[  847]='h00000d3c;  wr_data_rom[  847]='h00002c22;
    rd_cycle[  848] = 1'b0;  wr_cycle[  848] = 1'b1;  addr_rom[  848]='h00000d40;  wr_data_rom[  848]='h0000389a;
    rd_cycle[  849] = 1'b0;  wr_cycle[  849] = 1'b1;  addr_rom[  849]='h00000d44;  wr_data_rom[  849]='h000030e3;
    rd_cycle[  850] = 1'b0;  wr_cycle[  850] = 1'b1;  addr_rom[  850]='h00000d48;  wr_data_rom[  850]='h00002909;
    rd_cycle[  851] = 1'b0;  wr_cycle[  851] = 1'b1;  addr_rom[  851]='h00000d4c;  wr_data_rom[  851]='h00002e31;
    rd_cycle[  852] = 1'b0;  wr_cycle[  852] = 1'b1;  addr_rom[  852]='h00000d50;  wr_data_rom[  852]='h0000048a;
    rd_cycle[  853] = 1'b0;  wr_cycle[  853] = 1'b1;  addr_rom[  853]='h00000d54;  wr_data_rom[  853]='h000034f7;
    rd_cycle[  854] = 1'b0;  wr_cycle[  854] = 1'b1;  addr_rom[  854]='h00000d58;  wr_data_rom[  854]='h000020af;
    rd_cycle[  855] = 1'b0;  wr_cycle[  855] = 1'b1;  addr_rom[  855]='h00000d5c;  wr_data_rom[  855]='h000032e7;
    rd_cycle[  856] = 1'b0;  wr_cycle[  856] = 1'b1;  addr_rom[  856]='h00000d60;  wr_data_rom[  856]='h0000201e;
    rd_cycle[  857] = 1'b0;  wr_cycle[  857] = 1'b1;  addr_rom[  857]='h00000d64;  wr_data_rom[  857]='h0000169b;
    rd_cycle[  858] = 1'b0;  wr_cycle[  858] = 1'b1;  addr_rom[  858]='h00000d68;  wr_data_rom[  858]='h0000132c;
    rd_cycle[  859] = 1'b0;  wr_cycle[  859] = 1'b1;  addr_rom[  859]='h00000d6c;  wr_data_rom[  859]='h00002185;
    rd_cycle[  860] = 1'b0;  wr_cycle[  860] = 1'b1;  addr_rom[  860]='h00000d70;  wr_data_rom[  860]='h0000177f;
    rd_cycle[  861] = 1'b0;  wr_cycle[  861] = 1'b1;  addr_rom[  861]='h00000d74;  wr_data_rom[  861]='h00002bd5;
    rd_cycle[  862] = 1'b0;  wr_cycle[  862] = 1'b1;  addr_rom[  862]='h00000d78;  wr_data_rom[  862]='h00000159;
    rd_cycle[  863] = 1'b0;  wr_cycle[  863] = 1'b1;  addr_rom[  863]='h00000d7c;  wr_data_rom[  863]='h000034aa;
    rd_cycle[  864] = 1'b0;  wr_cycle[  864] = 1'b1;  addr_rom[  864]='h00000d80;  wr_data_rom[  864]='h00000b7c;
    rd_cycle[  865] = 1'b0;  wr_cycle[  865] = 1'b1;  addr_rom[  865]='h00000d84;  wr_data_rom[  865]='h000009d4;
    rd_cycle[  866] = 1'b0;  wr_cycle[  866] = 1'b1;  addr_rom[  866]='h00000d88;  wr_data_rom[  866]='h00002139;
    rd_cycle[  867] = 1'b0;  wr_cycle[  867] = 1'b1;  addr_rom[  867]='h00000d8c;  wr_data_rom[  867]='h00000d63;
    rd_cycle[  868] = 1'b0;  wr_cycle[  868] = 1'b1;  addr_rom[  868]='h00000d90;  wr_data_rom[  868]='h000012a7;
    rd_cycle[  869] = 1'b0;  wr_cycle[  869] = 1'b1;  addr_rom[  869]='h00000d94;  wr_data_rom[  869]='h00003014;
    rd_cycle[  870] = 1'b0;  wr_cycle[  870] = 1'b1;  addr_rom[  870]='h00000d98;  wr_data_rom[  870]='h00002b8f;
    rd_cycle[  871] = 1'b0;  wr_cycle[  871] = 1'b1;  addr_rom[  871]='h00000d9c;  wr_data_rom[  871]='h00003629;
    rd_cycle[  872] = 1'b0;  wr_cycle[  872] = 1'b1;  addr_rom[  872]='h00000da0;  wr_data_rom[  872]='h000026ec;
    rd_cycle[  873] = 1'b0;  wr_cycle[  873] = 1'b1;  addr_rom[  873]='h00000da4;  wr_data_rom[  873]='h0000065c;
    rd_cycle[  874] = 1'b0;  wr_cycle[  874] = 1'b1;  addr_rom[  874]='h00000da8;  wr_data_rom[  874]='h00003d5e;
    rd_cycle[  875] = 1'b0;  wr_cycle[  875] = 1'b1;  addr_rom[  875]='h00000dac;  wr_data_rom[  875]='h00002d95;
    rd_cycle[  876] = 1'b0;  wr_cycle[  876] = 1'b1;  addr_rom[  876]='h00000db0;  wr_data_rom[  876]='h000020e6;
    rd_cycle[  877] = 1'b0;  wr_cycle[  877] = 1'b1;  addr_rom[  877]='h00000db4;  wr_data_rom[  877]='h000003e3;
    rd_cycle[  878] = 1'b0;  wr_cycle[  878] = 1'b1;  addr_rom[  878]='h00000db8;  wr_data_rom[  878]='h00003e5d;
    rd_cycle[  879] = 1'b0;  wr_cycle[  879] = 1'b1;  addr_rom[  879]='h00000dbc;  wr_data_rom[  879]='h000033a2;
    rd_cycle[  880] = 1'b0;  wr_cycle[  880] = 1'b1;  addr_rom[  880]='h00000dc0;  wr_data_rom[  880]='h0000179d;
    rd_cycle[  881] = 1'b0;  wr_cycle[  881] = 1'b1;  addr_rom[  881]='h00000dc4;  wr_data_rom[  881]='h000001b4;
    rd_cycle[  882] = 1'b0;  wr_cycle[  882] = 1'b1;  addr_rom[  882]='h00000dc8;  wr_data_rom[  882]='h00000703;
    rd_cycle[  883] = 1'b0;  wr_cycle[  883] = 1'b1;  addr_rom[  883]='h00000dcc;  wr_data_rom[  883]='h000029c9;
    rd_cycle[  884] = 1'b0;  wr_cycle[  884] = 1'b1;  addr_rom[  884]='h00000dd0;  wr_data_rom[  884]='h0000323d;
    rd_cycle[  885] = 1'b0;  wr_cycle[  885] = 1'b1;  addr_rom[  885]='h00000dd4;  wr_data_rom[  885]='h00001c1e;
    rd_cycle[  886] = 1'b0;  wr_cycle[  886] = 1'b1;  addr_rom[  886]='h00000dd8;  wr_data_rom[  886]='h00003d9c;
    rd_cycle[  887] = 1'b0;  wr_cycle[  887] = 1'b1;  addr_rom[  887]='h00000ddc;  wr_data_rom[  887]='h0000070e;
    rd_cycle[  888] = 1'b0;  wr_cycle[  888] = 1'b1;  addr_rom[  888]='h00000de0;  wr_data_rom[  888]='h0000332f;
    rd_cycle[  889] = 1'b0;  wr_cycle[  889] = 1'b1;  addr_rom[  889]='h00000de4;  wr_data_rom[  889]='h000038ca;
    rd_cycle[  890] = 1'b0;  wr_cycle[  890] = 1'b1;  addr_rom[  890]='h00000de8;  wr_data_rom[  890]='h000036e0;
    rd_cycle[  891] = 1'b0;  wr_cycle[  891] = 1'b1;  addr_rom[  891]='h00000dec;  wr_data_rom[  891]='h00000593;
    rd_cycle[  892] = 1'b0;  wr_cycle[  892] = 1'b1;  addr_rom[  892]='h00000df0;  wr_data_rom[  892]='h000004a0;
    rd_cycle[  893] = 1'b0;  wr_cycle[  893] = 1'b1;  addr_rom[  893]='h00000df4;  wr_data_rom[  893]='h00003cc0;
    rd_cycle[  894] = 1'b0;  wr_cycle[  894] = 1'b1;  addr_rom[  894]='h00000df8;  wr_data_rom[  894]='h00001e4e;
    rd_cycle[  895] = 1'b0;  wr_cycle[  895] = 1'b1;  addr_rom[  895]='h00000dfc;  wr_data_rom[  895]='h00000734;
    rd_cycle[  896] = 1'b0;  wr_cycle[  896] = 1'b1;  addr_rom[  896]='h00000e00;  wr_data_rom[  896]='h00003733;
    rd_cycle[  897] = 1'b0;  wr_cycle[  897] = 1'b1;  addr_rom[  897]='h00000e04;  wr_data_rom[  897]='h000009a6;
    rd_cycle[  898] = 1'b0;  wr_cycle[  898] = 1'b1;  addr_rom[  898]='h00000e08;  wr_data_rom[  898]='h000015c9;
    rd_cycle[  899] = 1'b0;  wr_cycle[  899] = 1'b1;  addr_rom[  899]='h00000e0c;  wr_data_rom[  899]='h00002c5f;
    rd_cycle[  900] = 1'b0;  wr_cycle[  900] = 1'b1;  addr_rom[  900]='h00000e10;  wr_data_rom[  900]='h00003954;
    rd_cycle[  901] = 1'b0;  wr_cycle[  901] = 1'b1;  addr_rom[  901]='h00000e14;  wr_data_rom[  901]='h000003f4;
    rd_cycle[  902] = 1'b0;  wr_cycle[  902] = 1'b1;  addr_rom[  902]='h00000e18;  wr_data_rom[  902]='h00002ea8;
    rd_cycle[  903] = 1'b0;  wr_cycle[  903] = 1'b1;  addr_rom[  903]='h00000e1c;  wr_data_rom[  903]='h00003636;
    rd_cycle[  904] = 1'b0;  wr_cycle[  904] = 1'b1;  addr_rom[  904]='h00000e20;  wr_data_rom[  904]='h00003d94;
    rd_cycle[  905] = 1'b0;  wr_cycle[  905] = 1'b1;  addr_rom[  905]='h00000e24;  wr_data_rom[  905]='h00002bc7;
    rd_cycle[  906] = 1'b0;  wr_cycle[  906] = 1'b1;  addr_rom[  906]='h00000e28;  wr_data_rom[  906]='h000014b1;
    rd_cycle[  907] = 1'b0;  wr_cycle[  907] = 1'b1;  addr_rom[  907]='h00000e2c;  wr_data_rom[  907]='h000013db;
    rd_cycle[  908] = 1'b0;  wr_cycle[  908] = 1'b1;  addr_rom[  908]='h00000e30;  wr_data_rom[  908]='h00003c27;
    rd_cycle[  909] = 1'b0;  wr_cycle[  909] = 1'b1;  addr_rom[  909]='h00000e34;  wr_data_rom[  909]='h0000158f;
    rd_cycle[  910] = 1'b0;  wr_cycle[  910] = 1'b1;  addr_rom[  910]='h00000e38;  wr_data_rom[  910]='h00000a06;
    rd_cycle[  911] = 1'b0;  wr_cycle[  911] = 1'b1;  addr_rom[  911]='h00000e3c;  wr_data_rom[  911]='h000031f4;
    rd_cycle[  912] = 1'b0;  wr_cycle[  912] = 1'b1;  addr_rom[  912]='h00000e40;  wr_data_rom[  912]='h00001d0a;
    rd_cycle[  913] = 1'b0;  wr_cycle[  913] = 1'b1;  addr_rom[  913]='h00000e44;  wr_data_rom[  913]='h00001fa1;
    rd_cycle[  914] = 1'b0;  wr_cycle[  914] = 1'b1;  addr_rom[  914]='h00000e48;  wr_data_rom[  914]='h00003dc6;
    rd_cycle[  915] = 1'b0;  wr_cycle[  915] = 1'b1;  addr_rom[  915]='h00000e4c;  wr_data_rom[  915]='h00000218;
    rd_cycle[  916] = 1'b0;  wr_cycle[  916] = 1'b1;  addr_rom[  916]='h00000e50;  wr_data_rom[  916]='h000021b2;
    rd_cycle[  917] = 1'b0;  wr_cycle[  917] = 1'b1;  addr_rom[  917]='h00000e54;  wr_data_rom[  917]='h0000146c;
    rd_cycle[  918] = 1'b0;  wr_cycle[  918] = 1'b1;  addr_rom[  918]='h00000e58;  wr_data_rom[  918]='h000016a6;
    rd_cycle[  919] = 1'b0;  wr_cycle[  919] = 1'b1;  addr_rom[  919]='h00000e5c;  wr_data_rom[  919]='h00002a81;
    rd_cycle[  920] = 1'b0;  wr_cycle[  920] = 1'b1;  addr_rom[  920]='h00000e60;  wr_data_rom[  920]='h00001d20;
    rd_cycle[  921] = 1'b0;  wr_cycle[  921] = 1'b1;  addr_rom[  921]='h00000e64;  wr_data_rom[  921]='h000033ac;
    rd_cycle[  922] = 1'b0;  wr_cycle[  922] = 1'b1;  addr_rom[  922]='h00000e68;  wr_data_rom[  922]='h000031a7;
    rd_cycle[  923] = 1'b0;  wr_cycle[  923] = 1'b1;  addr_rom[  923]='h00000e6c;  wr_data_rom[  923]='h00001840;
    rd_cycle[  924] = 1'b0;  wr_cycle[  924] = 1'b1;  addr_rom[  924]='h00000e70;  wr_data_rom[  924]='h00000312;
    rd_cycle[  925] = 1'b0;  wr_cycle[  925] = 1'b1;  addr_rom[  925]='h00000e74;  wr_data_rom[  925]='h00001f6f;
    rd_cycle[  926] = 1'b0;  wr_cycle[  926] = 1'b1;  addr_rom[  926]='h00000e78;  wr_data_rom[  926]='h000028c2;
    rd_cycle[  927] = 1'b0;  wr_cycle[  927] = 1'b1;  addr_rom[  927]='h00000e7c;  wr_data_rom[  927]='h00001d5a;
    rd_cycle[  928] = 1'b0;  wr_cycle[  928] = 1'b1;  addr_rom[  928]='h00000e80;  wr_data_rom[  928]='h00003948;
    rd_cycle[  929] = 1'b0;  wr_cycle[  929] = 1'b1;  addr_rom[  929]='h00000e84;  wr_data_rom[  929]='h000002d3;
    rd_cycle[  930] = 1'b0;  wr_cycle[  930] = 1'b1;  addr_rom[  930]='h00000e88;  wr_data_rom[  930]='h00000cd1;
    rd_cycle[  931] = 1'b0;  wr_cycle[  931] = 1'b1;  addr_rom[  931]='h00000e8c;  wr_data_rom[  931]='h00000183;
    rd_cycle[  932] = 1'b0;  wr_cycle[  932] = 1'b1;  addr_rom[  932]='h00000e90;  wr_data_rom[  932]='h00002f37;
    rd_cycle[  933] = 1'b0;  wr_cycle[  933] = 1'b1;  addr_rom[  933]='h00000e94;  wr_data_rom[  933]='h00001024;
    rd_cycle[  934] = 1'b0;  wr_cycle[  934] = 1'b1;  addr_rom[  934]='h00000e98;  wr_data_rom[  934]='h00002132;
    rd_cycle[  935] = 1'b0;  wr_cycle[  935] = 1'b1;  addr_rom[  935]='h00000e9c;  wr_data_rom[  935]='h000035fa;
    rd_cycle[  936] = 1'b0;  wr_cycle[  936] = 1'b1;  addr_rom[  936]='h00000ea0;  wr_data_rom[  936]='h0000158d;
    rd_cycle[  937] = 1'b0;  wr_cycle[  937] = 1'b1;  addr_rom[  937]='h00000ea4;  wr_data_rom[  937]='h0000244e;
    rd_cycle[  938] = 1'b0;  wr_cycle[  938] = 1'b1;  addr_rom[  938]='h00000ea8;  wr_data_rom[  938]='h00003796;
    rd_cycle[  939] = 1'b0;  wr_cycle[  939] = 1'b1;  addr_rom[  939]='h00000eac;  wr_data_rom[  939]='h0000354e;
    rd_cycle[  940] = 1'b0;  wr_cycle[  940] = 1'b1;  addr_rom[  940]='h00000eb0;  wr_data_rom[  940]='h00002aed;
    rd_cycle[  941] = 1'b0;  wr_cycle[  941] = 1'b1;  addr_rom[  941]='h00000eb4;  wr_data_rom[  941]='h000010ec;
    rd_cycle[  942] = 1'b0;  wr_cycle[  942] = 1'b1;  addr_rom[  942]='h00000eb8;  wr_data_rom[  942]='h00000544;
    rd_cycle[  943] = 1'b0;  wr_cycle[  943] = 1'b1;  addr_rom[  943]='h00000ebc;  wr_data_rom[  943]='h000004c9;
    rd_cycle[  944] = 1'b0;  wr_cycle[  944] = 1'b1;  addr_rom[  944]='h00000ec0;  wr_data_rom[  944]='h00001cb6;
    rd_cycle[  945] = 1'b0;  wr_cycle[  945] = 1'b1;  addr_rom[  945]='h00000ec4;  wr_data_rom[  945]='h00000f13;
    rd_cycle[  946] = 1'b0;  wr_cycle[  946] = 1'b1;  addr_rom[  946]='h00000ec8;  wr_data_rom[  946]='h00000670;
    rd_cycle[  947] = 1'b0;  wr_cycle[  947] = 1'b1;  addr_rom[  947]='h00000ecc;  wr_data_rom[  947]='h0000091c;
    rd_cycle[  948] = 1'b0;  wr_cycle[  948] = 1'b1;  addr_rom[  948]='h00000ed0;  wr_data_rom[  948]='h000015ad;
    rd_cycle[  949] = 1'b0;  wr_cycle[  949] = 1'b1;  addr_rom[  949]='h00000ed4;  wr_data_rom[  949]='h00001a95;
    rd_cycle[  950] = 1'b0;  wr_cycle[  950] = 1'b1;  addr_rom[  950]='h00000ed8;  wr_data_rom[  950]='h00000700;
    rd_cycle[  951] = 1'b0;  wr_cycle[  951] = 1'b1;  addr_rom[  951]='h00000edc;  wr_data_rom[  951]='h00001116;
    rd_cycle[  952] = 1'b0;  wr_cycle[  952] = 1'b1;  addr_rom[  952]='h00000ee0;  wr_data_rom[  952]='h00001dad;
    rd_cycle[  953] = 1'b0;  wr_cycle[  953] = 1'b1;  addr_rom[  953]='h00000ee4;  wr_data_rom[  953]='h000036d5;
    rd_cycle[  954] = 1'b0;  wr_cycle[  954] = 1'b1;  addr_rom[  954]='h00000ee8;  wr_data_rom[  954]='h00002b0f;
    rd_cycle[  955] = 1'b0;  wr_cycle[  955] = 1'b1;  addr_rom[  955]='h00000eec;  wr_data_rom[  955]='h00002e39;
    rd_cycle[  956] = 1'b0;  wr_cycle[  956] = 1'b1;  addr_rom[  956]='h00000ef0;  wr_data_rom[  956]='h00001be2;
    rd_cycle[  957] = 1'b0;  wr_cycle[  957] = 1'b1;  addr_rom[  957]='h00000ef4;  wr_data_rom[  957]='h0000337f;
    rd_cycle[  958] = 1'b0;  wr_cycle[  958] = 1'b1;  addr_rom[  958]='h00000ef8;  wr_data_rom[  958]='h00001a93;
    rd_cycle[  959] = 1'b0;  wr_cycle[  959] = 1'b1;  addr_rom[  959]='h00000efc;  wr_data_rom[  959]='h00001f50;
    rd_cycle[  960] = 1'b0;  wr_cycle[  960] = 1'b1;  addr_rom[  960]='h00000f00;  wr_data_rom[  960]='h00003df7;
    rd_cycle[  961] = 1'b0;  wr_cycle[  961] = 1'b1;  addr_rom[  961]='h00000f04;  wr_data_rom[  961]='h00002fbc;
    rd_cycle[  962] = 1'b0;  wr_cycle[  962] = 1'b1;  addr_rom[  962]='h00000f08;  wr_data_rom[  962]='h00002326;
    rd_cycle[  963] = 1'b0;  wr_cycle[  963] = 1'b1;  addr_rom[  963]='h00000f0c;  wr_data_rom[  963]='h00002a0a;
    rd_cycle[  964] = 1'b0;  wr_cycle[  964] = 1'b1;  addr_rom[  964]='h00000f10;  wr_data_rom[  964]='h00002483;
    rd_cycle[  965] = 1'b0;  wr_cycle[  965] = 1'b1;  addr_rom[  965]='h00000f14;  wr_data_rom[  965]='h000018d9;
    rd_cycle[  966] = 1'b0;  wr_cycle[  966] = 1'b1;  addr_rom[  966]='h00000f18;  wr_data_rom[  966]='h00000b31;
    rd_cycle[  967] = 1'b0;  wr_cycle[  967] = 1'b1;  addr_rom[  967]='h00000f1c;  wr_data_rom[  967]='h00003f9f;
    rd_cycle[  968] = 1'b0;  wr_cycle[  968] = 1'b1;  addr_rom[  968]='h00000f20;  wr_data_rom[  968]='h0000028d;
    rd_cycle[  969] = 1'b0;  wr_cycle[  969] = 1'b1;  addr_rom[  969]='h00000f24;  wr_data_rom[  969]='h00003a1c;
    rd_cycle[  970] = 1'b0;  wr_cycle[  970] = 1'b1;  addr_rom[  970]='h00000f28;  wr_data_rom[  970]='h00003c66;
    rd_cycle[  971] = 1'b0;  wr_cycle[  971] = 1'b1;  addr_rom[  971]='h00000f2c;  wr_data_rom[  971]='h00001149;
    rd_cycle[  972] = 1'b0;  wr_cycle[  972] = 1'b1;  addr_rom[  972]='h00000f30;  wr_data_rom[  972]='h00002b32;
    rd_cycle[  973] = 1'b0;  wr_cycle[  973] = 1'b1;  addr_rom[  973]='h00000f34;  wr_data_rom[  973]='h000010bd;
    rd_cycle[  974] = 1'b0;  wr_cycle[  974] = 1'b1;  addr_rom[  974]='h00000f38;  wr_data_rom[  974]='h00000c96;
    rd_cycle[  975] = 1'b0;  wr_cycle[  975] = 1'b1;  addr_rom[  975]='h00000f3c;  wr_data_rom[  975]='h000021d3;
    rd_cycle[  976] = 1'b0;  wr_cycle[  976] = 1'b1;  addr_rom[  976]='h00000f40;  wr_data_rom[  976]='h00003bbe;
    rd_cycle[  977] = 1'b0;  wr_cycle[  977] = 1'b1;  addr_rom[  977]='h00000f44;  wr_data_rom[  977]='h00002d2f;
    rd_cycle[  978] = 1'b0;  wr_cycle[  978] = 1'b1;  addr_rom[  978]='h00000f48;  wr_data_rom[  978]='h000008cd;
    rd_cycle[  979] = 1'b0;  wr_cycle[  979] = 1'b1;  addr_rom[  979]='h00000f4c;  wr_data_rom[  979]='h00002539;
    rd_cycle[  980] = 1'b0;  wr_cycle[  980] = 1'b1;  addr_rom[  980]='h00000f50;  wr_data_rom[  980]='h0000217c;
    rd_cycle[  981] = 1'b0;  wr_cycle[  981] = 1'b1;  addr_rom[  981]='h00000f54;  wr_data_rom[  981]='h000016d9;
    rd_cycle[  982] = 1'b0;  wr_cycle[  982] = 1'b1;  addr_rom[  982]='h00000f58;  wr_data_rom[  982]='h0000392b;
    rd_cycle[  983] = 1'b0;  wr_cycle[  983] = 1'b1;  addr_rom[  983]='h00000f5c;  wr_data_rom[  983]='h000020f2;
    rd_cycle[  984] = 1'b0;  wr_cycle[  984] = 1'b1;  addr_rom[  984]='h00000f60;  wr_data_rom[  984]='h00001260;
    rd_cycle[  985] = 1'b0;  wr_cycle[  985] = 1'b1;  addr_rom[  985]='h00000f64;  wr_data_rom[  985]='h00000b02;
    rd_cycle[  986] = 1'b0;  wr_cycle[  986] = 1'b1;  addr_rom[  986]='h00000f68;  wr_data_rom[  986]='h00001b1d;
    rd_cycle[  987] = 1'b0;  wr_cycle[  987] = 1'b1;  addr_rom[  987]='h00000f6c;  wr_data_rom[  987]='h0000262f;
    rd_cycle[  988] = 1'b0;  wr_cycle[  988] = 1'b1;  addr_rom[  988]='h00000f70;  wr_data_rom[  988]='h00000a13;
    rd_cycle[  989] = 1'b0;  wr_cycle[  989] = 1'b1;  addr_rom[  989]='h00000f74;  wr_data_rom[  989]='h000039f5;
    rd_cycle[  990] = 1'b0;  wr_cycle[  990] = 1'b1;  addr_rom[  990]='h00000f78;  wr_data_rom[  990]='h00003f8c;
    rd_cycle[  991] = 1'b0;  wr_cycle[  991] = 1'b1;  addr_rom[  991]='h00000f7c;  wr_data_rom[  991]='h00003a8f;
    rd_cycle[  992] = 1'b0;  wr_cycle[  992] = 1'b1;  addr_rom[  992]='h00000f80;  wr_data_rom[  992]='h00003320;
    rd_cycle[  993] = 1'b0;  wr_cycle[  993] = 1'b1;  addr_rom[  993]='h00000f84;  wr_data_rom[  993]='h000020bd;
    rd_cycle[  994] = 1'b0;  wr_cycle[  994] = 1'b1;  addr_rom[  994]='h00000f88;  wr_data_rom[  994]='h00001994;
    rd_cycle[  995] = 1'b0;  wr_cycle[  995] = 1'b1;  addr_rom[  995]='h00000f8c;  wr_data_rom[  995]='h000032b3;
    rd_cycle[  996] = 1'b0;  wr_cycle[  996] = 1'b1;  addr_rom[  996]='h00000f90;  wr_data_rom[  996]='h000013fb;
    rd_cycle[  997] = 1'b0;  wr_cycle[  997] = 1'b1;  addr_rom[  997]='h00000f94;  wr_data_rom[  997]='h000028cc;
    rd_cycle[  998] = 1'b0;  wr_cycle[  998] = 1'b1;  addr_rom[  998]='h00000f98;  wr_data_rom[  998]='h00000973;
    rd_cycle[  999] = 1'b0;  wr_cycle[  999] = 1'b1;  addr_rom[  999]='h00000f9c;  wr_data_rom[  999]='h00000e9a;
    rd_cycle[ 1000] = 1'b0;  wr_cycle[ 1000] = 1'b1;  addr_rom[ 1000]='h00000fa0;  wr_data_rom[ 1000]='h00001d17;
    rd_cycle[ 1001] = 1'b0;  wr_cycle[ 1001] = 1'b1;  addr_rom[ 1001]='h00000fa4;  wr_data_rom[ 1001]='h000030e3;
    rd_cycle[ 1002] = 1'b0;  wr_cycle[ 1002] = 1'b1;  addr_rom[ 1002]='h00000fa8;  wr_data_rom[ 1002]='h0000192b;
    rd_cycle[ 1003] = 1'b0;  wr_cycle[ 1003] = 1'b1;  addr_rom[ 1003]='h00000fac;  wr_data_rom[ 1003]='h00000bb8;
    rd_cycle[ 1004] = 1'b0;  wr_cycle[ 1004] = 1'b1;  addr_rom[ 1004]='h00000fb0;  wr_data_rom[ 1004]='h00000138;
    rd_cycle[ 1005] = 1'b0;  wr_cycle[ 1005] = 1'b1;  addr_rom[ 1005]='h00000fb4;  wr_data_rom[ 1005]='h000022e9;
    rd_cycle[ 1006] = 1'b0;  wr_cycle[ 1006] = 1'b1;  addr_rom[ 1006]='h00000fb8;  wr_data_rom[ 1006]='h00001cfa;
    rd_cycle[ 1007] = 1'b0;  wr_cycle[ 1007] = 1'b1;  addr_rom[ 1007]='h00000fbc;  wr_data_rom[ 1007]='h00001c40;
    rd_cycle[ 1008] = 1'b0;  wr_cycle[ 1008] = 1'b1;  addr_rom[ 1008]='h00000fc0;  wr_data_rom[ 1008]='h0000220c;
    rd_cycle[ 1009] = 1'b0;  wr_cycle[ 1009] = 1'b1;  addr_rom[ 1009]='h00000fc4;  wr_data_rom[ 1009]='h00003403;
    rd_cycle[ 1010] = 1'b0;  wr_cycle[ 1010] = 1'b1;  addr_rom[ 1010]='h00000fc8;  wr_data_rom[ 1010]='h000037aa;
    rd_cycle[ 1011] = 1'b0;  wr_cycle[ 1011] = 1'b1;  addr_rom[ 1011]='h00000fcc;  wr_data_rom[ 1011]='h0000151b;
    rd_cycle[ 1012] = 1'b0;  wr_cycle[ 1012] = 1'b1;  addr_rom[ 1012]='h00000fd0;  wr_data_rom[ 1012]='h00002391;
    rd_cycle[ 1013] = 1'b0;  wr_cycle[ 1013] = 1'b1;  addr_rom[ 1013]='h00000fd4;  wr_data_rom[ 1013]='h0000228e;
    rd_cycle[ 1014] = 1'b0;  wr_cycle[ 1014] = 1'b1;  addr_rom[ 1014]='h00000fd8;  wr_data_rom[ 1014]='h0000353b;
    rd_cycle[ 1015] = 1'b0;  wr_cycle[ 1015] = 1'b1;  addr_rom[ 1015]='h00000fdc;  wr_data_rom[ 1015]='h000007f3;
    rd_cycle[ 1016] = 1'b0;  wr_cycle[ 1016] = 1'b1;  addr_rom[ 1016]='h00000fe0;  wr_data_rom[ 1016]='h00000f41;
    rd_cycle[ 1017] = 1'b0;  wr_cycle[ 1017] = 1'b1;  addr_rom[ 1017]='h00000fe4;  wr_data_rom[ 1017]='h000011c3;
    rd_cycle[ 1018] = 1'b0;  wr_cycle[ 1018] = 1'b1;  addr_rom[ 1018]='h00000fe8;  wr_data_rom[ 1018]='h00001208;
    rd_cycle[ 1019] = 1'b0;  wr_cycle[ 1019] = 1'b1;  addr_rom[ 1019]='h00000fec;  wr_data_rom[ 1019]='h00000e00;
    rd_cycle[ 1020] = 1'b0;  wr_cycle[ 1020] = 1'b1;  addr_rom[ 1020]='h00000ff0;  wr_data_rom[ 1020]='h00001009;
    rd_cycle[ 1021] = 1'b0;  wr_cycle[ 1021] = 1'b1;  addr_rom[ 1021]='h00000ff4;  wr_data_rom[ 1021]='h00003382;
    rd_cycle[ 1022] = 1'b0;  wr_cycle[ 1022] = 1'b1;  addr_rom[ 1022]='h00000ff8;  wr_data_rom[ 1022]='h000030ec;
    rd_cycle[ 1023] = 1'b0;  wr_cycle[ 1023] = 1'b1;  addr_rom[ 1023]='h00000ffc;  wr_data_rom[ 1023]='h00002b40;
    rd_cycle[ 1024] = 1'b0;  wr_cycle[ 1024] = 1'b1;  addr_rom[ 1024]='h00001000;  wr_data_rom[ 1024]='h000011a6;
    rd_cycle[ 1025] = 1'b0;  wr_cycle[ 1025] = 1'b1;  addr_rom[ 1025]='h00001004;  wr_data_rom[ 1025]='h00001941;
    rd_cycle[ 1026] = 1'b0;  wr_cycle[ 1026] = 1'b1;  addr_rom[ 1026]='h00001008;  wr_data_rom[ 1026]='h00001f1d;
    rd_cycle[ 1027] = 1'b0;  wr_cycle[ 1027] = 1'b1;  addr_rom[ 1027]='h0000100c;  wr_data_rom[ 1027]='h00003261;
    rd_cycle[ 1028] = 1'b0;  wr_cycle[ 1028] = 1'b1;  addr_rom[ 1028]='h00001010;  wr_data_rom[ 1028]='h00001ed5;
    rd_cycle[ 1029] = 1'b0;  wr_cycle[ 1029] = 1'b1;  addr_rom[ 1029]='h00001014;  wr_data_rom[ 1029]='h00003412;
    rd_cycle[ 1030] = 1'b0;  wr_cycle[ 1030] = 1'b1;  addr_rom[ 1030]='h00001018;  wr_data_rom[ 1030]='h00001097;
    rd_cycle[ 1031] = 1'b0;  wr_cycle[ 1031] = 1'b1;  addr_rom[ 1031]='h0000101c;  wr_data_rom[ 1031]='h0000055f;
    rd_cycle[ 1032] = 1'b0;  wr_cycle[ 1032] = 1'b1;  addr_rom[ 1032]='h00001020;  wr_data_rom[ 1032]='h000029cf;
    rd_cycle[ 1033] = 1'b0;  wr_cycle[ 1033] = 1'b1;  addr_rom[ 1033]='h00001024;  wr_data_rom[ 1033]='h00000af0;
    rd_cycle[ 1034] = 1'b0;  wr_cycle[ 1034] = 1'b1;  addr_rom[ 1034]='h00001028;  wr_data_rom[ 1034]='h00000038;
    rd_cycle[ 1035] = 1'b0;  wr_cycle[ 1035] = 1'b1;  addr_rom[ 1035]='h0000102c;  wr_data_rom[ 1035]='h00000a39;
    rd_cycle[ 1036] = 1'b0;  wr_cycle[ 1036] = 1'b1;  addr_rom[ 1036]='h00001030;  wr_data_rom[ 1036]='h000000a5;
    rd_cycle[ 1037] = 1'b0;  wr_cycle[ 1037] = 1'b1;  addr_rom[ 1037]='h00001034;  wr_data_rom[ 1037]='h000003d9;
    rd_cycle[ 1038] = 1'b0;  wr_cycle[ 1038] = 1'b1;  addr_rom[ 1038]='h00001038;  wr_data_rom[ 1038]='h0000035c;
    rd_cycle[ 1039] = 1'b0;  wr_cycle[ 1039] = 1'b1;  addr_rom[ 1039]='h0000103c;  wr_data_rom[ 1039]='h00003f0b;
    rd_cycle[ 1040] = 1'b0;  wr_cycle[ 1040] = 1'b1;  addr_rom[ 1040]='h00001040;  wr_data_rom[ 1040]='h00002c9e;
    rd_cycle[ 1041] = 1'b0;  wr_cycle[ 1041] = 1'b1;  addr_rom[ 1041]='h00001044;  wr_data_rom[ 1041]='h00002e0a;
    rd_cycle[ 1042] = 1'b0;  wr_cycle[ 1042] = 1'b1;  addr_rom[ 1042]='h00001048;  wr_data_rom[ 1042]='h00000dcb;
    rd_cycle[ 1043] = 1'b0;  wr_cycle[ 1043] = 1'b1;  addr_rom[ 1043]='h0000104c;  wr_data_rom[ 1043]='h00003777;
    rd_cycle[ 1044] = 1'b0;  wr_cycle[ 1044] = 1'b1;  addr_rom[ 1044]='h00001050;  wr_data_rom[ 1044]='h00001f3c;
    rd_cycle[ 1045] = 1'b0;  wr_cycle[ 1045] = 1'b1;  addr_rom[ 1045]='h00001054;  wr_data_rom[ 1045]='h000003b9;
    rd_cycle[ 1046] = 1'b0;  wr_cycle[ 1046] = 1'b1;  addr_rom[ 1046]='h00001058;  wr_data_rom[ 1046]='h00002e5d;
    rd_cycle[ 1047] = 1'b0;  wr_cycle[ 1047] = 1'b1;  addr_rom[ 1047]='h0000105c;  wr_data_rom[ 1047]='h0000105d;
    rd_cycle[ 1048] = 1'b0;  wr_cycle[ 1048] = 1'b1;  addr_rom[ 1048]='h00001060;  wr_data_rom[ 1048]='h000011f8;
    rd_cycle[ 1049] = 1'b0;  wr_cycle[ 1049] = 1'b1;  addr_rom[ 1049]='h00001064;  wr_data_rom[ 1049]='h00000234;
    rd_cycle[ 1050] = 1'b0;  wr_cycle[ 1050] = 1'b1;  addr_rom[ 1050]='h00001068;  wr_data_rom[ 1050]='h000014bf;
    rd_cycle[ 1051] = 1'b0;  wr_cycle[ 1051] = 1'b1;  addr_rom[ 1051]='h0000106c;  wr_data_rom[ 1051]='h00000449;
    rd_cycle[ 1052] = 1'b0;  wr_cycle[ 1052] = 1'b1;  addr_rom[ 1052]='h00001070;  wr_data_rom[ 1052]='h00001856;
    rd_cycle[ 1053] = 1'b0;  wr_cycle[ 1053] = 1'b1;  addr_rom[ 1053]='h00001074;  wr_data_rom[ 1053]='h000030d6;
    rd_cycle[ 1054] = 1'b0;  wr_cycle[ 1054] = 1'b1;  addr_rom[ 1054]='h00001078;  wr_data_rom[ 1054]='h00000d5f;
    rd_cycle[ 1055] = 1'b0;  wr_cycle[ 1055] = 1'b1;  addr_rom[ 1055]='h0000107c;  wr_data_rom[ 1055]='h000019da;
    rd_cycle[ 1056] = 1'b0;  wr_cycle[ 1056] = 1'b1;  addr_rom[ 1056]='h00001080;  wr_data_rom[ 1056]='h00000c31;
    rd_cycle[ 1057] = 1'b0;  wr_cycle[ 1057] = 1'b1;  addr_rom[ 1057]='h00001084;  wr_data_rom[ 1057]='h00002617;
    rd_cycle[ 1058] = 1'b0;  wr_cycle[ 1058] = 1'b1;  addr_rom[ 1058]='h00001088;  wr_data_rom[ 1058]='h00001d17;
    rd_cycle[ 1059] = 1'b0;  wr_cycle[ 1059] = 1'b1;  addr_rom[ 1059]='h0000108c;  wr_data_rom[ 1059]='h00001b2a;
    rd_cycle[ 1060] = 1'b0;  wr_cycle[ 1060] = 1'b1;  addr_rom[ 1060]='h00001090;  wr_data_rom[ 1060]='h00000151;
    rd_cycle[ 1061] = 1'b0;  wr_cycle[ 1061] = 1'b1;  addr_rom[ 1061]='h00001094;  wr_data_rom[ 1061]='h0000295a;
    rd_cycle[ 1062] = 1'b0;  wr_cycle[ 1062] = 1'b1;  addr_rom[ 1062]='h00001098;  wr_data_rom[ 1062]='h0000348f;
    rd_cycle[ 1063] = 1'b0;  wr_cycle[ 1063] = 1'b1;  addr_rom[ 1063]='h0000109c;  wr_data_rom[ 1063]='h00003d06;
    rd_cycle[ 1064] = 1'b0;  wr_cycle[ 1064] = 1'b1;  addr_rom[ 1064]='h000010a0;  wr_data_rom[ 1064]='h00003bf4;
    rd_cycle[ 1065] = 1'b0;  wr_cycle[ 1065] = 1'b1;  addr_rom[ 1065]='h000010a4;  wr_data_rom[ 1065]='h00002d65;
    rd_cycle[ 1066] = 1'b0;  wr_cycle[ 1066] = 1'b1;  addr_rom[ 1066]='h000010a8;  wr_data_rom[ 1066]='h00003b35;
    rd_cycle[ 1067] = 1'b0;  wr_cycle[ 1067] = 1'b1;  addr_rom[ 1067]='h000010ac;  wr_data_rom[ 1067]='h00002dbd;
    rd_cycle[ 1068] = 1'b0;  wr_cycle[ 1068] = 1'b1;  addr_rom[ 1068]='h000010b0;  wr_data_rom[ 1068]='h0000057c;
    rd_cycle[ 1069] = 1'b0;  wr_cycle[ 1069] = 1'b1;  addr_rom[ 1069]='h000010b4;  wr_data_rom[ 1069]='h00001669;
    rd_cycle[ 1070] = 1'b0;  wr_cycle[ 1070] = 1'b1;  addr_rom[ 1070]='h000010b8;  wr_data_rom[ 1070]='h00003505;
    rd_cycle[ 1071] = 1'b0;  wr_cycle[ 1071] = 1'b1;  addr_rom[ 1071]='h000010bc;  wr_data_rom[ 1071]='h00001634;
    rd_cycle[ 1072] = 1'b0;  wr_cycle[ 1072] = 1'b1;  addr_rom[ 1072]='h000010c0;  wr_data_rom[ 1072]='h000038bb;
    rd_cycle[ 1073] = 1'b0;  wr_cycle[ 1073] = 1'b1;  addr_rom[ 1073]='h000010c4;  wr_data_rom[ 1073]='h00003a8e;
    rd_cycle[ 1074] = 1'b0;  wr_cycle[ 1074] = 1'b1;  addr_rom[ 1074]='h000010c8;  wr_data_rom[ 1074]='h000017a0;
    rd_cycle[ 1075] = 1'b0;  wr_cycle[ 1075] = 1'b1;  addr_rom[ 1075]='h000010cc;  wr_data_rom[ 1075]='h00002fc1;
    rd_cycle[ 1076] = 1'b0;  wr_cycle[ 1076] = 1'b1;  addr_rom[ 1076]='h000010d0;  wr_data_rom[ 1076]='h00002d5f;
    rd_cycle[ 1077] = 1'b0;  wr_cycle[ 1077] = 1'b1;  addr_rom[ 1077]='h000010d4;  wr_data_rom[ 1077]='h00001963;
    rd_cycle[ 1078] = 1'b0;  wr_cycle[ 1078] = 1'b1;  addr_rom[ 1078]='h000010d8;  wr_data_rom[ 1078]='h000021a5;
    rd_cycle[ 1079] = 1'b0;  wr_cycle[ 1079] = 1'b1;  addr_rom[ 1079]='h000010dc;  wr_data_rom[ 1079]='h000023e1;
    rd_cycle[ 1080] = 1'b0;  wr_cycle[ 1080] = 1'b1;  addr_rom[ 1080]='h000010e0;  wr_data_rom[ 1080]='h00001e05;
    rd_cycle[ 1081] = 1'b0;  wr_cycle[ 1081] = 1'b1;  addr_rom[ 1081]='h000010e4;  wr_data_rom[ 1081]='h00002150;
    rd_cycle[ 1082] = 1'b0;  wr_cycle[ 1082] = 1'b1;  addr_rom[ 1082]='h000010e8;  wr_data_rom[ 1082]='h00003151;
    rd_cycle[ 1083] = 1'b0;  wr_cycle[ 1083] = 1'b1;  addr_rom[ 1083]='h000010ec;  wr_data_rom[ 1083]='h00003f2d;
    rd_cycle[ 1084] = 1'b0;  wr_cycle[ 1084] = 1'b1;  addr_rom[ 1084]='h000010f0;  wr_data_rom[ 1084]='h000013b4;
    rd_cycle[ 1085] = 1'b0;  wr_cycle[ 1085] = 1'b1;  addr_rom[ 1085]='h000010f4;  wr_data_rom[ 1085]='h00003c3b;
    rd_cycle[ 1086] = 1'b0;  wr_cycle[ 1086] = 1'b1;  addr_rom[ 1086]='h000010f8;  wr_data_rom[ 1086]='h000022f7;
    rd_cycle[ 1087] = 1'b0;  wr_cycle[ 1087] = 1'b1;  addr_rom[ 1087]='h000010fc;  wr_data_rom[ 1087]='h0000268e;
    rd_cycle[ 1088] = 1'b0;  wr_cycle[ 1088] = 1'b1;  addr_rom[ 1088]='h00001100;  wr_data_rom[ 1088]='h000021f4;
    rd_cycle[ 1089] = 1'b0;  wr_cycle[ 1089] = 1'b1;  addr_rom[ 1089]='h00001104;  wr_data_rom[ 1089]='h00002480;
    rd_cycle[ 1090] = 1'b0;  wr_cycle[ 1090] = 1'b1;  addr_rom[ 1090]='h00001108;  wr_data_rom[ 1090]='h000009e3;
    rd_cycle[ 1091] = 1'b0;  wr_cycle[ 1091] = 1'b1;  addr_rom[ 1091]='h0000110c;  wr_data_rom[ 1091]='h000012de;
    rd_cycle[ 1092] = 1'b0;  wr_cycle[ 1092] = 1'b1;  addr_rom[ 1092]='h00001110;  wr_data_rom[ 1092]='h0000242b;
    rd_cycle[ 1093] = 1'b0;  wr_cycle[ 1093] = 1'b1;  addr_rom[ 1093]='h00001114;  wr_data_rom[ 1093]='h000007ed;
    rd_cycle[ 1094] = 1'b0;  wr_cycle[ 1094] = 1'b1;  addr_rom[ 1094]='h00001118;  wr_data_rom[ 1094]='h0000068f;
    rd_cycle[ 1095] = 1'b0;  wr_cycle[ 1095] = 1'b1;  addr_rom[ 1095]='h0000111c;  wr_data_rom[ 1095]='h00001658;
    rd_cycle[ 1096] = 1'b0;  wr_cycle[ 1096] = 1'b1;  addr_rom[ 1096]='h00001120;  wr_data_rom[ 1096]='h000017c5;
    rd_cycle[ 1097] = 1'b0;  wr_cycle[ 1097] = 1'b1;  addr_rom[ 1097]='h00001124;  wr_data_rom[ 1097]='h00000cec;
    rd_cycle[ 1098] = 1'b0;  wr_cycle[ 1098] = 1'b1;  addr_rom[ 1098]='h00001128;  wr_data_rom[ 1098]='h00001382;
    rd_cycle[ 1099] = 1'b0;  wr_cycle[ 1099] = 1'b1;  addr_rom[ 1099]='h0000112c;  wr_data_rom[ 1099]='h00000a79;
    rd_cycle[ 1100] = 1'b0;  wr_cycle[ 1100] = 1'b1;  addr_rom[ 1100]='h00001130;  wr_data_rom[ 1100]='h00002187;
    rd_cycle[ 1101] = 1'b0;  wr_cycle[ 1101] = 1'b1;  addr_rom[ 1101]='h00001134;  wr_data_rom[ 1101]='h00003f85;
    rd_cycle[ 1102] = 1'b0;  wr_cycle[ 1102] = 1'b1;  addr_rom[ 1102]='h00001138;  wr_data_rom[ 1102]='h00002fc2;
    rd_cycle[ 1103] = 1'b0;  wr_cycle[ 1103] = 1'b1;  addr_rom[ 1103]='h0000113c;  wr_data_rom[ 1103]='h00000d04;
    rd_cycle[ 1104] = 1'b0;  wr_cycle[ 1104] = 1'b1;  addr_rom[ 1104]='h00001140;  wr_data_rom[ 1104]='h00003b4b;
    rd_cycle[ 1105] = 1'b0;  wr_cycle[ 1105] = 1'b1;  addr_rom[ 1105]='h00001144;  wr_data_rom[ 1105]='h00002faa;
    rd_cycle[ 1106] = 1'b0;  wr_cycle[ 1106] = 1'b1;  addr_rom[ 1106]='h00001148;  wr_data_rom[ 1106]='h0000173c;
    rd_cycle[ 1107] = 1'b0;  wr_cycle[ 1107] = 1'b1;  addr_rom[ 1107]='h0000114c;  wr_data_rom[ 1107]='h00001d48;
    rd_cycle[ 1108] = 1'b0;  wr_cycle[ 1108] = 1'b1;  addr_rom[ 1108]='h00001150;  wr_data_rom[ 1108]='h000018fd;
    rd_cycle[ 1109] = 1'b0;  wr_cycle[ 1109] = 1'b1;  addr_rom[ 1109]='h00001154;  wr_data_rom[ 1109]='h00000f8c;
    rd_cycle[ 1110] = 1'b0;  wr_cycle[ 1110] = 1'b1;  addr_rom[ 1110]='h00001158;  wr_data_rom[ 1110]='h00002316;
    rd_cycle[ 1111] = 1'b0;  wr_cycle[ 1111] = 1'b1;  addr_rom[ 1111]='h0000115c;  wr_data_rom[ 1111]='h00000bdb;
    rd_cycle[ 1112] = 1'b0;  wr_cycle[ 1112] = 1'b1;  addr_rom[ 1112]='h00001160;  wr_data_rom[ 1112]='h000036e5;
    rd_cycle[ 1113] = 1'b0;  wr_cycle[ 1113] = 1'b1;  addr_rom[ 1113]='h00001164;  wr_data_rom[ 1113]='h0000311a;
    rd_cycle[ 1114] = 1'b0;  wr_cycle[ 1114] = 1'b1;  addr_rom[ 1114]='h00001168;  wr_data_rom[ 1114]='h0000258d;
    rd_cycle[ 1115] = 1'b0;  wr_cycle[ 1115] = 1'b1;  addr_rom[ 1115]='h0000116c;  wr_data_rom[ 1115]='h00001609;
    rd_cycle[ 1116] = 1'b0;  wr_cycle[ 1116] = 1'b1;  addr_rom[ 1116]='h00001170;  wr_data_rom[ 1116]='h00001ef2;
    rd_cycle[ 1117] = 1'b0;  wr_cycle[ 1117] = 1'b1;  addr_rom[ 1117]='h00001174;  wr_data_rom[ 1117]='h00000fc7;
    rd_cycle[ 1118] = 1'b0;  wr_cycle[ 1118] = 1'b1;  addr_rom[ 1118]='h00001178;  wr_data_rom[ 1118]='h000012b9;
    rd_cycle[ 1119] = 1'b0;  wr_cycle[ 1119] = 1'b1;  addr_rom[ 1119]='h0000117c;  wr_data_rom[ 1119]='h00002097;
    rd_cycle[ 1120] = 1'b0;  wr_cycle[ 1120] = 1'b1;  addr_rom[ 1120]='h00001180;  wr_data_rom[ 1120]='h00003b4c;
    rd_cycle[ 1121] = 1'b0;  wr_cycle[ 1121] = 1'b1;  addr_rom[ 1121]='h00001184;  wr_data_rom[ 1121]='h00001244;
    rd_cycle[ 1122] = 1'b0;  wr_cycle[ 1122] = 1'b1;  addr_rom[ 1122]='h00001188;  wr_data_rom[ 1122]='h000033a9;
    rd_cycle[ 1123] = 1'b0;  wr_cycle[ 1123] = 1'b1;  addr_rom[ 1123]='h0000118c;  wr_data_rom[ 1123]='h00003cf3;
    rd_cycle[ 1124] = 1'b0;  wr_cycle[ 1124] = 1'b1;  addr_rom[ 1124]='h00001190;  wr_data_rom[ 1124]='h00003323;
    rd_cycle[ 1125] = 1'b0;  wr_cycle[ 1125] = 1'b1;  addr_rom[ 1125]='h00001194;  wr_data_rom[ 1125]='h0000073c;
    rd_cycle[ 1126] = 1'b0;  wr_cycle[ 1126] = 1'b1;  addr_rom[ 1126]='h00001198;  wr_data_rom[ 1126]='h00003994;
    rd_cycle[ 1127] = 1'b0;  wr_cycle[ 1127] = 1'b1;  addr_rom[ 1127]='h0000119c;  wr_data_rom[ 1127]='h00001c03;
    rd_cycle[ 1128] = 1'b0;  wr_cycle[ 1128] = 1'b1;  addr_rom[ 1128]='h000011a0;  wr_data_rom[ 1128]='h00001970;
    rd_cycle[ 1129] = 1'b0;  wr_cycle[ 1129] = 1'b1;  addr_rom[ 1129]='h000011a4;  wr_data_rom[ 1129]='h00003b80;
    rd_cycle[ 1130] = 1'b0;  wr_cycle[ 1130] = 1'b1;  addr_rom[ 1130]='h000011a8;  wr_data_rom[ 1130]='h000030ae;
    rd_cycle[ 1131] = 1'b0;  wr_cycle[ 1131] = 1'b1;  addr_rom[ 1131]='h000011ac;  wr_data_rom[ 1131]='h00000f7e;
    rd_cycle[ 1132] = 1'b0;  wr_cycle[ 1132] = 1'b1;  addr_rom[ 1132]='h000011b0;  wr_data_rom[ 1132]='h00002da0;
    rd_cycle[ 1133] = 1'b0;  wr_cycle[ 1133] = 1'b1;  addr_rom[ 1133]='h000011b4;  wr_data_rom[ 1133]='h0000106a;
    rd_cycle[ 1134] = 1'b0;  wr_cycle[ 1134] = 1'b1;  addr_rom[ 1134]='h000011b8;  wr_data_rom[ 1134]='h00002201;
    rd_cycle[ 1135] = 1'b0;  wr_cycle[ 1135] = 1'b1;  addr_rom[ 1135]='h000011bc;  wr_data_rom[ 1135]='h0000282d;
    rd_cycle[ 1136] = 1'b0;  wr_cycle[ 1136] = 1'b1;  addr_rom[ 1136]='h000011c0;  wr_data_rom[ 1136]='h00001da7;
    rd_cycle[ 1137] = 1'b0;  wr_cycle[ 1137] = 1'b1;  addr_rom[ 1137]='h000011c4;  wr_data_rom[ 1137]='h00000efd;
    rd_cycle[ 1138] = 1'b0;  wr_cycle[ 1138] = 1'b1;  addr_rom[ 1138]='h000011c8;  wr_data_rom[ 1138]='h0000208f;
    rd_cycle[ 1139] = 1'b0;  wr_cycle[ 1139] = 1'b1;  addr_rom[ 1139]='h000011cc;  wr_data_rom[ 1139]='h00003ab4;
    rd_cycle[ 1140] = 1'b0;  wr_cycle[ 1140] = 1'b1;  addr_rom[ 1140]='h000011d0;  wr_data_rom[ 1140]='h0000362b;
    rd_cycle[ 1141] = 1'b0;  wr_cycle[ 1141] = 1'b1;  addr_rom[ 1141]='h000011d4;  wr_data_rom[ 1141]='h00003f1d;
    rd_cycle[ 1142] = 1'b0;  wr_cycle[ 1142] = 1'b1;  addr_rom[ 1142]='h000011d8;  wr_data_rom[ 1142]='h000008d4;
    rd_cycle[ 1143] = 1'b0;  wr_cycle[ 1143] = 1'b1;  addr_rom[ 1143]='h000011dc;  wr_data_rom[ 1143]='h00000d67;
    rd_cycle[ 1144] = 1'b0;  wr_cycle[ 1144] = 1'b1;  addr_rom[ 1144]='h000011e0;  wr_data_rom[ 1144]='h0000065f;
    rd_cycle[ 1145] = 1'b0;  wr_cycle[ 1145] = 1'b1;  addr_rom[ 1145]='h000011e4;  wr_data_rom[ 1145]='h000024fe;
    rd_cycle[ 1146] = 1'b0;  wr_cycle[ 1146] = 1'b1;  addr_rom[ 1146]='h000011e8;  wr_data_rom[ 1146]='h00003041;
    rd_cycle[ 1147] = 1'b0;  wr_cycle[ 1147] = 1'b1;  addr_rom[ 1147]='h000011ec;  wr_data_rom[ 1147]='h000016ae;
    rd_cycle[ 1148] = 1'b0;  wr_cycle[ 1148] = 1'b1;  addr_rom[ 1148]='h000011f0;  wr_data_rom[ 1148]='h00000544;
    rd_cycle[ 1149] = 1'b0;  wr_cycle[ 1149] = 1'b1;  addr_rom[ 1149]='h000011f4;  wr_data_rom[ 1149]='h00003c12;
    rd_cycle[ 1150] = 1'b0;  wr_cycle[ 1150] = 1'b1;  addr_rom[ 1150]='h000011f8;  wr_data_rom[ 1150]='h00000be9;
    rd_cycle[ 1151] = 1'b0;  wr_cycle[ 1151] = 1'b1;  addr_rom[ 1151]='h000011fc;  wr_data_rom[ 1151]='h00003582;
    rd_cycle[ 1152] = 1'b0;  wr_cycle[ 1152] = 1'b1;  addr_rom[ 1152]='h00001200;  wr_data_rom[ 1152]='h00002f92;
    rd_cycle[ 1153] = 1'b0;  wr_cycle[ 1153] = 1'b1;  addr_rom[ 1153]='h00001204;  wr_data_rom[ 1153]='h00002eba;
    rd_cycle[ 1154] = 1'b0;  wr_cycle[ 1154] = 1'b1;  addr_rom[ 1154]='h00001208;  wr_data_rom[ 1154]='h00001337;
    rd_cycle[ 1155] = 1'b0;  wr_cycle[ 1155] = 1'b1;  addr_rom[ 1155]='h0000120c;  wr_data_rom[ 1155]='h0000165f;
    rd_cycle[ 1156] = 1'b0;  wr_cycle[ 1156] = 1'b1;  addr_rom[ 1156]='h00001210;  wr_data_rom[ 1156]='h00002537;
    rd_cycle[ 1157] = 1'b0;  wr_cycle[ 1157] = 1'b1;  addr_rom[ 1157]='h00001214;  wr_data_rom[ 1157]='h00001af0;
    rd_cycle[ 1158] = 1'b0;  wr_cycle[ 1158] = 1'b1;  addr_rom[ 1158]='h00001218;  wr_data_rom[ 1158]='h00003b4f;
    rd_cycle[ 1159] = 1'b0;  wr_cycle[ 1159] = 1'b1;  addr_rom[ 1159]='h0000121c;  wr_data_rom[ 1159]='h00000d10;
    rd_cycle[ 1160] = 1'b0;  wr_cycle[ 1160] = 1'b1;  addr_rom[ 1160]='h00001220;  wr_data_rom[ 1160]='h00003384;
    rd_cycle[ 1161] = 1'b0;  wr_cycle[ 1161] = 1'b1;  addr_rom[ 1161]='h00001224;  wr_data_rom[ 1161]='h0000331f;
    rd_cycle[ 1162] = 1'b0;  wr_cycle[ 1162] = 1'b1;  addr_rom[ 1162]='h00001228;  wr_data_rom[ 1162]='h00000298;
    rd_cycle[ 1163] = 1'b0;  wr_cycle[ 1163] = 1'b1;  addr_rom[ 1163]='h0000122c;  wr_data_rom[ 1163]='h000028a5;
    rd_cycle[ 1164] = 1'b0;  wr_cycle[ 1164] = 1'b1;  addr_rom[ 1164]='h00001230;  wr_data_rom[ 1164]='h00001eed;
    rd_cycle[ 1165] = 1'b0;  wr_cycle[ 1165] = 1'b1;  addr_rom[ 1165]='h00001234;  wr_data_rom[ 1165]='h00000673;
    rd_cycle[ 1166] = 1'b0;  wr_cycle[ 1166] = 1'b1;  addr_rom[ 1166]='h00001238;  wr_data_rom[ 1166]='h000030c9;
    rd_cycle[ 1167] = 1'b0;  wr_cycle[ 1167] = 1'b1;  addr_rom[ 1167]='h0000123c;  wr_data_rom[ 1167]='h00000b18;
    rd_cycle[ 1168] = 1'b0;  wr_cycle[ 1168] = 1'b1;  addr_rom[ 1168]='h00001240;  wr_data_rom[ 1168]='h000021d3;
    rd_cycle[ 1169] = 1'b0;  wr_cycle[ 1169] = 1'b1;  addr_rom[ 1169]='h00001244;  wr_data_rom[ 1169]='h00001cce;
    rd_cycle[ 1170] = 1'b0;  wr_cycle[ 1170] = 1'b1;  addr_rom[ 1170]='h00001248;  wr_data_rom[ 1170]='h00001255;
    rd_cycle[ 1171] = 1'b0;  wr_cycle[ 1171] = 1'b1;  addr_rom[ 1171]='h0000124c;  wr_data_rom[ 1171]='h00002e6a;
    rd_cycle[ 1172] = 1'b0;  wr_cycle[ 1172] = 1'b1;  addr_rom[ 1172]='h00001250;  wr_data_rom[ 1172]='h0000275f;
    rd_cycle[ 1173] = 1'b0;  wr_cycle[ 1173] = 1'b1;  addr_rom[ 1173]='h00001254;  wr_data_rom[ 1173]='h000016e1;
    rd_cycle[ 1174] = 1'b0;  wr_cycle[ 1174] = 1'b1;  addr_rom[ 1174]='h00001258;  wr_data_rom[ 1174]='h00002474;
    rd_cycle[ 1175] = 1'b0;  wr_cycle[ 1175] = 1'b1;  addr_rom[ 1175]='h0000125c;  wr_data_rom[ 1175]='h00000a83;
    rd_cycle[ 1176] = 1'b0;  wr_cycle[ 1176] = 1'b1;  addr_rom[ 1176]='h00001260;  wr_data_rom[ 1176]='h00002700;
    rd_cycle[ 1177] = 1'b0;  wr_cycle[ 1177] = 1'b1;  addr_rom[ 1177]='h00001264;  wr_data_rom[ 1177]='h00001fb2;
    rd_cycle[ 1178] = 1'b0;  wr_cycle[ 1178] = 1'b1;  addr_rom[ 1178]='h00001268;  wr_data_rom[ 1178]='h00000417;
    rd_cycle[ 1179] = 1'b0;  wr_cycle[ 1179] = 1'b1;  addr_rom[ 1179]='h0000126c;  wr_data_rom[ 1179]='h00003993;
    rd_cycle[ 1180] = 1'b0;  wr_cycle[ 1180] = 1'b1;  addr_rom[ 1180]='h00001270;  wr_data_rom[ 1180]='h00001534;
    rd_cycle[ 1181] = 1'b0;  wr_cycle[ 1181] = 1'b1;  addr_rom[ 1181]='h00001274;  wr_data_rom[ 1181]='h000021f6;
    rd_cycle[ 1182] = 1'b0;  wr_cycle[ 1182] = 1'b1;  addr_rom[ 1182]='h00001278;  wr_data_rom[ 1182]='h0000161e;
    rd_cycle[ 1183] = 1'b0;  wr_cycle[ 1183] = 1'b1;  addr_rom[ 1183]='h0000127c;  wr_data_rom[ 1183]='h00002a8c;
    rd_cycle[ 1184] = 1'b0;  wr_cycle[ 1184] = 1'b1;  addr_rom[ 1184]='h00001280;  wr_data_rom[ 1184]='h000016ea;
    rd_cycle[ 1185] = 1'b0;  wr_cycle[ 1185] = 1'b1;  addr_rom[ 1185]='h00001284;  wr_data_rom[ 1185]='h00001cde;
    rd_cycle[ 1186] = 1'b0;  wr_cycle[ 1186] = 1'b1;  addr_rom[ 1186]='h00001288;  wr_data_rom[ 1186]='h00002937;
    rd_cycle[ 1187] = 1'b0;  wr_cycle[ 1187] = 1'b1;  addr_rom[ 1187]='h0000128c;  wr_data_rom[ 1187]='h000020d5;
    rd_cycle[ 1188] = 1'b0;  wr_cycle[ 1188] = 1'b1;  addr_rom[ 1188]='h00001290;  wr_data_rom[ 1188]='h000029cf;
    rd_cycle[ 1189] = 1'b0;  wr_cycle[ 1189] = 1'b1;  addr_rom[ 1189]='h00001294;  wr_data_rom[ 1189]='h00001905;
    rd_cycle[ 1190] = 1'b0;  wr_cycle[ 1190] = 1'b1;  addr_rom[ 1190]='h00001298;  wr_data_rom[ 1190]='h00001a70;
    rd_cycle[ 1191] = 1'b0;  wr_cycle[ 1191] = 1'b1;  addr_rom[ 1191]='h0000129c;  wr_data_rom[ 1191]='h00002dfb;
    rd_cycle[ 1192] = 1'b0;  wr_cycle[ 1192] = 1'b1;  addr_rom[ 1192]='h000012a0;  wr_data_rom[ 1192]='h00003495;
    rd_cycle[ 1193] = 1'b0;  wr_cycle[ 1193] = 1'b1;  addr_rom[ 1193]='h000012a4;  wr_data_rom[ 1193]='h00001650;
    rd_cycle[ 1194] = 1'b0;  wr_cycle[ 1194] = 1'b1;  addr_rom[ 1194]='h000012a8;  wr_data_rom[ 1194]='h00001f45;
    rd_cycle[ 1195] = 1'b0;  wr_cycle[ 1195] = 1'b1;  addr_rom[ 1195]='h000012ac;  wr_data_rom[ 1195]='h0000373d;
    rd_cycle[ 1196] = 1'b0;  wr_cycle[ 1196] = 1'b1;  addr_rom[ 1196]='h000012b0;  wr_data_rom[ 1196]='h00002f73;
    rd_cycle[ 1197] = 1'b0;  wr_cycle[ 1197] = 1'b1;  addr_rom[ 1197]='h000012b4;  wr_data_rom[ 1197]='h000009c9;
    rd_cycle[ 1198] = 1'b0;  wr_cycle[ 1198] = 1'b1;  addr_rom[ 1198]='h000012b8;  wr_data_rom[ 1198]='h000002b8;
    rd_cycle[ 1199] = 1'b0;  wr_cycle[ 1199] = 1'b1;  addr_rom[ 1199]='h000012bc;  wr_data_rom[ 1199]='h00000f7f;
    rd_cycle[ 1200] = 1'b0;  wr_cycle[ 1200] = 1'b1;  addr_rom[ 1200]='h000012c0;  wr_data_rom[ 1200]='h0000053d;
    rd_cycle[ 1201] = 1'b0;  wr_cycle[ 1201] = 1'b1;  addr_rom[ 1201]='h000012c4;  wr_data_rom[ 1201]='h00001a42;
    rd_cycle[ 1202] = 1'b0;  wr_cycle[ 1202] = 1'b1;  addr_rom[ 1202]='h000012c8;  wr_data_rom[ 1202]='h0000098e;
    rd_cycle[ 1203] = 1'b0;  wr_cycle[ 1203] = 1'b1;  addr_rom[ 1203]='h000012cc;  wr_data_rom[ 1203]='h00003d36;
    rd_cycle[ 1204] = 1'b0;  wr_cycle[ 1204] = 1'b1;  addr_rom[ 1204]='h000012d0;  wr_data_rom[ 1204]='h0000023d;
    rd_cycle[ 1205] = 1'b0;  wr_cycle[ 1205] = 1'b1;  addr_rom[ 1205]='h000012d4;  wr_data_rom[ 1205]='h00000ef8;
    rd_cycle[ 1206] = 1'b0;  wr_cycle[ 1206] = 1'b1;  addr_rom[ 1206]='h000012d8;  wr_data_rom[ 1206]='h00000dd6;
    rd_cycle[ 1207] = 1'b0;  wr_cycle[ 1207] = 1'b1;  addr_rom[ 1207]='h000012dc;  wr_data_rom[ 1207]='h00002bb0;
    rd_cycle[ 1208] = 1'b0;  wr_cycle[ 1208] = 1'b1;  addr_rom[ 1208]='h000012e0;  wr_data_rom[ 1208]='h0000329d;
    rd_cycle[ 1209] = 1'b0;  wr_cycle[ 1209] = 1'b1;  addr_rom[ 1209]='h000012e4;  wr_data_rom[ 1209]='h0000191d;
    rd_cycle[ 1210] = 1'b0;  wr_cycle[ 1210] = 1'b1;  addr_rom[ 1210]='h000012e8;  wr_data_rom[ 1210]='h00003215;
    rd_cycle[ 1211] = 1'b0;  wr_cycle[ 1211] = 1'b1;  addr_rom[ 1211]='h000012ec;  wr_data_rom[ 1211]='h000006ae;
    rd_cycle[ 1212] = 1'b0;  wr_cycle[ 1212] = 1'b1;  addr_rom[ 1212]='h000012f0;  wr_data_rom[ 1212]='h0000117c;
    rd_cycle[ 1213] = 1'b0;  wr_cycle[ 1213] = 1'b1;  addr_rom[ 1213]='h000012f4;  wr_data_rom[ 1213]='h000008a3;
    rd_cycle[ 1214] = 1'b0;  wr_cycle[ 1214] = 1'b1;  addr_rom[ 1214]='h000012f8;  wr_data_rom[ 1214]='h00001541;
    rd_cycle[ 1215] = 1'b0;  wr_cycle[ 1215] = 1'b1;  addr_rom[ 1215]='h000012fc;  wr_data_rom[ 1215]='h000035fa;
    rd_cycle[ 1216] = 1'b0;  wr_cycle[ 1216] = 1'b1;  addr_rom[ 1216]='h00001300;  wr_data_rom[ 1216]='h00000368;
    rd_cycle[ 1217] = 1'b0;  wr_cycle[ 1217] = 1'b1;  addr_rom[ 1217]='h00001304;  wr_data_rom[ 1217]='h0000138b;
    rd_cycle[ 1218] = 1'b0;  wr_cycle[ 1218] = 1'b1;  addr_rom[ 1218]='h00001308;  wr_data_rom[ 1218]='h00001314;
    rd_cycle[ 1219] = 1'b0;  wr_cycle[ 1219] = 1'b1;  addr_rom[ 1219]='h0000130c;  wr_data_rom[ 1219]='h0000151a;
    rd_cycle[ 1220] = 1'b0;  wr_cycle[ 1220] = 1'b1;  addr_rom[ 1220]='h00001310;  wr_data_rom[ 1220]='h00000dc7;
    rd_cycle[ 1221] = 1'b0;  wr_cycle[ 1221] = 1'b1;  addr_rom[ 1221]='h00001314;  wr_data_rom[ 1221]='h00000227;
    rd_cycle[ 1222] = 1'b0;  wr_cycle[ 1222] = 1'b1;  addr_rom[ 1222]='h00001318;  wr_data_rom[ 1222]='h00001bf7;
    rd_cycle[ 1223] = 1'b0;  wr_cycle[ 1223] = 1'b1;  addr_rom[ 1223]='h0000131c;  wr_data_rom[ 1223]='h00003c9d;
    rd_cycle[ 1224] = 1'b0;  wr_cycle[ 1224] = 1'b1;  addr_rom[ 1224]='h00001320;  wr_data_rom[ 1224]='h00001e5a;
    rd_cycle[ 1225] = 1'b0;  wr_cycle[ 1225] = 1'b1;  addr_rom[ 1225]='h00001324;  wr_data_rom[ 1225]='h000022b9;
    rd_cycle[ 1226] = 1'b0;  wr_cycle[ 1226] = 1'b1;  addr_rom[ 1226]='h00001328;  wr_data_rom[ 1226]='h00000f7f;
    rd_cycle[ 1227] = 1'b0;  wr_cycle[ 1227] = 1'b1;  addr_rom[ 1227]='h0000132c;  wr_data_rom[ 1227]='h00002665;
    rd_cycle[ 1228] = 1'b0;  wr_cycle[ 1228] = 1'b1;  addr_rom[ 1228]='h00001330;  wr_data_rom[ 1228]='h0000115d;
    rd_cycle[ 1229] = 1'b0;  wr_cycle[ 1229] = 1'b1;  addr_rom[ 1229]='h00001334;  wr_data_rom[ 1229]='h00002536;
    rd_cycle[ 1230] = 1'b0;  wr_cycle[ 1230] = 1'b1;  addr_rom[ 1230]='h00001338;  wr_data_rom[ 1230]='h00003f76;
    rd_cycle[ 1231] = 1'b0;  wr_cycle[ 1231] = 1'b1;  addr_rom[ 1231]='h0000133c;  wr_data_rom[ 1231]='h00000250;
    rd_cycle[ 1232] = 1'b0;  wr_cycle[ 1232] = 1'b1;  addr_rom[ 1232]='h00001340;  wr_data_rom[ 1232]='h000008c0;
    rd_cycle[ 1233] = 1'b0;  wr_cycle[ 1233] = 1'b1;  addr_rom[ 1233]='h00001344;  wr_data_rom[ 1233]='h00003c6e;
    rd_cycle[ 1234] = 1'b0;  wr_cycle[ 1234] = 1'b1;  addr_rom[ 1234]='h00001348;  wr_data_rom[ 1234]='h00002c52;
    rd_cycle[ 1235] = 1'b0;  wr_cycle[ 1235] = 1'b1;  addr_rom[ 1235]='h0000134c;  wr_data_rom[ 1235]='h000031b7;
    rd_cycle[ 1236] = 1'b0;  wr_cycle[ 1236] = 1'b1;  addr_rom[ 1236]='h00001350;  wr_data_rom[ 1236]='h000035ee;
    rd_cycle[ 1237] = 1'b0;  wr_cycle[ 1237] = 1'b1;  addr_rom[ 1237]='h00001354;  wr_data_rom[ 1237]='h00003210;
    rd_cycle[ 1238] = 1'b0;  wr_cycle[ 1238] = 1'b1;  addr_rom[ 1238]='h00001358;  wr_data_rom[ 1238]='h000023db;
    rd_cycle[ 1239] = 1'b0;  wr_cycle[ 1239] = 1'b1;  addr_rom[ 1239]='h0000135c;  wr_data_rom[ 1239]='h00003e76;
    rd_cycle[ 1240] = 1'b0;  wr_cycle[ 1240] = 1'b1;  addr_rom[ 1240]='h00001360;  wr_data_rom[ 1240]='h000010ac;
    rd_cycle[ 1241] = 1'b0;  wr_cycle[ 1241] = 1'b1;  addr_rom[ 1241]='h00001364;  wr_data_rom[ 1241]='h00003066;
    rd_cycle[ 1242] = 1'b0;  wr_cycle[ 1242] = 1'b1;  addr_rom[ 1242]='h00001368;  wr_data_rom[ 1242]='h00001805;
    rd_cycle[ 1243] = 1'b0;  wr_cycle[ 1243] = 1'b1;  addr_rom[ 1243]='h0000136c;  wr_data_rom[ 1243]='h00000d8c;
    rd_cycle[ 1244] = 1'b0;  wr_cycle[ 1244] = 1'b1;  addr_rom[ 1244]='h00001370;  wr_data_rom[ 1244]='h00002a69;
    rd_cycle[ 1245] = 1'b0;  wr_cycle[ 1245] = 1'b1;  addr_rom[ 1245]='h00001374;  wr_data_rom[ 1245]='h000002b2;
    rd_cycle[ 1246] = 1'b0;  wr_cycle[ 1246] = 1'b1;  addr_rom[ 1246]='h00001378;  wr_data_rom[ 1246]='h00003758;
    rd_cycle[ 1247] = 1'b0;  wr_cycle[ 1247] = 1'b1;  addr_rom[ 1247]='h0000137c;  wr_data_rom[ 1247]='h00003620;
    rd_cycle[ 1248] = 1'b0;  wr_cycle[ 1248] = 1'b1;  addr_rom[ 1248]='h00001380;  wr_data_rom[ 1248]='h00001a33;
    rd_cycle[ 1249] = 1'b0;  wr_cycle[ 1249] = 1'b1;  addr_rom[ 1249]='h00001384;  wr_data_rom[ 1249]='h00001fe6;
    rd_cycle[ 1250] = 1'b0;  wr_cycle[ 1250] = 1'b1;  addr_rom[ 1250]='h00001388;  wr_data_rom[ 1250]='h00003695;
    rd_cycle[ 1251] = 1'b0;  wr_cycle[ 1251] = 1'b1;  addr_rom[ 1251]='h0000138c;  wr_data_rom[ 1251]='h00003eb3;
    rd_cycle[ 1252] = 1'b0;  wr_cycle[ 1252] = 1'b1;  addr_rom[ 1252]='h00001390;  wr_data_rom[ 1252]='h00000aa7;
    rd_cycle[ 1253] = 1'b0;  wr_cycle[ 1253] = 1'b1;  addr_rom[ 1253]='h00001394;  wr_data_rom[ 1253]='h00003901;
    rd_cycle[ 1254] = 1'b0;  wr_cycle[ 1254] = 1'b1;  addr_rom[ 1254]='h00001398;  wr_data_rom[ 1254]='h00002e6b;
    rd_cycle[ 1255] = 1'b0;  wr_cycle[ 1255] = 1'b1;  addr_rom[ 1255]='h0000139c;  wr_data_rom[ 1255]='h0000162b;
    rd_cycle[ 1256] = 1'b0;  wr_cycle[ 1256] = 1'b1;  addr_rom[ 1256]='h000013a0;  wr_data_rom[ 1256]='h00002367;
    rd_cycle[ 1257] = 1'b0;  wr_cycle[ 1257] = 1'b1;  addr_rom[ 1257]='h000013a4;  wr_data_rom[ 1257]='h00002f96;
    rd_cycle[ 1258] = 1'b0;  wr_cycle[ 1258] = 1'b1;  addr_rom[ 1258]='h000013a8;  wr_data_rom[ 1258]='h00001791;
    rd_cycle[ 1259] = 1'b0;  wr_cycle[ 1259] = 1'b1;  addr_rom[ 1259]='h000013ac;  wr_data_rom[ 1259]='h00003eb1;
    rd_cycle[ 1260] = 1'b0;  wr_cycle[ 1260] = 1'b1;  addr_rom[ 1260]='h000013b0;  wr_data_rom[ 1260]='h000029ee;
    rd_cycle[ 1261] = 1'b0;  wr_cycle[ 1261] = 1'b1;  addr_rom[ 1261]='h000013b4;  wr_data_rom[ 1261]='h00001427;
    rd_cycle[ 1262] = 1'b0;  wr_cycle[ 1262] = 1'b1;  addr_rom[ 1262]='h000013b8;  wr_data_rom[ 1262]='h000007cd;
    rd_cycle[ 1263] = 1'b0;  wr_cycle[ 1263] = 1'b1;  addr_rom[ 1263]='h000013bc;  wr_data_rom[ 1263]='h00002638;
    rd_cycle[ 1264] = 1'b0;  wr_cycle[ 1264] = 1'b1;  addr_rom[ 1264]='h000013c0;  wr_data_rom[ 1264]='h0000137b;
    rd_cycle[ 1265] = 1'b0;  wr_cycle[ 1265] = 1'b1;  addr_rom[ 1265]='h000013c4;  wr_data_rom[ 1265]='h00003d21;
    rd_cycle[ 1266] = 1'b0;  wr_cycle[ 1266] = 1'b1;  addr_rom[ 1266]='h000013c8;  wr_data_rom[ 1266]='h00000cf6;
    rd_cycle[ 1267] = 1'b0;  wr_cycle[ 1267] = 1'b1;  addr_rom[ 1267]='h000013cc;  wr_data_rom[ 1267]='h0000122d;
    rd_cycle[ 1268] = 1'b0;  wr_cycle[ 1268] = 1'b1;  addr_rom[ 1268]='h000013d0;  wr_data_rom[ 1268]='h00001f03;
    rd_cycle[ 1269] = 1'b0;  wr_cycle[ 1269] = 1'b1;  addr_rom[ 1269]='h000013d4;  wr_data_rom[ 1269]='h00003e4c;
    rd_cycle[ 1270] = 1'b0;  wr_cycle[ 1270] = 1'b1;  addr_rom[ 1270]='h000013d8;  wr_data_rom[ 1270]='h00000631;
    rd_cycle[ 1271] = 1'b0;  wr_cycle[ 1271] = 1'b1;  addr_rom[ 1271]='h000013dc;  wr_data_rom[ 1271]='h00000651;
    rd_cycle[ 1272] = 1'b0;  wr_cycle[ 1272] = 1'b1;  addr_rom[ 1272]='h000013e0;  wr_data_rom[ 1272]='h0000372c;
    rd_cycle[ 1273] = 1'b0;  wr_cycle[ 1273] = 1'b1;  addr_rom[ 1273]='h000013e4;  wr_data_rom[ 1273]='h000024e8;
    rd_cycle[ 1274] = 1'b0;  wr_cycle[ 1274] = 1'b1;  addr_rom[ 1274]='h000013e8;  wr_data_rom[ 1274]='h000013fc;
    rd_cycle[ 1275] = 1'b0;  wr_cycle[ 1275] = 1'b1;  addr_rom[ 1275]='h000013ec;  wr_data_rom[ 1275]='h00001ca0;
    rd_cycle[ 1276] = 1'b0;  wr_cycle[ 1276] = 1'b1;  addr_rom[ 1276]='h000013f0;  wr_data_rom[ 1276]='h000002ba;
    rd_cycle[ 1277] = 1'b0;  wr_cycle[ 1277] = 1'b1;  addr_rom[ 1277]='h000013f4;  wr_data_rom[ 1277]='h000009c4;
    rd_cycle[ 1278] = 1'b0;  wr_cycle[ 1278] = 1'b1;  addr_rom[ 1278]='h000013f8;  wr_data_rom[ 1278]='h0000331d;
    rd_cycle[ 1279] = 1'b0;  wr_cycle[ 1279] = 1'b1;  addr_rom[ 1279]='h000013fc;  wr_data_rom[ 1279]='h00000e24;
    rd_cycle[ 1280] = 1'b0;  wr_cycle[ 1280] = 1'b1;  addr_rom[ 1280]='h00001400;  wr_data_rom[ 1280]='h00002511;
    rd_cycle[ 1281] = 1'b0;  wr_cycle[ 1281] = 1'b1;  addr_rom[ 1281]='h00001404;  wr_data_rom[ 1281]='h00002764;
    rd_cycle[ 1282] = 1'b0;  wr_cycle[ 1282] = 1'b1;  addr_rom[ 1282]='h00001408;  wr_data_rom[ 1282]='h00001fc8;
    rd_cycle[ 1283] = 1'b0;  wr_cycle[ 1283] = 1'b1;  addr_rom[ 1283]='h0000140c;  wr_data_rom[ 1283]='h000016b0;
    rd_cycle[ 1284] = 1'b0;  wr_cycle[ 1284] = 1'b1;  addr_rom[ 1284]='h00001410;  wr_data_rom[ 1284]='h00003cce;
    rd_cycle[ 1285] = 1'b0;  wr_cycle[ 1285] = 1'b1;  addr_rom[ 1285]='h00001414;  wr_data_rom[ 1285]='h00002590;
    rd_cycle[ 1286] = 1'b0;  wr_cycle[ 1286] = 1'b1;  addr_rom[ 1286]='h00001418;  wr_data_rom[ 1286]='h00001e78;
    rd_cycle[ 1287] = 1'b0;  wr_cycle[ 1287] = 1'b1;  addr_rom[ 1287]='h0000141c;  wr_data_rom[ 1287]='h000027be;
    rd_cycle[ 1288] = 1'b0;  wr_cycle[ 1288] = 1'b1;  addr_rom[ 1288]='h00001420;  wr_data_rom[ 1288]='h0000038c;
    rd_cycle[ 1289] = 1'b0;  wr_cycle[ 1289] = 1'b1;  addr_rom[ 1289]='h00001424;  wr_data_rom[ 1289]='h0000121a;
    rd_cycle[ 1290] = 1'b0;  wr_cycle[ 1290] = 1'b1;  addr_rom[ 1290]='h00001428;  wr_data_rom[ 1290]='h00002409;
    rd_cycle[ 1291] = 1'b0;  wr_cycle[ 1291] = 1'b1;  addr_rom[ 1291]='h0000142c;  wr_data_rom[ 1291]='h0000224f;
    rd_cycle[ 1292] = 1'b0;  wr_cycle[ 1292] = 1'b1;  addr_rom[ 1292]='h00001430;  wr_data_rom[ 1292]='h00001132;
    rd_cycle[ 1293] = 1'b0;  wr_cycle[ 1293] = 1'b1;  addr_rom[ 1293]='h00001434;  wr_data_rom[ 1293]='h000010ba;
    rd_cycle[ 1294] = 1'b0;  wr_cycle[ 1294] = 1'b1;  addr_rom[ 1294]='h00001438;  wr_data_rom[ 1294]='h0000372f;
    rd_cycle[ 1295] = 1'b0;  wr_cycle[ 1295] = 1'b1;  addr_rom[ 1295]='h0000143c;  wr_data_rom[ 1295]='h00002f51;
    rd_cycle[ 1296] = 1'b0;  wr_cycle[ 1296] = 1'b1;  addr_rom[ 1296]='h00001440;  wr_data_rom[ 1296]='h00001124;
    rd_cycle[ 1297] = 1'b0;  wr_cycle[ 1297] = 1'b1;  addr_rom[ 1297]='h00001444;  wr_data_rom[ 1297]='h000004ab;
    rd_cycle[ 1298] = 1'b0;  wr_cycle[ 1298] = 1'b1;  addr_rom[ 1298]='h00001448;  wr_data_rom[ 1298]='h00001f38;
    rd_cycle[ 1299] = 1'b0;  wr_cycle[ 1299] = 1'b1;  addr_rom[ 1299]='h0000144c;  wr_data_rom[ 1299]='h00003734;
    rd_cycle[ 1300] = 1'b0;  wr_cycle[ 1300] = 1'b1;  addr_rom[ 1300]='h00001450;  wr_data_rom[ 1300]='h00002517;
    rd_cycle[ 1301] = 1'b0;  wr_cycle[ 1301] = 1'b1;  addr_rom[ 1301]='h00001454;  wr_data_rom[ 1301]='h000010a3;
    rd_cycle[ 1302] = 1'b0;  wr_cycle[ 1302] = 1'b1;  addr_rom[ 1302]='h00001458;  wr_data_rom[ 1302]='h00000553;
    rd_cycle[ 1303] = 1'b0;  wr_cycle[ 1303] = 1'b1;  addr_rom[ 1303]='h0000145c;  wr_data_rom[ 1303]='h00001cc6;
    rd_cycle[ 1304] = 1'b0;  wr_cycle[ 1304] = 1'b1;  addr_rom[ 1304]='h00001460;  wr_data_rom[ 1304]='h00001f56;
    rd_cycle[ 1305] = 1'b0;  wr_cycle[ 1305] = 1'b1;  addr_rom[ 1305]='h00001464;  wr_data_rom[ 1305]='h00001abc;
    rd_cycle[ 1306] = 1'b0;  wr_cycle[ 1306] = 1'b1;  addr_rom[ 1306]='h00001468;  wr_data_rom[ 1306]='h000006d9;
    rd_cycle[ 1307] = 1'b0;  wr_cycle[ 1307] = 1'b1;  addr_rom[ 1307]='h0000146c;  wr_data_rom[ 1307]='h00003025;
    rd_cycle[ 1308] = 1'b0;  wr_cycle[ 1308] = 1'b1;  addr_rom[ 1308]='h00001470;  wr_data_rom[ 1308]='h00001b53;
    rd_cycle[ 1309] = 1'b0;  wr_cycle[ 1309] = 1'b1;  addr_rom[ 1309]='h00001474;  wr_data_rom[ 1309]='h00000823;
    rd_cycle[ 1310] = 1'b0;  wr_cycle[ 1310] = 1'b1;  addr_rom[ 1310]='h00001478;  wr_data_rom[ 1310]='h00000880;
    rd_cycle[ 1311] = 1'b0;  wr_cycle[ 1311] = 1'b1;  addr_rom[ 1311]='h0000147c;  wr_data_rom[ 1311]='h0000045b;
    rd_cycle[ 1312] = 1'b0;  wr_cycle[ 1312] = 1'b1;  addr_rom[ 1312]='h00001480;  wr_data_rom[ 1312]='h00003667;
    rd_cycle[ 1313] = 1'b0;  wr_cycle[ 1313] = 1'b1;  addr_rom[ 1313]='h00001484;  wr_data_rom[ 1313]='h00003702;
    rd_cycle[ 1314] = 1'b0;  wr_cycle[ 1314] = 1'b1;  addr_rom[ 1314]='h00001488;  wr_data_rom[ 1314]='h000002cf;
    rd_cycle[ 1315] = 1'b0;  wr_cycle[ 1315] = 1'b1;  addr_rom[ 1315]='h0000148c;  wr_data_rom[ 1315]='h00000685;
    rd_cycle[ 1316] = 1'b0;  wr_cycle[ 1316] = 1'b1;  addr_rom[ 1316]='h00001490;  wr_data_rom[ 1316]='h00001916;
    rd_cycle[ 1317] = 1'b0;  wr_cycle[ 1317] = 1'b1;  addr_rom[ 1317]='h00001494;  wr_data_rom[ 1317]='h00000346;
    rd_cycle[ 1318] = 1'b0;  wr_cycle[ 1318] = 1'b1;  addr_rom[ 1318]='h00001498;  wr_data_rom[ 1318]='h0000363e;
    rd_cycle[ 1319] = 1'b0;  wr_cycle[ 1319] = 1'b1;  addr_rom[ 1319]='h0000149c;  wr_data_rom[ 1319]='h0000070d;
    rd_cycle[ 1320] = 1'b0;  wr_cycle[ 1320] = 1'b1;  addr_rom[ 1320]='h000014a0;  wr_data_rom[ 1320]='h00003c3b;
    rd_cycle[ 1321] = 1'b0;  wr_cycle[ 1321] = 1'b1;  addr_rom[ 1321]='h000014a4;  wr_data_rom[ 1321]='h00001217;
    rd_cycle[ 1322] = 1'b0;  wr_cycle[ 1322] = 1'b1;  addr_rom[ 1322]='h000014a8;  wr_data_rom[ 1322]='h0000284b;
    rd_cycle[ 1323] = 1'b0;  wr_cycle[ 1323] = 1'b1;  addr_rom[ 1323]='h000014ac;  wr_data_rom[ 1323]='h00003c6b;
    rd_cycle[ 1324] = 1'b0;  wr_cycle[ 1324] = 1'b1;  addr_rom[ 1324]='h000014b0;  wr_data_rom[ 1324]='h0000217f;
    rd_cycle[ 1325] = 1'b0;  wr_cycle[ 1325] = 1'b1;  addr_rom[ 1325]='h000014b4;  wr_data_rom[ 1325]='h00001408;
    rd_cycle[ 1326] = 1'b0;  wr_cycle[ 1326] = 1'b1;  addr_rom[ 1326]='h000014b8;  wr_data_rom[ 1326]='h00000a33;
    rd_cycle[ 1327] = 1'b0;  wr_cycle[ 1327] = 1'b1;  addr_rom[ 1327]='h000014bc;  wr_data_rom[ 1327]='h00001eca;
    rd_cycle[ 1328] = 1'b0;  wr_cycle[ 1328] = 1'b1;  addr_rom[ 1328]='h000014c0;  wr_data_rom[ 1328]='h00003fcc;
    rd_cycle[ 1329] = 1'b0;  wr_cycle[ 1329] = 1'b1;  addr_rom[ 1329]='h000014c4;  wr_data_rom[ 1329]='h0000241d;
    rd_cycle[ 1330] = 1'b0;  wr_cycle[ 1330] = 1'b1;  addr_rom[ 1330]='h000014c8;  wr_data_rom[ 1330]='h000033b6;
    rd_cycle[ 1331] = 1'b0;  wr_cycle[ 1331] = 1'b1;  addr_rom[ 1331]='h000014cc;  wr_data_rom[ 1331]='h00003115;
    rd_cycle[ 1332] = 1'b0;  wr_cycle[ 1332] = 1'b1;  addr_rom[ 1332]='h000014d0;  wr_data_rom[ 1332]='h00001012;
    rd_cycle[ 1333] = 1'b0;  wr_cycle[ 1333] = 1'b1;  addr_rom[ 1333]='h000014d4;  wr_data_rom[ 1333]='h00000772;
    rd_cycle[ 1334] = 1'b0;  wr_cycle[ 1334] = 1'b1;  addr_rom[ 1334]='h000014d8;  wr_data_rom[ 1334]='h00000add;
    rd_cycle[ 1335] = 1'b0;  wr_cycle[ 1335] = 1'b1;  addr_rom[ 1335]='h000014dc;  wr_data_rom[ 1335]='h00002e4d;
    rd_cycle[ 1336] = 1'b0;  wr_cycle[ 1336] = 1'b1;  addr_rom[ 1336]='h000014e0;  wr_data_rom[ 1336]='h00000cea;
    rd_cycle[ 1337] = 1'b0;  wr_cycle[ 1337] = 1'b1;  addr_rom[ 1337]='h000014e4;  wr_data_rom[ 1337]='h00001f33;
    rd_cycle[ 1338] = 1'b0;  wr_cycle[ 1338] = 1'b1;  addr_rom[ 1338]='h000014e8;  wr_data_rom[ 1338]='h00000cc5;
    rd_cycle[ 1339] = 1'b0;  wr_cycle[ 1339] = 1'b1;  addr_rom[ 1339]='h000014ec;  wr_data_rom[ 1339]='h0000254b;
    rd_cycle[ 1340] = 1'b0;  wr_cycle[ 1340] = 1'b1;  addr_rom[ 1340]='h000014f0;  wr_data_rom[ 1340]='h00003285;
    rd_cycle[ 1341] = 1'b0;  wr_cycle[ 1341] = 1'b1;  addr_rom[ 1341]='h000014f4;  wr_data_rom[ 1341]='h000035a5;
    rd_cycle[ 1342] = 1'b0;  wr_cycle[ 1342] = 1'b1;  addr_rom[ 1342]='h000014f8;  wr_data_rom[ 1342]='h00003b7f;
    rd_cycle[ 1343] = 1'b0;  wr_cycle[ 1343] = 1'b1;  addr_rom[ 1343]='h000014fc;  wr_data_rom[ 1343]='h00002e8d;
    rd_cycle[ 1344] = 1'b0;  wr_cycle[ 1344] = 1'b1;  addr_rom[ 1344]='h00001500;  wr_data_rom[ 1344]='h0000181c;
    rd_cycle[ 1345] = 1'b0;  wr_cycle[ 1345] = 1'b1;  addr_rom[ 1345]='h00001504;  wr_data_rom[ 1345]='h00003fd7;
    rd_cycle[ 1346] = 1'b0;  wr_cycle[ 1346] = 1'b1;  addr_rom[ 1346]='h00001508;  wr_data_rom[ 1346]='h000001d5;
    rd_cycle[ 1347] = 1'b0;  wr_cycle[ 1347] = 1'b1;  addr_rom[ 1347]='h0000150c;  wr_data_rom[ 1347]='h0000284a;
    rd_cycle[ 1348] = 1'b0;  wr_cycle[ 1348] = 1'b1;  addr_rom[ 1348]='h00001510;  wr_data_rom[ 1348]='h00001bff;
    rd_cycle[ 1349] = 1'b0;  wr_cycle[ 1349] = 1'b1;  addr_rom[ 1349]='h00001514;  wr_data_rom[ 1349]='h00000da8;
    rd_cycle[ 1350] = 1'b0;  wr_cycle[ 1350] = 1'b1;  addr_rom[ 1350]='h00001518;  wr_data_rom[ 1350]='h00003d79;
    rd_cycle[ 1351] = 1'b0;  wr_cycle[ 1351] = 1'b1;  addr_rom[ 1351]='h0000151c;  wr_data_rom[ 1351]='h00000cbc;
    rd_cycle[ 1352] = 1'b0;  wr_cycle[ 1352] = 1'b1;  addr_rom[ 1352]='h00001520;  wr_data_rom[ 1352]='h00001c81;
    rd_cycle[ 1353] = 1'b0;  wr_cycle[ 1353] = 1'b1;  addr_rom[ 1353]='h00001524;  wr_data_rom[ 1353]='h000010f6;
    rd_cycle[ 1354] = 1'b0;  wr_cycle[ 1354] = 1'b1;  addr_rom[ 1354]='h00001528;  wr_data_rom[ 1354]='h0000309c;
    rd_cycle[ 1355] = 1'b0;  wr_cycle[ 1355] = 1'b1;  addr_rom[ 1355]='h0000152c;  wr_data_rom[ 1355]='h000027c7;
    rd_cycle[ 1356] = 1'b0;  wr_cycle[ 1356] = 1'b1;  addr_rom[ 1356]='h00001530;  wr_data_rom[ 1356]='h00000694;
    rd_cycle[ 1357] = 1'b0;  wr_cycle[ 1357] = 1'b1;  addr_rom[ 1357]='h00001534;  wr_data_rom[ 1357]='h00002454;
    rd_cycle[ 1358] = 1'b0;  wr_cycle[ 1358] = 1'b1;  addr_rom[ 1358]='h00001538;  wr_data_rom[ 1358]='h00000dbd;
    rd_cycle[ 1359] = 1'b0;  wr_cycle[ 1359] = 1'b1;  addr_rom[ 1359]='h0000153c;  wr_data_rom[ 1359]='h00001c90;
    rd_cycle[ 1360] = 1'b0;  wr_cycle[ 1360] = 1'b1;  addr_rom[ 1360]='h00001540;  wr_data_rom[ 1360]='h00002ef1;
    rd_cycle[ 1361] = 1'b0;  wr_cycle[ 1361] = 1'b1;  addr_rom[ 1361]='h00001544;  wr_data_rom[ 1361]='h00001fc4;
    rd_cycle[ 1362] = 1'b0;  wr_cycle[ 1362] = 1'b1;  addr_rom[ 1362]='h00001548;  wr_data_rom[ 1362]='h000034f1;
    rd_cycle[ 1363] = 1'b0;  wr_cycle[ 1363] = 1'b1;  addr_rom[ 1363]='h0000154c;  wr_data_rom[ 1363]='h00000b97;
    rd_cycle[ 1364] = 1'b0;  wr_cycle[ 1364] = 1'b1;  addr_rom[ 1364]='h00001550;  wr_data_rom[ 1364]='h00002233;
    rd_cycle[ 1365] = 1'b0;  wr_cycle[ 1365] = 1'b1;  addr_rom[ 1365]='h00001554;  wr_data_rom[ 1365]='h00003cf9;
    rd_cycle[ 1366] = 1'b0;  wr_cycle[ 1366] = 1'b1;  addr_rom[ 1366]='h00001558;  wr_data_rom[ 1366]='h00001f07;
    rd_cycle[ 1367] = 1'b0;  wr_cycle[ 1367] = 1'b1;  addr_rom[ 1367]='h0000155c;  wr_data_rom[ 1367]='h000027e6;
    rd_cycle[ 1368] = 1'b0;  wr_cycle[ 1368] = 1'b1;  addr_rom[ 1368]='h00001560;  wr_data_rom[ 1368]='h00001a78;
    rd_cycle[ 1369] = 1'b0;  wr_cycle[ 1369] = 1'b1;  addr_rom[ 1369]='h00001564;  wr_data_rom[ 1369]='h000021ba;
    rd_cycle[ 1370] = 1'b0;  wr_cycle[ 1370] = 1'b1;  addr_rom[ 1370]='h00001568;  wr_data_rom[ 1370]='h0000206f;
    rd_cycle[ 1371] = 1'b0;  wr_cycle[ 1371] = 1'b1;  addr_rom[ 1371]='h0000156c;  wr_data_rom[ 1371]='h00002446;
    rd_cycle[ 1372] = 1'b0;  wr_cycle[ 1372] = 1'b1;  addr_rom[ 1372]='h00001570;  wr_data_rom[ 1372]='h00003bdb;
    rd_cycle[ 1373] = 1'b0;  wr_cycle[ 1373] = 1'b1;  addr_rom[ 1373]='h00001574;  wr_data_rom[ 1373]='h00002696;
    rd_cycle[ 1374] = 1'b0;  wr_cycle[ 1374] = 1'b1;  addr_rom[ 1374]='h00001578;  wr_data_rom[ 1374]='h00002709;
    rd_cycle[ 1375] = 1'b0;  wr_cycle[ 1375] = 1'b1;  addr_rom[ 1375]='h0000157c;  wr_data_rom[ 1375]='h00000c81;
    rd_cycle[ 1376] = 1'b0;  wr_cycle[ 1376] = 1'b1;  addr_rom[ 1376]='h00001580;  wr_data_rom[ 1376]='h00002f05;
    rd_cycle[ 1377] = 1'b0;  wr_cycle[ 1377] = 1'b1;  addr_rom[ 1377]='h00001584;  wr_data_rom[ 1377]='h000029db;
    rd_cycle[ 1378] = 1'b0;  wr_cycle[ 1378] = 1'b1;  addr_rom[ 1378]='h00001588;  wr_data_rom[ 1378]='h00002056;
    rd_cycle[ 1379] = 1'b0;  wr_cycle[ 1379] = 1'b1;  addr_rom[ 1379]='h0000158c;  wr_data_rom[ 1379]='h00002bb0;
    rd_cycle[ 1380] = 1'b0;  wr_cycle[ 1380] = 1'b1;  addr_rom[ 1380]='h00001590;  wr_data_rom[ 1380]='h00002870;
    rd_cycle[ 1381] = 1'b0;  wr_cycle[ 1381] = 1'b1;  addr_rom[ 1381]='h00001594;  wr_data_rom[ 1381]='h00003d74;
    rd_cycle[ 1382] = 1'b0;  wr_cycle[ 1382] = 1'b1;  addr_rom[ 1382]='h00001598;  wr_data_rom[ 1382]='h00003c90;
    rd_cycle[ 1383] = 1'b0;  wr_cycle[ 1383] = 1'b1;  addr_rom[ 1383]='h0000159c;  wr_data_rom[ 1383]='h00000919;
    rd_cycle[ 1384] = 1'b0;  wr_cycle[ 1384] = 1'b1;  addr_rom[ 1384]='h000015a0;  wr_data_rom[ 1384]='h00002242;
    rd_cycle[ 1385] = 1'b0;  wr_cycle[ 1385] = 1'b1;  addr_rom[ 1385]='h000015a4;  wr_data_rom[ 1385]='h00002720;
    rd_cycle[ 1386] = 1'b0;  wr_cycle[ 1386] = 1'b1;  addr_rom[ 1386]='h000015a8;  wr_data_rom[ 1386]='h00000127;
    rd_cycle[ 1387] = 1'b0;  wr_cycle[ 1387] = 1'b1;  addr_rom[ 1387]='h000015ac;  wr_data_rom[ 1387]='h00000e09;
    rd_cycle[ 1388] = 1'b0;  wr_cycle[ 1388] = 1'b1;  addr_rom[ 1388]='h000015b0;  wr_data_rom[ 1388]='h00003da3;
    rd_cycle[ 1389] = 1'b0;  wr_cycle[ 1389] = 1'b1;  addr_rom[ 1389]='h000015b4;  wr_data_rom[ 1389]='h00001fcd;
    rd_cycle[ 1390] = 1'b0;  wr_cycle[ 1390] = 1'b1;  addr_rom[ 1390]='h000015b8;  wr_data_rom[ 1390]='h00000123;
    rd_cycle[ 1391] = 1'b0;  wr_cycle[ 1391] = 1'b1;  addr_rom[ 1391]='h000015bc;  wr_data_rom[ 1391]='h000008d9;
    rd_cycle[ 1392] = 1'b0;  wr_cycle[ 1392] = 1'b1;  addr_rom[ 1392]='h000015c0;  wr_data_rom[ 1392]='h00003eb1;
    rd_cycle[ 1393] = 1'b0;  wr_cycle[ 1393] = 1'b1;  addr_rom[ 1393]='h000015c4;  wr_data_rom[ 1393]='h00000013;
    rd_cycle[ 1394] = 1'b0;  wr_cycle[ 1394] = 1'b1;  addr_rom[ 1394]='h000015c8;  wr_data_rom[ 1394]='h00000b34;
    rd_cycle[ 1395] = 1'b0;  wr_cycle[ 1395] = 1'b1;  addr_rom[ 1395]='h000015cc;  wr_data_rom[ 1395]='h00000aef;
    rd_cycle[ 1396] = 1'b0;  wr_cycle[ 1396] = 1'b1;  addr_rom[ 1396]='h000015d0;  wr_data_rom[ 1396]='h00000c4d;
    rd_cycle[ 1397] = 1'b0;  wr_cycle[ 1397] = 1'b1;  addr_rom[ 1397]='h000015d4;  wr_data_rom[ 1397]='h000016c4;
    rd_cycle[ 1398] = 1'b0;  wr_cycle[ 1398] = 1'b1;  addr_rom[ 1398]='h000015d8;  wr_data_rom[ 1398]='h00002aba;
    rd_cycle[ 1399] = 1'b0;  wr_cycle[ 1399] = 1'b1;  addr_rom[ 1399]='h000015dc;  wr_data_rom[ 1399]='h00001901;
    rd_cycle[ 1400] = 1'b0;  wr_cycle[ 1400] = 1'b1;  addr_rom[ 1400]='h000015e0;  wr_data_rom[ 1400]='h0000272e;
    rd_cycle[ 1401] = 1'b0;  wr_cycle[ 1401] = 1'b1;  addr_rom[ 1401]='h000015e4;  wr_data_rom[ 1401]='h00000962;
    rd_cycle[ 1402] = 1'b0;  wr_cycle[ 1402] = 1'b1;  addr_rom[ 1402]='h000015e8;  wr_data_rom[ 1402]='h000004a6;
    rd_cycle[ 1403] = 1'b0;  wr_cycle[ 1403] = 1'b1;  addr_rom[ 1403]='h000015ec;  wr_data_rom[ 1403]='h00002121;
    rd_cycle[ 1404] = 1'b0;  wr_cycle[ 1404] = 1'b1;  addr_rom[ 1404]='h000015f0;  wr_data_rom[ 1404]='h00003606;
    rd_cycle[ 1405] = 1'b0;  wr_cycle[ 1405] = 1'b1;  addr_rom[ 1405]='h000015f4;  wr_data_rom[ 1405]='h000020f0;
    rd_cycle[ 1406] = 1'b0;  wr_cycle[ 1406] = 1'b1;  addr_rom[ 1406]='h000015f8;  wr_data_rom[ 1406]='h0000147a;
    rd_cycle[ 1407] = 1'b0;  wr_cycle[ 1407] = 1'b1;  addr_rom[ 1407]='h000015fc;  wr_data_rom[ 1407]='h00000dbb;
    rd_cycle[ 1408] = 1'b0;  wr_cycle[ 1408] = 1'b1;  addr_rom[ 1408]='h00001600;  wr_data_rom[ 1408]='h00001d55;
    rd_cycle[ 1409] = 1'b0;  wr_cycle[ 1409] = 1'b1;  addr_rom[ 1409]='h00001604;  wr_data_rom[ 1409]='h00002f24;
    rd_cycle[ 1410] = 1'b0;  wr_cycle[ 1410] = 1'b1;  addr_rom[ 1410]='h00001608;  wr_data_rom[ 1410]='h000031d2;
    rd_cycle[ 1411] = 1'b0;  wr_cycle[ 1411] = 1'b1;  addr_rom[ 1411]='h0000160c;  wr_data_rom[ 1411]='h00001274;
    rd_cycle[ 1412] = 1'b0;  wr_cycle[ 1412] = 1'b1;  addr_rom[ 1412]='h00001610;  wr_data_rom[ 1412]='h00003fd3;
    rd_cycle[ 1413] = 1'b0;  wr_cycle[ 1413] = 1'b1;  addr_rom[ 1413]='h00001614;  wr_data_rom[ 1413]='h00001cec;
    rd_cycle[ 1414] = 1'b0;  wr_cycle[ 1414] = 1'b1;  addr_rom[ 1414]='h00001618;  wr_data_rom[ 1414]='h00002a06;
    rd_cycle[ 1415] = 1'b0;  wr_cycle[ 1415] = 1'b1;  addr_rom[ 1415]='h0000161c;  wr_data_rom[ 1415]='h000007e3;
    rd_cycle[ 1416] = 1'b0;  wr_cycle[ 1416] = 1'b1;  addr_rom[ 1416]='h00001620;  wr_data_rom[ 1416]='h00002059;
    rd_cycle[ 1417] = 1'b0;  wr_cycle[ 1417] = 1'b1;  addr_rom[ 1417]='h00001624;  wr_data_rom[ 1417]='h00003ba8;
    rd_cycle[ 1418] = 1'b0;  wr_cycle[ 1418] = 1'b1;  addr_rom[ 1418]='h00001628;  wr_data_rom[ 1418]='h000037a1;
    rd_cycle[ 1419] = 1'b0;  wr_cycle[ 1419] = 1'b1;  addr_rom[ 1419]='h0000162c;  wr_data_rom[ 1419]='h00001269;
    rd_cycle[ 1420] = 1'b0;  wr_cycle[ 1420] = 1'b1;  addr_rom[ 1420]='h00001630;  wr_data_rom[ 1420]='h00001c38;
    rd_cycle[ 1421] = 1'b0;  wr_cycle[ 1421] = 1'b1;  addr_rom[ 1421]='h00001634;  wr_data_rom[ 1421]='h00000dcd;
    rd_cycle[ 1422] = 1'b0;  wr_cycle[ 1422] = 1'b1;  addr_rom[ 1422]='h00001638;  wr_data_rom[ 1422]='h000021f1;
    rd_cycle[ 1423] = 1'b0;  wr_cycle[ 1423] = 1'b1;  addr_rom[ 1423]='h0000163c;  wr_data_rom[ 1423]='h00001130;
    rd_cycle[ 1424] = 1'b0;  wr_cycle[ 1424] = 1'b1;  addr_rom[ 1424]='h00001640;  wr_data_rom[ 1424]='h000004c1;
    rd_cycle[ 1425] = 1'b0;  wr_cycle[ 1425] = 1'b1;  addr_rom[ 1425]='h00001644;  wr_data_rom[ 1425]='h000015a3;
    rd_cycle[ 1426] = 1'b0;  wr_cycle[ 1426] = 1'b1;  addr_rom[ 1426]='h00001648;  wr_data_rom[ 1426]='h000029ad;
    rd_cycle[ 1427] = 1'b0;  wr_cycle[ 1427] = 1'b1;  addr_rom[ 1427]='h0000164c;  wr_data_rom[ 1427]='h0000350f;
    rd_cycle[ 1428] = 1'b0;  wr_cycle[ 1428] = 1'b1;  addr_rom[ 1428]='h00001650;  wr_data_rom[ 1428]='h00000e80;
    rd_cycle[ 1429] = 1'b0;  wr_cycle[ 1429] = 1'b1;  addr_rom[ 1429]='h00001654;  wr_data_rom[ 1429]='h00000a0d;
    rd_cycle[ 1430] = 1'b0;  wr_cycle[ 1430] = 1'b1;  addr_rom[ 1430]='h00001658;  wr_data_rom[ 1430]='h00003a10;
    rd_cycle[ 1431] = 1'b0;  wr_cycle[ 1431] = 1'b1;  addr_rom[ 1431]='h0000165c;  wr_data_rom[ 1431]='h0000325c;
    rd_cycle[ 1432] = 1'b0;  wr_cycle[ 1432] = 1'b1;  addr_rom[ 1432]='h00001660;  wr_data_rom[ 1432]='h00003c47;
    rd_cycle[ 1433] = 1'b0;  wr_cycle[ 1433] = 1'b1;  addr_rom[ 1433]='h00001664;  wr_data_rom[ 1433]='h00003755;
    rd_cycle[ 1434] = 1'b0;  wr_cycle[ 1434] = 1'b1;  addr_rom[ 1434]='h00001668;  wr_data_rom[ 1434]='h00000a4a;
    rd_cycle[ 1435] = 1'b0;  wr_cycle[ 1435] = 1'b1;  addr_rom[ 1435]='h0000166c;  wr_data_rom[ 1435]='h0000135f;
    rd_cycle[ 1436] = 1'b0;  wr_cycle[ 1436] = 1'b1;  addr_rom[ 1436]='h00001670;  wr_data_rom[ 1436]='h000002f8;
    rd_cycle[ 1437] = 1'b0;  wr_cycle[ 1437] = 1'b1;  addr_rom[ 1437]='h00001674;  wr_data_rom[ 1437]='h0000028b;
    rd_cycle[ 1438] = 1'b0;  wr_cycle[ 1438] = 1'b1;  addr_rom[ 1438]='h00001678;  wr_data_rom[ 1438]='h0000119e;
    rd_cycle[ 1439] = 1'b0;  wr_cycle[ 1439] = 1'b1;  addr_rom[ 1439]='h0000167c;  wr_data_rom[ 1439]='h00001bd8;
    rd_cycle[ 1440] = 1'b0;  wr_cycle[ 1440] = 1'b1;  addr_rom[ 1440]='h00001680;  wr_data_rom[ 1440]='h000025ff;
    rd_cycle[ 1441] = 1'b0;  wr_cycle[ 1441] = 1'b1;  addr_rom[ 1441]='h00001684;  wr_data_rom[ 1441]='h00001f6d;
    rd_cycle[ 1442] = 1'b0;  wr_cycle[ 1442] = 1'b1;  addr_rom[ 1442]='h00001688;  wr_data_rom[ 1442]='h00003a6c;
    rd_cycle[ 1443] = 1'b0;  wr_cycle[ 1443] = 1'b1;  addr_rom[ 1443]='h0000168c;  wr_data_rom[ 1443]='h000009be;
    rd_cycle[ 1444] = 1'b0;  wr_cycle[ 1444] = 1'b1;  addr_rom[ 1444]='h00001690;  wr_data_rom[ 1444]='h00003a1a;
    rd_cycle[ 1445] = 1'b0;  wr_cycle[ 1445] = 1'b1;  addr_rom[ 1445]='h00001694;  wr_data_rom[ 1445]='h00002876;
    rd_cycle[ 1446] = 1'b0;  wr_cycle[ 1446] = 1'b1;  addr_rom[ 1446]='h00001698;  wr_data_rom[ 1446]='h00003a9b;
    rd_cycle[ 1447] = 1'b0;  wr_cycle[ 1447] = 1'b1;  addr_rom[ 1447]='h0000169c;  wr_data_rom[ 1447]='h00001af6;
    rd_cycle[ 1448] = 1'b0;  wr_cycle[ 1448] = 1'b1;  addr_rom[ 1448]='h000016a0;  wr_data_rom[ 1448]='h0000274a;
    rd_cycle[ 1449] = 1'b0;  wr_cycle[ 1449] = 1'b1;  addr_rom[ 1449]='h000016a4;  wr_data_rom[ 1449]='h00000b6b;
    rd_cycle[ 1450] = 1'b0;  wr_cycle[ 1450] = 1'b1;  addr_rom[ 1450]='h000016a8;  wr_data_rom[ 1450]='h00002897;
    rd_cycle[ 1451] = 1'b0;  wr_cycle[ 1451] = 1'b1;  addr_rom[ 1451]='h000016ac;  wr_data_rom[ 1451]='h00003c87;
    rd_cycle[ 1452] = 1'b0;  wr_cycle[ 1452] = 1'b1;  addr_rom[ 1452]='h000016b0;  wr_data_rom[ 1452]='h00001149;
    rd_cycle[ 1453] = 1'b0;  wr_cycle[ 1453] = 1'b1;  addr_rom[ 1453]='h000016b4;  wr_data_rom[ 1453]='h00000471;
    rd_cycle[ 1454] = 1'b0;  wr_cycle[ 1454] = 1'b1;  addr_rom[ 1454]='h000016b8;  wr_data_rom[ 1454]='h00001af9;
    rd_cycle[ 1455] = 1'b0;  wr_cycle[ 1455] = 1'b1;  addr_rom[ 1455]='h000016bc;  wr_data_rom[ 1455]='h00001752;
    rd_cycle[ 1456] = 1'b0;  wr_cycle[ 1456] = 1'b1;  addr_rom[ 1456]='h000016c0;  wr_data_rom[ 1456]='h000027d5;
    rd_cycle[ 1457] = 1'b0;  wr_cycle[ 1457] = 1'b1;  addr_rom[ 1457]='h000016c4;  wr_data_rom[ 1457]='h0000007e;
    rd_cycle[ 1458] = 1'b0;  wr_cycle[ 1458] = 1'b1;  addr_rom[ 1458]='h000016c8;  wr_data_rom[ 1458]='h00003719;
    rd_cycle[ 1459] = 1'b0;  wr_cycle[ 1459] = 1'b1;  addr_rom[ 1459]='h000016cc;  wr_data_rom[ 1459]='h000029af;
    rd_cycle[ 1460] = 1'b0;  wr_cycle[ 1460] = 1'b1;  addr_rom[ 1460]='h000016d0;  wr_data_rom[ 1460]='h00003419;
    rd_cycle[ 1461] = 1'b0;  wr_cycle[ 1461] = 1'b1;  addr_rom[ 1461]='h000016d4;  wr_data_rom[ 1461]='h000024fc;
    rd_cycle[ 1462] = 1'b0;  wr_cycle[ 1462] = 1'b1;  addr_rom[ 1462]='h000016d8;  wr_data_rom[ 1462]='h00003ee4;
    rd_cycle[ 1463] = 1'b0;  wr_cycle[ 1463] = 1'b1;  addr_rom[ 1463]='h000016dc;  wr_data_rom[ 1463]='h000004a6;
    rd_cycle[ 1464] = 1'b0;  wr_cycle[ 1464] = 1'b1;  addr_rom[ 1464]='h000016e0;  wr_data_rom[ 1464]='h00001078;
    rd_cycle[ 1465] = 1'b0;  wr_cycle[ 1465] = 1'b1;  addr_rom[ 1465]='h000016e4;  wr_data_rom[ 1465]='h00001c94;
    rd_cycle[ 1466] = 1'b0;  wr_cycle[ 1466] = 1'b1;  addr_rom[ 1466]='h000016e8;  wr_data_rom[ 1466]='h0000153d;
    rd_cycle[ 1467] = 1'b0;  wr_cycle[ 1467] = 1'b1;  addr_rom[ 1467]='h000016ec;  wr_data_rom[ 1467]='h00002a51;
    rd_cycle[ 1468] = 1'b0;  wr_cycle[ 1468] = 1'b1;  addr_rom[ 1468]='h000016f0;  wr_data_rom[ 1468]='h00002687;
    rd_cycle[ 1469] = 1'b0;  wr_cycle[ 1469] = 1'b1;  addr_rom[ 1469]='h000016f4;  wr_data_rom[ 1469]='h00000c05;
    rd_cycle[ 1470] = 1'b0;  wr_cycle[ 1470] = 1'b1;  addr_rom[ 1470]='h000016f8;  wr_data_rom[ 1470]='h000032ca;
    rd_cycle[ 1471] = 1'b0;  wr_cycle[ 1471] = 1'b1;  addr_rom[ 1471]='h000016fc;  wr_data_rom[ 1471]='h00000695;
    rd_cycle[ 1472] = 1'b0;  wr_cycle[ 1472] = 1'b1;  addr_rom[ 1472]='h00001700;  wr_data_rom[ 1472]='h00003320;
    rd_cycle[ 1473] = 1'b0;  wr_cycle[ 1473] = 1'b1;  addr_rom[ 1473]='h00001704;  wr_data_rom[ 1473]='h00000af1;
    rd_cycle[ 1474] = 1'b0;  wr_cycle[ 1474] = 1'b1;  addr_rom[ 1474]='h00001708;  wr_data_rom[ 1474]='h00000815;
    rd_cycle[ 1475] = 1'b0;  wr_cycle[ 1475] = 1'b1;  addr_rom[ 1475]='h0000170c;  wr_data_rom[ 1475]='h00003169;
    rd_cycle[ 1476] = 1'b0;  wr_cycle[ 1476] = 1'b1;  addr_rom[ 1476]='h00001710;  wr_data_rom[ 1476]='h00002800;
    rd_cycle[ 1477] = 1'b0;  wr_cycle[ 1477] = 1'b1;  addr_rom[ 1477]='h00001714;  wr_data_rom[ 1477]='h000002af;
    rd_cycle[ 1478] = 1'b0;  wr_cycle[ 1478] = 1'b1;  addr_rom[ 1478]='h00001718;  wr_data_rom[ 1478]='h000004c2;
    rd_cycle[ 1479] = 1'b0;  wr_cycle[ 1479] = 1'b1;  addr_rom[ 1479]='h0000171c;  wr_data_rom[ 1479]='h000037b4;
    rd_cycle[ 1480] = 1'b0;  wr_cycle[ 1480] = 1'b1;  addr_rom[ 1480]='h00001720;  wr_data_rom[ 1480]='h000008f1;
    rd_cycle[ 1481] = 1'b0;  wr_cycle[ 1481] = 1'b1;  addr_rom[ 1481]='h00001724;  wr_data_rom[ 1481]='h00003251;
    rd_cycle[ 1482] = 1'b0;  wr_cycle[ 1482] = 1'b1;  addr_rom[ 1482]='h00001728;  wr_data_rom[ 1482]='h00001789;
    rd_cycle[ 1483] = 1'b0;  wr_cycle[ 1483] = 1'b1;  addr_rom[ 1483]='h0000172c;  wr_data_rom[ 1483]='h00000d54;
    rd_cycle[ 1484] = 1'b0;  wr_cycle[ 1484] = 1'b1;  addr_rom[ 1484]='h00001730;  wr_data_rom[ 1484]='h00003e80;
    rd_cycle[ 1485] = 1'b0;  wr_cycle[ 1485] = 1'b1;  addr_rom[ 1485]='h00001734;  wr_data_rom[ 1485]='h00002eb3;
    rd_cycle[ 1486] = 1'b0;  wr_cycle[ 1486] = 1'b1;  addr_rom[ 1486]='h00001738;  wr_data_rom[ 1486]='h000016fa;
    rd_cycle[ 1487] = 1'b0;  wr_cycle[ 1487] = 1'b1;  addr_rom[ 1487]='h0000173c;  wr_data_rom[ 1487]='h00001fd7;
    rd_cycle[ 1488] = 1'b0;  wr_cycle[ 1488] = 1'b1;  addr_rom[ 1488]='h00001740;  wr_data_rom[ 1488]='h00000713;
    rd_cycle[ 1489] = 1'b0;  wr_cycle[ 1489] = 1'b1;  addr_rom[ 1489]='h00001744;  wr_data_rom[ 1489]='h000018e1;
    rd_cycle[ 1490] = 1'b0;  wr_cycle[ 1490] = 1'b1;  addr_rom[ 1490]='h00001748;  wr_data_rom[ 1490]='h00002350;
    rd_cycle[ 1491] = 1'b0;  wr_cycle[ 1491] = 1'b1;  addr_rom[ 1491]='h0000174c;  wr_data_rom[ 1491]='h00000269;
    rd_cycle[ 1492] = 1'b0;  wr_cycle[ 1492] = 1'b1;  addr_rom[ 1492]='h00001750;  wr_data_rom[ 1492]='h00003d68;
    rd_cycle[ 1493] = 1'b0;  wr_cycle[ 1493] = 1'b1;  addr_rom[ 1493]='h00001754;  wr_data_rom[ 1493]='h00000b84;
    rd_cycle[ 1494] = 1'b0;  wr_cycle[ 1494] = 1'b1;  addr_rom[ 1494]='h00001758;  wr_data_rom[ 1494]='h00000f7b;
    rd_cycle[ 1495] = 1'b0;  wr_cycle[ 1495] = 1'b1;  addr_rom[ 1495]='h0000175c;  wr_data_rom[ 1495]='h00000a45;
    rd_cycle[ 1496] = 1'b0;  wr_cycle[ 1496] = 1'b1;  addr_rom[ 1496]='h00001760;  wr_data_rom[ 1496]='h00002904;
    rd_cycle[ 1497] = 1'b0;  wr_cycle[ 1497] = 1'b1;  addr_rom[ 1497]='h00001764;  wr_data_rom[ 1497]='h000004fb;
    rd_cycle[ 1498] = 1'b0;  wr_cycle[ 1498] = 1'b1;  addr_rom[ 1498]='h00001768;  wr_data_rom[ 1498]='h000033f6;
    rd_cycle[ 1499] = 1'b0;  wr_cycle[ 1499] = 1'b1;  addr_rom[ 1499]='h0000176c;  wr_data_rom[ 1499]='h00000e19;
    rd_cycle[ 1500] = 1'b0;  wr_cycle[ 1500] = 1'b1;  addr_rom[ 1500]='h00001770;  wr_data_rom[ 1500]='h0000310f;
    rd_cycle[ 1501] = 1'b0;  wr_cycle[ 1501] = 1'b1;  addr_rom[ 1501]='h00001774;  wr_data_rom[ 1501]='h000000f3;
    rd_cycle[ 1502] = 1'b0;  wr_cycle[ 1502] = 1'b1;  addr_rom[ 1502]='h00001778;  wr_data_rom[ 1502]='h00002de8;
    rd_cycle[ 1503] = 1'b0;  wr_cycle[ 1503] = 1'b1;  addr_rom[ 1503]='h0000177c;  wr_data_rom[ 1503]='h00001819;
    rd_cycle[ 1504] = 1'b0;  wr_cycle[ 1504] = 1'b1;  addr_rom[ 1504]='h00001780;  wr_data_rom[ 1504]='h00000886;
    rd_cycle[ 1505] = 1'b0;  wr_cycle[ 1505] = 1'b1;  addr_rom[ 1505]='h00001784;  wr_data_rom[ 1505]='h00003bfc;
    rd_cycle[ 1506] = 1'b0;  wr_cycle[ 1506] = 1'b1;  addr_rom[ 1506]='h00001788;  wr_data_rom[ 1506]='h00003940;
    rd_cycle[ 1507] = 1'b0;  wr_cycle[ 1507] = 1'b1;  addr_rom[ 1507]='h0000178c;  wr_data_rom[ 1507]='h00003194;
    rd_cycle[ 1508] = 1'b0;  wr_cycle[ 1508] = 1'b1;  addr_rom[ 1508]='h00001790;  wr_data_rom[ 1508]='h00002f5c;
    rd_cycle[ 1509] = 1'b0;  wr_cycle[ 1509] = 1'b1;  addr_rom[ 1509]='h00001794;  wr_data_rom[ 1509]='h0000075a;
    rd_cycle[ 1510] = 1'b0;  wr_cycle[ 1510] = 1'b1;  addr_rom[ 1510]='h00001798;  wr_data_rom[ 1510]='h000030c5;
    rd_cycle[ 1511] = 1'b0;  wr_cycle[ 1511] = 1'b1;  addr_rom[ 1511]='h0000179c;  wr_data_rom[ 1511]='h000003df;
    rd_cycle[ 1512] = 1'b0;  wr_cycle[ 1512] = 1'b1;  addr_rom[ 1512]='h000017a0;  wr_data_rom[ 1512]='h00002425;
    rd_cycle[ 1513] = 1'b0;  wr_cycle[ 1513] = 1'b1;  addr_rom[ 1513]='h000017a4;  wr_data_rom[ 1513]='h00001864;
    rd_cycle[ 1514] = 1'b0;  wr_cycle[ 1514] = 1'b1;  addr_rom[ 1514]='h000017a8;  wr_data_rom[ 1514]='h000033d2;
    rd_cycle[ 1515] = 1'b0;  wr_cycle[ 1515] = 1'b1;  addr_rom[ 1515]='h000017ac;  wr_data_rom[ 1515]='h00000c96;
    rd_cycle[ 1516] = 1'b0;  wr_cycle[ 1516] = 1'b1;  addr_rom[ 1516]='h000017b0;  wr_data_rom[ 1516]='h000003b0;
    rd_cycle[ 1517] = 1'b0;  wr_cycle[ 1517] = 1'b1;  addr_rom[ 1517]='h000017b4;  wr_data_rom[ 1517]='h000015df;
    rd_cycle[ 1518] = 1'b0;  wr_cycle[ 1518] = 1'b1;  addr_rom[ 1518]='h000017b8;  wr_data_rom[ 1518]='h00001839;
    rd_cycle[ 1519] = 1'b0;  wr_cycle[ 1519] = 1'b1;  addr_rom[ 1519]='h000017bc;  wr_data_rom[ 1519]='h00001817;
    rd_cycle[ 1520] = 1'b0;  wr_cycle[ 1520] = 1'b1;  addr_rom[ 1520]='h000017c0;  wr_data_rom[ 1520]='h00000862;
    rd_cycle[ 1521] = 1'b0;  wr_cycle[ 1521] = 1'b1;  addr_rom[ 1521]='h000017c4;  wr_data_rom[ 1521]='h0000380d;
    rd_cycle[ 1522] = 1'b0;  wr_cycle[ 1522] = 1'b1;  addr_rom[ 1522]='h000017c8;  wr_data_rom[ 1522]='h00003f5b;
    rd_cycle[ 1523] = 1'b0;  wr_cycle[ 1523] = 1'b1;  addr_rom[ 1523]='h000017cc;  wr_data_rom[ 1523]='h00000fb7;
    rd_cycle[ 1524] = 1'b0;  wr_cycle[ 1524] = 1'b1;  addr_rom[ 1524]='h000017d0;  wr_data_rom[ 1524]='h000024c9;
    rd_cycle[ 1525] = 1'b0;  wr_cycle[ 1525] = 1'b1;  addr_rom[ 1525]='h000017d4;  wr_data_rom[ 1525]='h00002f54;
    rd_cycle[ 1526] = 1'b0;  wr_cycle[ 1526] = 1'b1;  addr_rom[ 1526]='h000017d8;  wr_data_rom[ 1526]='h00001580;
    rd_cycle[ 1527] = 1'b0;  wr_cycle[ 1527] = 1'b1;  addr_rom[ 1527]='h000017dc;  wr_data_rom[ 1527]='h0000279d;
    rd_cycle[ 1528] = 1'b0;  wr_cycle[ 1528] = 1'b1;  addr_rom[ 1528]='h000017e0;  wr_data_rom[ 1528]='h00001527;
    rd_cycle[ 1529] = 1'b0;  wr_cycle[ 1529] = 1'b1;  addr_rom[ 1529]='h000017e4;  wr_data_rom[ 1529]='h00001f8f;
    rd_cycle[ 1530] = 1'b0;  wr_cycle[ 1530] = 1'b1;  addr_rom[ 1530]='h000017e8;  wr_data_rom[ 1530]='h00000c1d;
    rd_cycle[ 1531] = 1'b0;  wr_cycle[ 1531] = 1'b1;  addr_rom[ 1531]='h000017ec;  wr_data_rom[ 1531]='h000013f8;
    rd_cycle[ 1532] = 1'b0;  wr_cycle[ 1532] = 1'b1;  addr_rom[ 1532]='h000017f0;  wr_data_rom[ 1532]='h00000853;
    rd_cycle[ 1533] = 1'b0;  wr_cycle[ 1533] = 1'b1;  addr_rom[ 1533]='h000017f4;  wr_data_rom[ 1533]='h00002005;
    rd_cycle[ 1534] = 1'b0;  wr_cycle[ 1534] = 1'b1;  addr_rom[ 1534]='h000017f8;  wr_data_rom[ 1534]='h00003ac2;
    rd_cycle[ 1535] = 1'b0;  wr_cycle[ 1535] = 1'b1;  addr_rom[ 1535]='h000017fc;  wr_data_rom[ 1535]='h000017eb;
    rd_cycle[ 1536] = 1'b0;  wr_cycle[ 1536] = 1'b1;  addr_rom[ 1536]='h00001800;  wr_data_rom[ 1536]='h00000af2;
    rd_cycle[ 1537] = 1'b0;  wr_cycle[ 1537] = 1'b1;  addr_rom[ 1537]='h00001804;  wr_data_rom[ 1537]='h00003ab1;
    rd_cycle[ 1538] = 1'b0;  wr_cycle[ 1538] = 1'b1;  addr_rom[ 1538]='h00001808;  wr_data_rom[ 1538]='h00002a7b;
    rd_cycle[ 1539] = 1'b0;  wr_cycle[ 1539] = 1'b1;  addr_rom[ 1539]='h0000180c;  wr_data_rom[ 1539]='h000002c9;
    rd_cycle[ 1540] = 1'b0;  wr_cycle[ 1540] = 1'b1;  addr_rom[ 1540]='h00001810;  wr_data_rom[ 1540]='h00002f45;
    rd_cycle[ 1541] = 1'b0;  wr_cycle[ 1541] = 1'b1;  addr_rom[ 1541]='h00001814;  wr_data_rom[ 1541]='h00003e78;
    rd_cycle[ 1542] = 1'b0;  wr_cycle[ 1542] = 1'b1;  addr_rom[ 1542]='h00001818;  wr_data_rom[ 1542]='h00003954;
    rd_cycle[ 1543] = 1'b0;  wr_cycle[ 1543] = 1'b1;  addr_rom[ 1543]='h0000181c;  wr_data_rom[ 1543]='h00000157;
    rd_cycle[ 1544] = 1'b0;  wr_cycle[ 1544] = 1'b1;  addr_rom[ 1544]='h00001820;  wr_data_rom[ 1544]='h00002e06;
    rd_cycle[ 1545] = 1'b0;  wr_cycle[ 1545] = 1'b1;  addr_rom[ 1545]='h00001824;  wr_data_rom[ 1545]='h0000083f;
    rd_cycle[ 1546] = 1'b0;  wr_cycle[ 1546] = 1'b1;  addr_rom[ 1546]='h00001828;  wr_data_rom[ 1546]='h00001b7d;
    rd_cycle[ 1547] = 1'b0;  wr_cycle[ 1547] = 1'b1;  addr_rom[ 1547]='h0000182c;  wr_data_rom[ 1547]='h00003f36;
    rd_cycle[ 1548] = 1'b0;  wr_cycle[ 1548] = 1'b1;  addr_rom[ 1548]='h00001830;  wr_data_rom[ 1548]='h00003818;
    rd_cycle[ 1549] = 1'b0;  wr_cycle[ 1549] = 1'b1;  addr_rom[ 1549]='h00001834;  wr_data_rom[ 1549]='h00003ca6;
    rd_cycle[ 1550] = 1'b0;  wr_cycle[ 1550] = 1'b1;  addr_rom[ 1550]='h00001838;  wr_data_rom[ 1550]='h00003792;
    rd_cycle[ 1551] = 1'b0;  wr_cycle[ 1551] = 1'b1;  addr_rom[ 1551]='h0000183c;  wr_data_rom[ 1551]='h000020b6;
    rd_cycle[ 1552] = 1'b0;  wr_cycle[ 1552] = 1'b1;  addr_rom[ 1552]='h00001840;  wr_data_rom[ 1552]='h00002d3c;
    rd_cycle[ 1553] = 1'b0;  wr_cycle[ 1553] = 1'b1;  addr_rom[ 1553]='h00001844;  wr_data_rom[ 1553]='h00002cb6;
    rd_cycle[ 1554] = 1'b0;  wr_cycle[ 1554] = 1'b1;  addr_rom[ 1554]='h00001848;  wr_data_rom[ 1554]='h00003f41;
    rd_cycle[ 1555] = 1'b0;  wr_cycle[ 1555] = 1'b1;  addr_rom[ 1555]='h0000184c;  wr_data_rom[ 1555]='h00002460;
    rd_cycle[ 1556] = 1'b0;  wr_cycle[ 1556] = 1'b1;  addr_rom[ 1556]='h00001850;  wr_data_rom[ 1556]='h00000251;
    rd_cycle[ 1557] = 1'b0;  wr_cycle[ 1557] = 1'b1;  addr_rom[ 1557]='h00001854;  wr_data_rom[ 1557]='h0000086d;
    rd_cycle[ 1558] = 1'b0;  wr_cycle[ 1558] = 1'b1;  addr_rom[ 1558]='h00001858;  wr_data_rom[ 1558]='h00003d5d;
    rd_cycle[ 1559] = 1'b0;  wr_cycle[ 1559] = 1'b1;  addr_rom[ 1559]='h0000185c;  wr_data_rom[ 1559]='h0000235d;
    rd_cycle[ 1560] = 1'b0;  wr_cycle[ 1560] = 1'b1;  addr_rom[ 1560]='h00001860;  wr_data_rom[ 1560]='h00002eb5;
    rd_cycle[ 1561] = 1'b0;  wr_cycle[ 1561] = 1'b1;  addr_rom[ 1561]='h00001864;  wr_data_rom[ 1561]='h00003b46;
    rd_cycle[ 1562] = 1'b0;  wr_cycle[ 1562] = 1'b1;  addr_rom[ 1562]='h00001868;  wr_data_rom[ 1562]='h000022c5;
    rd_cycle[ 1563] = 1'b0;  wr_cycle[ 1563] = 1'b1;  addr_rom[ 1563]='h0000186c;  wr_data_rom[ 1563]='h00002c75;
    rd_cycle[ 1564] = 1'b0;  wr_cycle[ 1564] = 1'b1;  addr_rom[ 1564]='h00001870;  wr_data_rom[ 1564]='h0000151e;
    rd_cycle[ 1565] = 1'b0;  wr_cycle[ 1565] = 1'b1;  addr_rom[ 1565]='h00001874;  wr_data_rom[ 1565]='h000008d2;
    rd_cycle[ 1566] = 1'b0;  wr_cycle[ 1566] = 1'b1;  addr_rom[ 1566]='h00001878;  wr_data_rom[ 1566]='h00000a6a;
    rd_cycle[ 1567] = 1'b0;  wr_cycle[ 1567] = 1'b1;  addr_rom[ 1567]='h0000187c;  wr_data_rom[ 1567]='h000034c4;
    rd_cycle[ 1568] = 1'b0;  wr_cycle[ 1568] = 1'b1;  addr_rom[ 1568]='h00001880;  wr_data_rom[ 1568]='h000013c8;
    rd_cycle[ 1569] = 1'b0;  wr_cycle[ 1569] = 1'b1;  addr_rom[ 1569]='h00001884;  wr_data_rom[ 1569]='h00000d53;
    rd_cycle[ 1570] = 1'b0;  wr_cycle[ 1570] = 1'b1;  addr_rom[ 1570]='h00001888;  wr_data_rom[ 1570]='h0000290a;
    rd_cycle[ 1571] = 1'b0;  wr_cycle[ 1571] = 1'b1;  addr_rom[ 1571]='h0000188c;  wr_data_rom[ 1571]='h00002b8d;
    rd_cycle[ 1572] = 1'b0;  wr_cycle[ 1572] = 1'b1;  addr_rom[ 1572]='h00001890;  wr_data_rom[ 1572]='h00003051;
    rd_cycle[ 1573] = 1'b0;  wr_cycle[ 1573] = 1'b1;  addr_rom[ 1573]='h00001894;  wr_data_rom[ 1573]='h00000442;
    rd_cycle[ 1574] = 1'b0;  wr_cycle[ 1574] = 1'b1;  addr_rom[ 1574]='h00001898;  wr_data_rom[ 1574]='h000014f9;
    rd_cycle[ 1575] = 1'b0;  wr_cycle[ 1575] = 1'b1;  addr_rom[ 1575]='h0000189c;  wr_data_rom[ 1575]='h0000393f;
    rd_cycle[ 1576] = 1'b0;  wr_cycle[ 1576] = 1'b1;  addr_rom[ 1576]='h000018a0;  wr_data_rom[ 1576]='h000003c6;
    rd_cycle[ 1577] = 1'b0;  wr_cycle[ 1577] = 1'b1;  addr_rom[ 1577]='h000018a4;  wr_data_rom[ 1577]='h000037a9;
    rd_cycle[ 1578] = 1'b0;  wr_cycle[ 1578] = 1'b1;  addr_rom[ 1578]='h000018a8;  wr_data_rom[ 1578]='h0000015d;
    rd_cycle[ 1579] = 1'b0;  wr_cycle[ 1579] = 1'b1;  addr_rom[ 1579]='h000018ac;  wr_data_rom[ 1579]='h000001b9;
    rd_cycle[ 1580] = 1'b0;  wr_cycle[ 1580] = 1'b1;  addr_rom[ 1580]='h000018b0;  wr_data_rom[ 1580]='h00002d1e;
    rd_cycle[ 1581] = 1'b0;  wr_cycle[ 1581] = 1'b1;  addr_rom[ 1581]='h000018b4;  wr_data_rom[ 1581]='h00003522;
    rd_cycle[ 1582] = 1'b0;  wr_cycle[ 1582] = 1'b1;  addr_rom[ 1582]='h000018b8;  wr_data_rom[ 1582]='h000032d4;
    rd_cycle[ 1583] = 1'b0;  wr_cycle[ 1583] = 1'b1;  addr_rom[ 1583]='h000018bc;  wr_data_rom[ 1583]='h0000383a;
    rd_cycle[ 1584] = 1'b0;  wr_cycle[ 1584] = 1'b1;  addr_rom[ 1584]='h000018c0;  wr_data_rom[ 1584]='h000037a0;
    rd_cycle[ 1585] = 1'b0;  wr_cycle[ 1585] = 1'b1;  addr_rom[ 1585]='h000018c4;  wr_data_rom[ 1585]='h00000f2c;
    rd_cycle[ 1586] = 1'b0;  wr_cycle[ 1586] = 1'b1;  addr_rom[ 1586]='h000018c8;  wr_data_rom[ 1586]='h00001efe;
    rd_cycle[ 1587] = 1'b0;  wr_cycle[ 1587] = 1'b1;  addr_rom[ 1587]='h000018cc;  wr_data_rom[ 1587]='h00000dff;
    rd_cycle[ 1588] = 1'b0;  wr_cycle[ 1588] = 1'b1;  addr_rom[ 1588]='h000018d0;  wr_data_rom[ 1588]='h000035ca;
    rd_cycle[ 1589] = 1'b0;  wr_cycle[ 1589] = 1'b1;  addr_rom[ 1589]='h000018d4;  wr_data_rom[ 1589]='h0000326f;
    rd_cycle[ 1590] = 1'b0;  wr_cycle[ 1590] = 1'b1;  addr_rom[ 1590]='h000018d8;  wr_data_rom[ 1590]='h0000233c;
    rd_cycle[ 1591] = 1'b0;  wr_cycle[ 1591] = 1'b1;  addr_rom[ 1591]='h000018dc;  wr_data_rom[ 1591]='h000032e8;
    rd_cycle[ 1592] = 1'b0;  wr_cycle[ 1592] = 1'b1;  addr_rom[ 1592]='h000018e0;  wr_data_rom[ 1592]='h00002655;
    rd_cycle[ 1593] = 1'b0;  wr_cycle[ 1593] = 1'b1;  addr_rom[ 1593]='h000018e4;  wr_data_rom[ 1593]='h00000770;
    rd_cycle[ 1594] = 1'b0;  wr_cycle[ 1594] = 1'b1;  addr_rom[ 1594]='h000018e8;  wr_data_rom[ 1594]='h000014b0;
    rd_cycle[ 1595] = 1'b0;  wr_cycle[ 1595] = 1'b1;  addr_rom[ 1595]='h000018ec;  wr_data_rom[ 1595]='h00000839;
    rd_cycle[ 1596] = 1'b0;  wr_cycle[ 1596] = 1'b1;  addr_rom[ 1596]='h000018f0;  wr_data_rom[ 1596]='h000038f8;
    rd_cycle[ 1597] = 1'b0;  wr_cycle[ 1597] = 1'b1;  addr_rom[ 1597]='h000018f4;  wr_data_rom[ 1597]='h00000e37;
    rd_cycle[ 1598] = 1'b0;  wr_cycle[ 1598] = 1'b1;  addr_rom[ 1598]='h000018f8;  wr_data_rom[ 1598]='h00000644;
    rd_cycle[ 1599] = 1'b0;  wr_cycle[ 1599] = 1'b1;  addr_rom[ 1599]='h000018fc;  wr_data_rom[ 1599]='h00002f03;
    rd_cycle[ 1600] = 1'b0;  wr_cycle[ 1600] = 1'b1;  addr_rom[ 1600]='h00001900;  wr_data_rom[ 1600]='h00001616;
    rd_cycle[ 1601] = 1'b0;  wr_cycle[ 1601] = 1'b1;  addr_rom[ 1601]='h00001904;  wr_data_rom[ 1601]='h000015b0;
    rd_cycle[ 1602] = 1'b0;  wr_cycle[ 1602] = 1'b1;  addr_rom[ 1602]='h00001908;  wr_data_rom[ 1602]='h00000b6b;
    rd_cycle[ 1603] = 1'b0;  wr_cycle[ 1603] = 1'b1;  addr_rom[ 1603]='h0000190c;  wr_data_rom[ 1603]='h00001777;
    rd_cycle[ 1604] = 1'b0;  wr_cycle[ 1604] = 1'b1;  addr_rom[ 1604]='h00001910;  wr_data_rom[ 1604]='h00003b1f;
    rd_cycle[ 1605] = 1'b0;  wr_cycle[ 1605] = 1'b1;  addr_rom[ 1605]='h00001914;  wr_data_rom[ 1605]='h00001858;
    rd_cycle[ 1606] = 1'b0;  wr_cycle[ 1606] = 1'b1;  addr_rom[ 1606]='h00001918;  wr_data_rom[ 1606]='h000024b1;
    rd_cycle[ 1607] = 1'b0;  wr_cycle[ 1607] = 1'b1;  addr_rom[ 1607]='h0000191c;  wr_data_rom[ 1607]='h000031a2;
    rd_cycle[ 1608] = 1'b0;  wr_cycle[ 1608] = 1'b1;  addr_rom[ 1608]='h00001920;  wr_data_rom[ 1608]='h000034a9;
    rd_cycle[ 1609] = 1'b0;  wr_cycle[ 1609] = 1'b1;  addr_rom[ 1609]='h00001924;  wr_data_rom[ 1609]='h0000145c;
    rd_cycle[ 1610] = 1'b0;  wr_cycle[ 1610] = 1'b1;  addr_rom[ 1610]='h00001928;  wr_data_rom[ 1610]='h00001ab3;
    rd_cycle[ 1611] = 1'b0;  wr_cycle[ 1611] = 1'b1;  addr_rom[ 1611]='h0000192c;  wr_data_rom[ 1611]='h00000936;
    rd_cycle[ 1612] = 1'b0;  wr_cycle[ 1612] = 1'b1;  addr_rom[ 1612]='h00001930;  wr_data_rom[ 1612]='h00000671;
    rd_cycle[ 1613] = 1'b0;  wr_cycle[ 1613] = 1'b1;  addr_rom[ 1613]='h00001934;  wr_data_rom[ 1613]='h000019ad;
    rd_cycle[ 1614] = 1'b0;  wr_cycle[ 1614] = 1'b1;  addr_rom[ 1614]='h00001938;  wr_data_rom[ 1614]='h00003763;
    rd_cycle[ 1615] = 1'b0;  wr_cycle[ 1615] = 1'b1;  addr_rom[ 1615]='h0000193c;  wr_data_rom[ 1615]='h00000f7f;
    rd_cycle[ 1616] = 1'b0;  wr_cycle[ 1616] = 1'b1;  addr_rom[ 1616]='h00001940;  wr_data_rom[ 1616]='h00003bcf;
    rd_cycle[ 1617] = 1'b0;  wr_cycle[ 1617] = 1'b1;  addr_rom[ 1617]='h00001944;  wr_data_rom[ 1617]='h0000333f;
    rd_cycle[ 1618] = 1'b0;  wr_cycle[ 1618] = 1'b1;  addr_rom[ 1618]='h00001948;  wr_data_rom[ 1618]='h00003165;
    rd_cycle[ 1619] = 1'b0;  wr_cycle[ 1619] = 1'b1;  addr_rom[ 1619]='h0000194c;  wr_data_rom[ 1619]='h00003f1f;
    rd_cycle[ 1620] = 1'b0;  wr_cycle[ 1620] = 1'b1;  addr_rom[ 1620]='h00001950;  wr_data_rom[ 1620]='h000034d7;
    rd_cycle[ 1621] = 1'b0;  wr_cycle[ 1621] = 1'b1;  addr_rom[ 1621]='h00001954;  wr_data_rom[ 1621]='h0000372a;
    rd_cycle[ 1622] = 1'b0;  wr_cycle[ 1622] = 1'b1;  addr_rom[ 1622]='h00001958;  wr_data_rom[ 1622]='h000004d8;
    rd_cycle[ 1623] = 1'b0;  wr_cycle[ 1623] = 1'b1;  addr_rom[ 1623]='h0000195c;  wr_data_rom[ 1623]='h000016c5;
    rd_cycle[ 1624] = 1'b0;  wr_cycle[ 1624] = 1'b1;  addr_rom[ 1624]='h00001960;  wr_data_rom[ 1624]='h000005f9;
    rd_cycle[ 1625] = 1'b0;  wr_cycle[ 1625] = 1'b1;  addr_rom[ 1625]='h00001964;  wr_data_rom[ 1625]='h000010e2;
    rd_cycle[ 1626] = 1'b0;  wr_cycle[ 1626] = 1'b1;  addr_rom[ 1626]='h00001968;  wr_data_rom[ 1626]='h00002269;
    rd_cycle[ 1627] = 1'b0;  wr_cycle[ 1627] = 1'b1;  addr_rom[ 1627]='h0000196c;  wr_data_rom[ 1627]='h00003b5b;
    rd_cycle[ 1628] = 1'b0;  wr_cycle[ 1628] = 1'b1;  addr_rom[ 1628]='h00001970;  wr_data_rom[ 1628]='h00001813;
    rd_cycle[ 1629] = 1'b0;  wr_cycle[ 1629] = 1'b1;  addr_rom[ 1629]='h00001974;  wr_data_rom[ 1629]='h00001966;
    rd_cycle[ 1630] = 1'b0;  wr_cycle[ 1630] = 1'b1;  addr_rom[ 1630]='h00001978;  wr_data_rom[ 1630]='h00001bca;
    rd_cycle[ 1631] = 1'b0;  wr_cycle[ 1631] = 1'b1;  addr_rom[ 1631]='h0000197c;  wr_data_rom[ 1631]='h00002d3a;
    rd_cycle[ 1632] = 1'b0;  wr_cycle[ 1632] = 1'b1;  addr_rom[ 1632]='h00001980;  wr_data_rom[ 1632]='h00001231;
    rd_cycle[ 1633] = 1'b0;  wr_cycle[ 1633] = 1'b1;  addr_rom[ 1633]='h00001984;  wr_data_rom[ 1633]='h000035f7;
    rd_cycle[ 1634] = 1'b0;  wr_cycle[ 1634] = 1'b1;  addr_rom[ 1634]='h00001988;  wr_data_rom[ 1634]='h0000065e;
    rd_cycle[ 1635] = 1'b0;  wr_cycle[ 1635] = 1'b1;  addr_rom[ 1635]='h0000198c;  wr_data_rom[ 1635]='h00001558;
    rd_cycle[ 1636] = 1'b0;  wr_cycle[ 1636] = 1'b1;  addr_rom[ 1636]='h00001990;  wr_data_rom[ 1636]='h00003ce0;
    rd_cycle[ 1637] = 1'b0;  wr_cycle[ 1637] = 1'b1;  addr_rom[ 1637]='h00001994;  wr_data_rom[ 1637]='h00000c50;
    rd_cycle[ 1638] = 1'b0;  wr_cycle[ 1638] = 1'b1;  addr_rom[ 1638]='h00001998;  wr_data_rom[ 1638]='h000007e8;
    rd_cycle[ 1639] = 1'b0;  wr_cycle[ 1639] = 1'b1;  addr_rom[ 1639]='h0000199c;  wr_data_rom[ 1639]='h00003b40;
    rd_cycle[ 1640] = 1'b0;  wr_cycle[ 1640] = 1'b1;  addr_rom[ 1640]='h000019a0;  wr_data_rom[ 1640]='h00002226;
    rd_cycle[ 1641] = 1'b0;  wr_cycle[ 1641] = 1'b1;  addr_rom[ 1641]='h000019a4;  wr_data_rom[ 1641]='h00001e92;
    rd_cycle[ 1642] = 1'b0;  wr_cycle[ 1642] = 1'b1;  addr_rom[ 1642]='h000019a8;  wr_data_rom[ 1642]='h00000915;
    rd_cycle[ 1643] = 1'b0;  wr_cycle[ 1643] = 1'b1;  addr_rom[ 1643]='h000019ac;  wr_data_rom[ 1643]='h000012ee;
    rd_cycle[ 1644] = 1'b0;  wr_cycle[ 1644] = 1'b1;  addr_rom[ 1644]='h000019b0;  wr_data_rom[ 1644]='h00002506;
    rd_cycle[ 1645] = 1'b0;  wr_cycle[ 1645] = 1'b1;  addr_rom[ 1645]='h000019b4;  wr_data_rom[ 1645]='h00002e00;
    rd_cycle[ 1646] = 1'b0;  wr_cycle[ 1646] = 1'b1;  addr_rom[ 1646]='h000019b8;  wr_data_rom[ 1646]='h00003615;
    rd_cycle[ 1647] = 1'b0;  wr_cycle[ 1647] = 1'b1;  addr_rom[ 1647]='h000019bc;  wr_data_rom[ 1647]='h00000e22;
    rd_cycle[ 1648] = 1'b0;  wr_cycle[ 1648] = 1'b1;  addr_rom[ 1648]='h000019c0;  wr_data_rom[ 1648]='h000037fd;
    rd_cycle[ 1649] = 1'b0;  wr_cycle[ 1649] = 1'b1;  addr_rom[ 1649]='h000019c4;  wr_data_rom[ 1649]='h0000142b;
    rd_cycle[ 1650] = 1'b0;  wr_cycle[ 1650] = 1'b1;  addr_rom[ 1650]='h000019c8;  wr_data_rom[ 1650]='h000030a5;
    rd_cycle[ 1651] = 1'b0;  wr_cycle[ 1651] = 1'b1;  addr_rom[ 1651]='h000019cc;  wr_data_rom[ 1651]='h000004c0;
    rd_cycle[ 1652] = 1'b0;  wr_cycle[ 1652] = 1'b1;  addr_rom[ 1652]='h000019d0;  wr_data_rom[ 1652]='h00002e60;
    rd_cycle[ 1653] = 1'b0;  wr_cycle[ 1653] = 1'b1;  addr_rom[ 1653]='h000019d4;  wr_data_rom[ 1653]='h00001391;
    rd_cycle[ 1654] = 1'b0;  wr_cycle[ 1654] = 1'b1;  addr_rom[ 1654]='h000019d8;  wr_data_rom[ 1654]='h00000523;
    rd_cycle[ 1655] = 1'b0;  wr_cycle[ 1655] = 1'b1;  addr_rom[ 1655]='h000019dc;  wr_data_rom[ 1655]='h000010fb;
    rd_cycle[ 1656] = 1'b0;  wr_cycle[ 1656] = 1'b1;  addr_rom[ 1656]='h000019e0;  wr_data_rom[ 1656]='h00003d42;
    rd_cycle[ 1657] = 1'b0;  wr_cycle[ 1657] = 1'b1;  addr_rom[ 1657]='h000019e4;  wr_data_rom[ 1657]='h00003652;
    rd_cycle[ 1658] = 1'b0;  wr_cycle[ 1658] = 1'b1;  addr_rom[ 1658]='h000019e8;  wr_data_rom[ 1658]='h000018ed;
    rd_cycle[ 1659] = 1'b0;  wr_cycle[ 1659] = 1'b1;  addr_rom[ 1659]='h000019ec;  wr_data_rom[ 1659]='h00003e5c;
    rd_cycle[ 1660] = 1'b0;  wr_cycle[ 1660] = 1'b1;  addr_rom[ 1660]='h000019f0;  wr_data_rom[ 1660]='h000000fd;
    rd_cycle[ 1661] = 1'b0;  wr_cycle[ 1661] = 1'b1;  addr_rom[ 1661]='h000019f4;  wr_data_rom[ 1661]='h00002bbd;
    rd_cycle[ 1662] = 1'b0;  wr_cycle[ 1662] = 1'b1;  addr_rom[ 1662]='h000019f8;  wr_data_rom[ 1662]='h00001b74;
    rd_cycle[ 1663] = 1'b0;  wr_cycle[ 1663] = 1'b1;  addr_rom[ 1663]='h000019fc;  wr_data_rom[ 1663]='h000008b6;
    rd_cycle[ 1664] = 1'b0;  wr_cycle[ 1664] = 1'b1;  addr_rom[ 1664]='h00001a00;  wr_data_rom[ 1664]='h00003975;
    rd_cycle[ 1665] = 1'b0;  wr_cycle[ 1665] = 1'b1;  addr_rom[ 1665]='h00001a04;  wr_data_rom[ 1665]='h00001b3f;
    rd_cycle[ 1666] = 1'b0;  wr_cycle[ 1666] = 1'b1;  addr_rom[ 1666]='h00001a08;  wr_data_rom[ 1666]='h00000bef;
    rd_cycle[ 1667] = 1'b0;  wr_cycle[ 1667] = 1'b1;  addr_rom[ 1667]='h00001a0c;  wr_data_rom[ 1667]='h00001831;
    rd_cycle[ 1668] = 1'b0;  wr_cycle[ 1668] = 1'b1;  addr_rom[ 1668]='h00001a10;  wr_data_rom[ 1668]='h00000b45;
    rd_cycle[ 1669] = 1'b0;  wr_cycle[ 1669] = 1'b1;  addr_rom[ 1669]='h00001a14;  wr_data_rom[ 1669]='h00000d01;
    rd_cycle[ 1670] = 1'b0;  wr_cycle[ 1670] = 1'b1;  addr_rom[ 1670]='h00001a18;  wr_data_rom[ 1670]='h0000327e;
    rd_cycle[ 1671] = 1'b0;  wr_cycle[ 1671] = 1'b1;  addr_rom[ 1671]='h00001a1c;  wr_data_rom[ 1671]='h0000201e;
    rd_cycle[ 1672] = 1'b0;  wr_cycle[ 1672] = 1'b1;  addr_rom[ 1672]='h00001a20;  wr_data_rom[ 1672]='h00003ea6;
    rd_cycle[ 1673] = 1'b0;  wr_cycle[ 1673] = 1'b1;  addr_rom[ 1673]='h00001a24;  wr_data_rom[ 1673]='h000024c7;
    rd_cycle[ 1674] = 1'b0;  wr_cycle[ 1674] = 1'b1;  addr_rom[ 1674]='h00001a28;  wr_data_rom[ 1674]='h00003100;
    rd_cycle[ 1675] = 1'b0;  wr_cycle[ 1675] = 1'b1;  addr_rom[ 1675]='h00001a2c;  wr_data_rom[ 1675]='h0000396f;
    rd_cycle[ 1676] = 1'b0;  wr_cycle[ 1676] = 1'b1;  addr_rom[ 1676]='h00001a30;  wr_data_rom[ 1676]='h000034f1;
    rd_cycle[ 1677] = 1'b0;  wr_cycle[ 1677] = 1'b1;  addr_rom[ 1677]='h00001a34;  wr_data_rom[ 1677]='h00000cc1;
    rd_cycle[ 1678] = 1'b0;  wr_cycle[ 1678] = 1'b1;  addr_rom[ 1678]='h00001a38;  wr_data_rom[ 1678]='h0000143e;
    rd_cycle[ 1679] = 1'b0;  wr_cycle[ 1679] = 1'b1;  addr_rom[ 1679]='h00001a3c;  wr_data_rom[ 1679]='h000028fc;
    rd_cycle[ 1680] = 1'b0;  wr_cycle[ 1680] = 1'b1;  addr_rom[ 1680]='h00001a40;  wr_data_rom[ 1680]='h00001263;
    rd_cycle[ 1681] = 1'b0;  wr_cycle[ 1681] = 1'b1;  addr_rom[ 1681]='h00001a44;  wr_data_rom[ 1681]='h0000246e;
    rd_cycle[ 1682] = 1'b0;  wr_cycle[ 1682] = 1'b1;  addr_rom[ 1682]='h00001a48;  wr_data_rom[ 1682]='h0000239f;
    rd_cycle[ 1683] = 1'b0;  wr_cycle[ 1683] = 1'b1;  addr_rom[ 1683]='h00001a4c;  wr_data_rom[ 1683]='h00002260;
    rd_cycle[ 1684] = 1'b0;  wr_cycle[ 1684] = 1'b1;  addr_rom[ 1684]='h00001a50;  wr_data_rom[ 1684]='h00001956;
    rd_cycle[ 1685] = 1'b0;  wr_cycle[ 1685] = 1'b1;  addr_rom[ 1685]='h00001a54;  wr_data_rom[ 1685]='h0000289b;
    rd_cycle[ 1686] = 1'b0;  wr_cycle[ 1686] = 1'b1;  addr_rom[ 1686]='h00001a58;  wr_data_rom[ 1686]='h00000d58;
    rd_cycle[ 1687] = 1'b0;  wr_cycle[ 1687] = 1'b1;  addr_rom[ 1687]='h00001a5c;  wr_data_rom[ 1687]='h000033be;
    rd_cycle[ 1688] = 1'b0;  wr_cycle[ 1688] = 1'b1;  addr_rom[ 1688]='h00001a60;  wr_data_rom[ 1688]='h00000236;
    rd_cycle[ 1689] = 1'b0;  wr_cycle[ 1689] = 1'b1;  addr_rom[ 1689]='h00001a64;  wr_data_rom[ 1689]='h00002f40;
    rd_cycle[ 1690] = 1'b0;  wr_cycle[ 1690] = 1'b1;  addr_rom[ 1690]='h00001a68;  wr_data_rom[ 1690]='h00002177;
    rd_cycle[ 1691] = 1'b0;  wr_cycle[ 1691] = 1'b1;  addr_rom[ 1691]='h00001a6c;  wr_data_rom[ 1691]='h00001891;
    rd_cycle[ 1692] = 1'b0;  wr_cycle[ 1692] = 1'b1;  addr_rom[ 1692]='h00001a70;  wr_data_rom[ 1692]='h000006ce;
    rd_cycle[ 1693] = 1'b0;  wr_cycle[ 1693] = 1'b1;  addr_rom[ 1693]='h00001a74;  wr_data_rom[ 1693]='h0000277f;
    rd_cycle[ 1694] = 1'b0;  wr_cycle[ 1694] = 1'b1;  addr_rom[ 1694]='h00001a78;  wr_data_rom[ 1694]='h0000038d;
    rd_cycle[ 1695] = 1'b0;  wr_cycle[ 1695] = 1'b1;  addr_rom[ 1695]='h00001a7c;  wr_data_rom[ 1695]='h00000472;
    rd_cycle[ 1696] = 1'b0;  wr_cycle[ 1696] = 1'b1;  addr_rom[ 1696]='h00001a80;  wr_data_rom[ 1696]='h00003eb5;
    rd_cycle[ 1697] = 1'b0;  wr_cycle[ 1697] = 1'b1;  addr_rom[ 1697]='h00001a84;  wr_data_rom[ 1697]='h000000c0;
    rd_cycle[ 1698] = 1'b0;  wr_cycle[ 1698] = 1'b1;  addr_rom[ 1698]='h00001a88;  wr_data_rom[ 1698]='h000022c2;
    rd_cycle[ 1699] = 1'b0;  wr_cycle[ 1699] = 1'b1;  addr_rom[ 1699]='h00001a8c;  wr_data_rom[ 1699]='h00002bbd;
    rd_cycle[ 1700] = 1'b0;  wr_cycle[ 1700] = 1'b1;  addr_rom[ 1700]='h00001a90;  wr_data_rom[ 1700]='h00001747;
    rd_cycle[ 1701] = 1'b0;  wr_cycle[ 1701] = 1'b1;  addr_rom[ 1701]='h00001a94;  wr_data_rom[ 1701]='h00000c4a;
    rd_cycle[ 1702] = 1'b0;  wr_cycle[ 1702] = 1'b1;  addr_rom[ 1702]='h00001a98;  wr_data_rom[ 1702]='h00001027;
    rd_cycle[ 1703] = 1'b0;  wr_cycle[ 1703] = 1'b1;  addr_rom[ 1703]='h00001a9c;  wr_data_rom[ 1703]='h0000053b;
    rd_cycle[ 1704] = 1'b0;  wr_cycle[ 1704] = 1'b1;  addr_rom[ 1704]='h00001aa0;  wr_data_rom[ 1704]='h00002355;
    rd_cycle[ 1705] = 1'b0;  wr_cycle[ 1705] = 1'b1;  addr_rom[ 1705]='h00001aa4;  wr_data_rom[ 1705]='h0000372a;
    rd_cycle[ 1706] = 1'b0;  wr_cycle[ 1706] = 1'b1;  addr_rom[ 1706]='h00001aa8;  wr_data_rom[ 1706]='h00000b98;
    rd_cycle[ 1707] = 1'b0;  wr_cycle[ 1707] = 1'b1;  addr_rom[ 1707]='h00001aac;  wr_data_rom[ 1707]='h00002088;
    rd_cycle[ 1708] = 1'b0;  wr_cycle[ 1708] = 1'b1;  addr_rom[ 1708]='h00001ab0;  wr_data_rom[ 1708]='h00003c6b;
    rd_cycle[ 1709] = 1'b0;  wr_cycle[ 1709] = 1'b1;  addr_rom[ 1709]='h00001ab4;  wr_data_rom[ 1709]='h00002b22;
    rd_cycle[ 1710] = 1'b0;  wr_cycle[ 1710] = 1'b1;  addr_rom[ 1710]='h00001ab8;  wr_data_rom[ 1710]='h00000de4;
    rd_cycle[ 1711] = 1'b0;  wr_cycle[ 1711] = 1'b1;  addr_rom[ 1711]='h00001abc;  wr_data_rom[ 1711]='h0000052e;
    rd_cycle[ 1712] = 1'b0;  wr_cycle[ 1712] = 1'b1;  addr_rom[ 1712]='h00001ac0;  wr_data_rom[ 1712]='h00001181;
    rd_cycle[ 1713] = 1'b0;  wr_cycle[ 1713] = 1'b1;  addr_rom[ 1713]='h00001ac4;  wr_data_rom[ 1713]='h00001507;
    rd_cycle[ 1714] = 1'b0;  wr_cycle[ 1714] = 1'b1;  addr_rom[ 1714]='h00001ac8;  wr_data_rom[ 1714]='h000004c1;
    rd_cycle[ 1715] = 1'b0;  wr_cycle[ 1715] = 1'b1;  addr_rom[ 1715]='h00001acc;  wr_data_rom[ 1715]='h0000105b;
    rd_cycle[ 1716] = 1'b0;  wr_cycle[ 1716] = 1'b1;  addr_rom[ 1716]='h00001ad0;  wr_data_rom[ 1716]='h00003c0f;
    rd_cycle[ 1717] = 1'b0;  wr_cycle[ 1717] = 1'b1;  addr_rom[ 1717]='h00001ad4;  wr_data_rom[ 1717]='h00003823;
    rd_cycle[ 1718] = 1'b0;  wr_cycle[ 1718] = 1'b1;  addr_rom[ 1718]='h00001ad8;  wr_data_rom[ 1718]='h00001c8d;
    rd_cycle[ 1719] = 1'b0;  wr_cycle[ 1719] = 1'b1;  addr_rom[ 1719]='h00001adc;  wr_data_rom[ 1719]='h00000fcb;
    rd_cycle[ 1720] = 1'b0;  wr_cycle[ 1720] = 1'b1;  addr_rom[ 1720]='h00001ae0;  wr_data_rom[ 1720]='h0000190e;
    rd_cycle[ 1721] = 1'b0;  wr_cycle[ 1721] = 1'b1;  addr_rom[ 1721]='h00001ae4;  wr_data_rom[ 1721]='h00003f39;
    rd_cycle[ 1722] = 1'b0;  wr_cycle[ 1722] = 1'b1;  addr_rom[ 1722]='h00001ae8;  wr_data_rom[ 1722]='h00002260;
    rd_cycle[ 1723] = 1'b0;  wr_cycle[ 1723] = 1'b1;  addr_rom[ 1723]='h00001aec;  wr_data_rom[ 1723]='h00001cd6;
    rd_cycle[ 1724] = 1'b0;  wr_cycle[ 1724] = 1'b1;  addr_rom[ 1724]='h00001af0;  wr_data_rom[ 1724]='h000031fd;
    rd_cycle[ 1725] = 1'b0;  wr_cycle[ 1725] = 1'b1;  addr_rom[ 1725]='h00001af4;  wr_data_rom[ 1725]='h00003570;
    rd_cycle[ 1726] = 1'b0;  wr_cycle[ 1726] = 1'b1;  addr_rom[ 1726]='h00001af8;  wr_data_rom[ 1726]='h00000fe4;
    rd_cycle[ 1727] = 1'b0;  wr_cycle[ 1727] = 1'b1;  addr_rom[ 1727]='h00001afc;  wr_data_rom[ 1727]='h00002347;
    rd_cycle[ 1728] = 1'b0;  wr_cycle[ 1728] = 1'b1;  addr_rom[ 1728]='h00001b00;  wr_data_rom[ 1728]='h00001229;
    rd_cycle[ 1729] = 1'b0;  wr_cycle[ 1729] = 1'b1;  addr_rom[ 1729]='h00001b04;  wr_data_rom[ 1729]='h0000275b;
    rd_cycle[ 1730] = 1'b0;  wr_cycle[ 1730] = 1'b1;  addr_rom[ 1730]='h00001b08;  wr_data_rom[ 1730]='h00001700;
    rd_cycle[ 1731] = 1'b0;  wr_cycle[ 1731] = 1'b1;  addr_rom[ 1731]='h00001b0c;  wr_data_rom[ 1731]='h00002551;
    rd_cycle[ 1732] = 1'b0;  wr_cycle[ 1732] = 1'b1;  addr_rom[ 1732]='h00001b10;  wr_data_rom[ 1732]='h00003851;
    rd_cycle[ 1733] = 1'b0;  wr_cycle[ 1733] = 1'b1;  addr_rom[ 1733]='h00001b14;  wr_data_rom[ 1733]='h00003ee6;
    rd_cycle[ 1734] = 1'b0;  wr_cycle[ 1734] = 1'b1;  addr_rom[ 1734]='h00001b18;  wr_data_rom[ 1734]='h00002a53;
    rd_cycle[ 1735] = 1'b0;  wr_cycle[ 1735] = 1'b1;  addr_rom[ 1735]='h00001b1c;  wr_data_rom[ 1735]='h000011f2;
    rd_cycle[ 1736] = 1'b0;  wr_cycle[ 1736] = 1'b1;  addr_rom[ 1736]='h00001b20;  wr_data_rom[ 1736]='h00002a9b;
    rd_cycle[ 1737] = 1'b0;  wr_cycle[ 1737] = 1'b1;  addr_rom[ 1737]='h00001b24;  wr_data_rom[ 1737]='h00002500;
    rd_cycle[ 1738] = 1'b0;  wr_cycle[ 1738] = 1'b1;  addr_rom[ 1738]='h00001b28;  wr_data_rom[ 1738]='h000030c2;
    rd_cycle[ 1739] = 1'b0;  wr_cycle[ 1739] = 1'b1;  addr_rom[ 1739]='h00001b2c;  wr_data_rom[ 1739]='h00000115;
    rd_cycle[ 1740] = 1'b0;  wr_cycle[ 1740] = 1'b1;  addr_rom[ 1740]='h00001b30;  wr_data_rom[ 1740]='h000031c1;
    rd_cycle[ 1741] = 1'b0;  wr_cycle[ 1741] = 1'b1;  addr_rom[ 1741]='h00001b34;  wr_data_rom[ 1741]='h00001d06;
    rd_cycle[ 1742] = 1'b0;  wr_cycle[ 1742] = 1'b1;  addr_rom[ 1742]='h00001b38;  wr_data_rom[ 1742]='h000028dd;
    rd_cycle[ 1743] = 1'b0;  wr_cycle[ 1743] = 1'b1;  addr_rom[ 1743]='h00001b3c;  wr_data_rom[ 1743]='h000038f7;
    rd_cycle[ 1744] = 1'b0;  wr_cycle[ 1744] = 1'b1;  addr_rom[ 1744]='h00001b40;  wr_data_rom[ 1744]='h00000fbd;
    rd_cycle[ 1745] = 1'b0;  wr_cycle[ 1745] = 1'b1;  addr_rom[ 1745]='h00001b44;  wr_data_rom[ 1745]='h0000352d;
    rd_cycle[ 1746] = 1'b0;  wr_cycle[ 1746] = 1'b1;  addr_rom[ 1746]='h00001b48;  wr_data_rom[ 1746]='h000023f8;
    rd_cycle[ 1747] = 1'b0;  wr_cycle[ 1747] = 1'b1;  addr_rom[ 1747]='h00001b4c;  wr_data_rom[ 1747]='h00003015;
    rd_cycle[ 1748] = 1'b0;  wr_cycle[ 1748] = 1'b1;  addr_rom[ 1748]='h00001b50;  wr_data_rom[ 1748]='h00001d31;
    rd_cycle[ 1749] = 1'b0;  wr_cycle[ 1749] = 1'b1;  addr_rom[ 1749]='h00001b54;  wr_data_rom[ 1749]='h000028a3;
    rd_cycle[ 1750] = 1'b0;  wr_cycle[ 1750] = 1'b1;  addr_rom[ 1750]='h00001b58;  wr_data_rom[ 1750]='h00001483;
    rd_cycle[ 1751] = 1'b0;  wr_cycle[ 1751] = 1'b1;  addr_rom[ 1751]='h00001b5c;  wr_data_rom[ 1751]='h00000dce;
    rd_cycle[ 1752] = 1'b0;  wr_cycle[ 1752] = 1'b1;  addr_rom[ 1752]='h00001b60;  wr_data_rom[ 1752]='h00001ae5;
    rd_cycle[ 1753] = 1'b0;  wr_cycle[ 1753] = 1'b1;  addr_rom[ 1753]='h00001b64;  wr_data_rom[ 1753]='h00003cb0;
    rd_cycle[ 1754] = 1'b0;  wr_cycle[ 1754] = 1'b1;  addr_rom[ 1754]='h00001b68;  wr_data_rom[ 1754]='h00000804;
    rd_cycle[ 1755] = 1'b0;  wr_cycle[ 1755] = 1'b1;  addr_rom[ 1755]='h00001b6c;  wr_data_rom[ 1755]='h00002a57;
    rd_cycle[ 1756] = 1'b0;  wr_cycle[ 1756] = 1'b1;  addr_rom[ 1756]='h00001b70;  wr_data_rom[ 1756]='h00000683;
    rd_cycle[ 1757] = 1'b0;  wr_cycle[ 1757] = 1'b1;  addr_rom[ 1757]='h00001b74;  wr_data_rom[ 1757]='h00002509;
    rd_cycle[ 1758] = 1'b0;  wr_cycle[ 1758] = 1'b1;  addr_rom[ 1758]='h00001b78;  wr_data_rom[ 1758]='h0000113d;
    rd_cycle[ 1759] = 1'b0;  wr_cycle[ 1759] = 1'b1;  addr_rom[ 1759]='h00001b7c;  wr_data_rom[ 1759]='h00000f01;
    rd_cycle[ 1760] = 1'b0;  wr_cycle[ 1760] = 1'b1;  addr_rom[ 1760]='h00001b80;  wr_data_rom[ 1760]='h000013cb;
    rd_cycle[ 1761] = 1'b0;  wr_cycle[ 1761] = 1'b1;  addr_rom[ 1761]='h00001b84;  wr_data_rom[ 1761]='h000020b3;
    rd_cycle[ 1762] = 1'b0;  wr_cycle[ 1762] = 1'b1;  addr_rom[ 1762]='h00001b88;  wr_data_rom[ 1762]='h00002b8b;
    rd_cycle[ 1763] = 1'b0;  wr_cycle[ 1763] = 1'b1;  addr_rom[ 1763]='h00001b8c;  wr_data_rom[ 1763]='h00003527;
    rd_cycle[ 1764] = 1'b0;  wr_cycle[ 1764] = 1'b1;  addr_rom[ 1764]='h00001b90;  wr_data_rom[ 1764]='h000009b5;
    rd_cycle[ 1765] = 1'b0;  wr_cycle[ 1765] = 1'b1;  addr_rom[ 1765]='h00001b94;  wr_data_rom[ 1765]='h00002731;
    rd_cycle[ 1766] = 1'b0;  wr_cycle[ 1766] = 1'b1;  addr_rom[ 1766]='h00001b98;  wr_data_rom[ 1766]='h00002625;
    rd_cycle[ 1767] = 1'b0;  wr_cycle[ 1767] = 1'b1;  addr_rom[ 1767]='h00001b9c;  wr_data_rom[ 1767]='h00001c48;
    rd_cycle[ 1768] = 1'b0;  wr_cycle[ 1768] = 1'b1;  addr_rom[ 1768]='h00001ba0;  wr_data_rom[ 1768]='h00002ada;
    rd_cycle[ 1769] = 1'b0;  wr_cycle[ 1769] = 1'b1;  addr_rom[ 1769]='h00001ba4;  wr_data_rom[ 1769]='h00003249;
    rd_cycle[ 1770] = 1'b0;  wr_cycle[ 1770] = 1'b1;  addr_rom[ 1770]='h00001ba8;  wr_data_rom[ 1770]='h00003fa6;
    rd_cycle[ 1771] = 1'b0;  wr_cycle[ 1771] = 1'b1;  addr_rom[ 1771]='h00001bac;  wr_data_rom[ 1771]='h0000238e;
    rd_cycle[ 1772] = 1'b0;  wr_cycle[ 1772] = 1'b1;  addr_rom[ 1772]='h00001bb0;  wr_data_rom[ 1772]='h00003916;
    rd_cycle[ 1773] = 1'b0;  wr_cycle[ 1773] = 1'b1;  addr_rom[ 1773]='h00001bb4;  wr_data_rom[ 1773]='h0000173a;
    rd_cycle[ 1774] = 1'b0;  wr_cycle[ 1774] = 1'b1;  addr_rom[ 1774]='h00001bb8;  wr_data_rom[ 1774]='h00002598;
    rd_cycle[ 1775] = 1'b0;  wr_cycle[ 1775] = 1'b1;  addr_rom[ 1775]='h00001bbc;  wr_data_rom[ 1775]='h000023d3;
    rd_cycle[ 1776] = 1'b0;  wr_cycle[ 1776] = 1'b1;  addr_rom[ 1776]='h00001bc0;  wr_data_rom[ 1776]='h00000654;
    rd_cycle[ 1777] = 1'b0;  wr_cycle[ 1777] = 1'b1;  addr_rom[ 1777]='h00001bc4;  wr_data_rom[ 1777]='h000003d9;
    rd_cycle[ 1778] = 1'b0;  wr_cycle[ 1778] = 1'b1;  addr_rom[ 1778]='h00001bc8;  wr_data_rom[ 1778]='h000018cd;
    rd_cycle[ 1779] = 1'b0;  wr_cycle[ 1779] = 1'b1;  addr_rom[ 1779]='h00001bcc;  wr_data_rom[ 1779]='h00002919;
    rd_cycle[ 1780] = 1'b0;  wr_cycle[ 1780] = 1'b1;  addr_rom[ 1780]='h00001bd0;  wr_data_rom[ 1780]='h00001360;
    rd_cycle[ 1781] = 1'b0;  wr_cycle[ 1781] = 1'b1;  addr_rom[ 1781]='h00001bd4;  wr_data_rom[ 1781]='h000022e5;
    rd_cycle[ 1782] = 1'b0;  wr_cycle[ 1782] = 1'b1;  addr_rom[ 1782]='h00001bd8;  wr_data_rom[ 1782]='h000014ee;
    rd_cycle[ 1783] = 1'b0;  wr_cycle[ 1783] = 1'b1;  addr_rom[ 1783]='h00001bdc;  wr_data_rom[ 1783]='h00002eb1;
    rd_cycle[ 1784] = 1'b0;  wr_cycle[ 1784] = 1'b1;  addr_rom[ 1784]='h00001be0;  wr_data_rom[ 1784]='h0000365a;
    rd_cycle[ 1785] = 1'b0;  wr_cycle[ 1785] = 1'b1;  addr_rom[ 1785]='h00001be4;  wr_data_rom[ 1785]='h00000834;
    rd_cycle[ 1786] = 1'b0;  wr_cycle[ 1786] = 1'b1;  addr_rom[ 1786]='h00001be8;  wr_data_rom[ 1786]='h000019f1;
    rd_cycle[ 1787] = 1'b0;  wr_cycle[ 1787] = 1'b1;  addr_rom[ 1787]='h00001bec;  wr_data_rom[ 1787]='h00003e87;
    rd_cycle[ 1788] = 1'b0;  wr_cycle[ 1788] = 1'b1;  addr_rom[ 1788]='h00001bf0;  wr_data_rom[ 1788]='h00002fc2;
    rd_cycle[ 1789] = 1'b0;  wr_cycle[ 1789] = 1'b1;  addr_rom[ 1789]='h00001bf4;  wr_data_rom[ 1789]='h00003e94;
    rd_cycle[ 1790] = 1'b0;  wr_cycle[ 1790] = 1'b1;  addr_rom[ 1790]='h00001bf8;  wr_data_rom[ 1790]='h00002ab8;
    rd_cycle[ 1791] = 1'b0;  wr_cycle[ 1791] = 1'b1;  addr_rom[ 1791]='h00001bfc;  wr_data_rom[ 1791]='h00000dae;
    rd_cycle[ 1792] = 1'b0;  wr_cycle[ 1792] = 1'b1;  addr_rom[ 1792]='h00001c00;  wr_data_rom[ 1792]='h0000308c;
    rd_cycle[ 1793] = 1'b0;  wr_cycle[ 1793] = 1'b1;  addr_rom[ 1793]='h00001c04;  wr_data_rom[ 1793]='h00001183;
    rd_cycle[ 1794] = 1'b0;  wr_cycle[ 1794] = 1'b1;  addr_rom[ 1794]='h00001c08;  wr_data_rom[ 1794]='h00003fcf;
    rd_cycle[ 1795] = 1'b0;  wr_cycle[ 1795] = 1'b1;  addr_rom[ 1795]='h00001c0c;  wr_data_rom[ 1795]='h00003aed;
    rd_cycle[ 1796] = 1'b0;  wr_cycle[ 1796] = 1'b1;  addr_rom[ 1796]='h00001c10;  wr_data_rom[ 1796]='h0000063e;
    rd_cycle[ 1797] = 1'b0;  wr_cycle[ 1797] = 1'b1;  addr_rom[ 1797]='h00001c14;  wr_data_rom[ 1797]='h00000001;
    rd_cycle[ 1798] = 1'b0;  wr_cycle[ 1798] = 1'b1;  addr_rom[ 1798]='h00001c18;  wr_data_rom[ 1798]='h00000bb7;
    rd_cycle[ 1799] = 1'b0;  wr_cycle[ 1799] = 1'b1;  addr_rom[ 1799]='h00001c1c;  wr_data_rom[ 1799]='h00000af9;
    rd_cycle[ 1800] = 1'b0;  wr_cycle[ 1800] = 1'b1;  addr_rom[ 1800]='h00001c20;  wr_data_rom[ 1800]='h00003d7b;
    rd_cycle[ 1801] = 1'b0;  wr_cycle[ 1801] = 1'b1;  addr_rom[ 1801]='h00001c24;  wr_data_rom[ 1801]='h0000210c;
    rd_cycle[ 1802] = 1'b0;  wr_cycle[ 1802] = 1'b1;  addr_rom[ 1802]='h00001c28;  wr_data_rom[ 1802]='h00002c4e;
    rd_cycle[ 1803] = 1'b0;  wr_cycle[ 1803] = 1'b1;  addr_rom[ 1803]='h00001c2c;  wr_data_rom[ 1803]='h00002b3e;
    rd_cycle[ 1804] = 1'b0;  wr_cycle[ 1804] = 1'b1;  addr_rom[ 1804]='h00001c30;  wr_data_rom[ 1804]='h00002929;
    rd_cycle[ 1805] = 1'b0;  wr_cycle[ 1805] = 1'b1;  addr_rom[ 1805]='h00001c34;  wr_data_rom[ 1805]='h00002bcb;
    rd_cycle[ 1806] = 1'b0;  wr_cycle[ 1806] = 1'b1;  addr_rom[ 1806]='h00001c38;  wr_data_rom[ 1806]='h0000156b;
    rd_cycle[ 1807] = 1'b0;  wr_cycle[ 1807] = 1'b1;  addr_rom[ 1807]='h00001c3c;  wr_data_rom[ 1807]='h000015e1;
    rd_cycle[ 1808] = 1'b0;  wr_cycle[ 1808] = 1'b1;  addr_rom[ 1808]='h00001c40;  wr_data_rom[ 1808]='h00002395;
    rd_cycle[ 1809] = 1'b0;  wr_cycle[ 1809] = 1'b1;  addr_rom[ 1809]='h00001c44;  wr_data_rom[ 1809]='h00003c5a;
    rd_cycle[ 1810] = 1'b0;  wr_cycle[ 1810] = 1'b1;  addr_rom[ 1810]='h00001c48;  wr_data_rom[ 1810]='h00003233;
    rd_cycle[ 1811] = 1'b0;  wr_cycle[ 1811] = 1'b1;  addr_rom[ 1811]='h00001c4c;  wr_data_rom[ 1811]='h00002cf4;
    rd_cycle[ 1812] = 1'b0;  wr_cycle[ 1812] = 1'b1;  addr_rom[ 1812]='h00001c50;  wr_data_rom[ 1812]='h00002130;
    rd_cycle[ 1813] = 1'b0;  wr_cycle[ 1813] = 1'b1;  addr_rom[ 1813]='h00001c54;  wr_data_rom[ 1813]='h00002fae;
    rd_cycle[ 1814] = 1'b0;  wr_cycle[ 1814] = 1'b1;  addr_rom[ 1814]='h00001c58;  wr_data_rom[ 1814]='h0000034e;
    rd_cycle[ 1815] = 1'b0;  wr_cycle[ 1815] = 1'b1;  addr_rom[ 1815]='h00001c5c;  wr_data_rom[ 1815]='h00002047;
    rd_cycle[ 1816] = 1'b0;  wr_cycle[ 1816] = 1'b1;  addr_rom[ 1816]='h00001c60;  wr_data_rom[ 1816]='h000001af;
    rd_cycle[ 1817] = 1'b0;  wr_cycle[ 1817] = 1'b1;  addr_rom[ 1817]='h00001c64;  wr_data_rom[ 1817]='h000028ad;
    rd_cycle[ 1818] = 1'b0;  wr_cycle[ 1818] = 1'b1;  addr_rom[ 1818]='h00001c68;  wr_data_rom[ 1818]='h00003616;
    rd_cycle[ 1819] = 1'b0;  wr_cycle[ 1819] = 1'b1;  addr_rom[ 1819]='h00001c6c;  wr_data_rom[ 1819]='h00002c70;
    rd_cycle[ 1820] = 1'b0;  wr_cycle[ 1820] = 1'b1;  addr_rom[ 1820]='h00001c70;  wr_data_rom[ 1820]='h00000532;
    rd_cycle[ 1821] = 1'b0;  wr_cycle[ 1821] = 1'b1;  addr_rom[ 1821]='h00001c74;  wr_data_rom[ 1821]='h000035f8;
    rd_cycle[ 1822] = 1'b0;  wr_cycle[ 1822] = 1'b1;  addr_rom[ 1822]='h00001c78;  wr_data_rom[ 1822]='h00001088;
    rd_cycle[ 1823] = 1'b0;  wr_cycle[ 1823] = 1'b1;  addr_rom[ 1823]='h00001c7c;  wr_data_rom[ 1823]='h000036d9;
    rd_cycle[ 1824] = 1'b0;  wr_cycle[ 1824] = 1'b1;  addr_rom[ 1824]='h00001c80;  wr_data_rom[ 1824]='h00000227;
    rd_cycle[ 1825] = 1'b0;  wr_cycle[ 1825] = 1'b1;  addr_rom[ 1825]='h00001c84;  wr_data_rom[ 1825]='h00003b3d;
    rd_cycle[ 1826] = 1'b0;  wr_cycle[ 1826] = 1'b1;  addr_rom[ 1826]='h00001c88;  wr_data_rom[ 1826]='h000022ef;
    rd_cycle[ 1827] = 1'b0;  wr_cycle[ 1827] = 1'b1;  addr_rom[ 1827]='h00001c8c;  wr_data_rom[ 1827]='h00003ca4;
    rd_cycle[ 1828] = 1'b0;  wr_cycle[ 1828] = 1'b1;  addr_rom[ 1828]='h00001c90;  wr_data_rom[ 1828]='h000019d5;
    rd_cycle[ 1829] = 1'b0;  wr_cycle[ 1829] = 1'b1;  addr_rom[ 1829]='h00001c94;  wr_data_rom[ 1829]='h00003f61;
    rd_cycle[ 1830] = 1'b0;  wr_cycle[ 1830] = 1'b1;  addr_rom[ 1830]='h00001c98;  wr_data_rom[ 1830]='h00001a8b;
    rd_cycle[ 1831] = 1'b0;  wr_cycle[ 1831] = 1'b1;  addr_rom[ 1831]='h00001c9c;  wr_data_rom[ 1831]='h00001985;
    rd_cycle[ 1832] = 1'b0;  wr_cycle[ 1832] = 1'b1;  addr_rom[ 1832]='h00001ca0;  wr_data_rom[ 1832]='h00003f16;
    rd_cycle[ 1833] = 1'b0;  wr_cycle[ 1833] = 1'b1;  addr_rom[ 1833]='h00001ca4;  wr_data_rom[ 1833]='h00002def;
    rd_cycle[ 1834] = 1'b0;  wr_cycle[ 1834] = 1'b1;  addr_rom[ 1834]='h00001ca8;  wr_data_rom[ 1834]='h00001812;
    rd_cycle[ 1835] = 1'b0;  wr_cycle[ 1835] = 1'b1;  addr_rom[ 1835]='h00001cac;  wr_data_rom[ 1835]='h00000205;
    rd_cycle[ 1836] = 1'b0;  wr_cycle[ 1836] = 1'b1;  addr_rom[ 1836]='h00001cb0;  wr_data_rom[ 1836]='h00001fc1;
    rd_cycle[ 1837] = 1'b0;  wr_cycle[ 1837] = 1'b1;  addr_rom[ 1837]='h00001cb4;  wr_data_rom[ 1837]='h00002a35;
    rd_cycle[ 1838] = 1'b0;  wr_cycle[ 1838] = 1'b1;  addr_rom[ 1838]='h00001cb8;  wr_data_rom[ 1838]='h000014b2;
    rd_cycle[ 1839] = 1'b0;  wr_cycle[ 1839] = 1'b1;  addr_rom[ 1839]='h00001cbc;  wr_data_rom[ 1839]='h00001704;
    rd_cycle[ 1840] = 1'b0;  wr_cycle[ 1840] = 1'b1;  addr_rom[ 1840]='h00001cc0;  wr_data_rom[ 1840]='h000018f4;
    rd_cycle[ 1841] = 1'b0;  wr_cycle[ 1841] = 1'b1;  addr_rom[ 1841]='h00001cc4;  wr_data_rom[ 1841]='h00003e3c;
    rd_cycle[ 1842] = 1'b0;  wr_cycle[ 1842] = 1'b1;  addr_rom[ 1842]='h00001cc8;  wr_data_rom[ 1842]='h00002d9b;
    rd_cycle[ 1843] = 1'b0;  wr_cycle[ 1843] = 1'b1;  addr_rom[ 1843]='h00001ccc;  wr_data_rom[ 1843]='h00001c87;
    rd_cycle[ 1844] = 1'b0;  wr_cycle[ 1844] = 1'b1;  addr_rom[ 1844]='h00001cd0;  wr_data_rom[ 1844]='h00000810;
    rd_cycle[ 1845] = 1'b0;  wr_cycle[ 1845] = 1'b1;  addr_rom[ 1845]='h00001cd4;  wr_data_rom[ 1845]='h00000e2f;
    rd_cycle[ 1846] = 1'b0;  wr_cycle[ 1846] = 1'b1;  addr_rom[ 1846]='h00001cd8;  wr_data_rom[ 1846]='h000034a1;
    rd_cycle[ 1847] = 1'b0;  wr_cycle[ 1847] = 1'b1;  addr_rom[ 1847]='h00001cdc;  wr_data_rom[ 1847]='h00003c5c;
    rd_cycle[ 1848] = 1'b0;  wr_cycle[ 1848] = 1'b1;  addr_rom[ 1848]='h00001ce0;  wr_data_rom[ 1848]='h00001851;
    rd_cycle[ 1849] = 1'b0;  wr_cycle[ 1849] = 1'b1;  addr_rom[ 1849]='h00001ce4;  wr_data_rom[ 1849]='h0000053b;
    rd_cycle[ 1850] = 1'b0;  wr_cycle[ 1850] = 1'b1;  addr_rom[ 1850]='h00001ce8;  wr_data_rom[ 1850]='h00001496;
    rd_cycle[ 1851] = 1'b0;  wr_cycle[ 1851] = 1'b1;  addr_rom[ 1851]='h00001cec;  wr_data_rom[ 1851]='h0000059c;
    rd_cycle[ 1852] = 1'b0;  wr_cycle[ 1852] = 1'b1;  addr_rom[ 1852]='h00001cf0;  wr_data_rom[ 1852]='h00000d0d;
    rd_cycle[ 1853] = 1'b0;  wr_cycle[ 1853] = 1'b1;  addr_rom[ 1853]='h00001cf4;  wr_data_rom[ 1853]='h00001114;
    rd_cycle[ 1854] = 1'b0;  wr_cycle[ 1854] = 1'b1;  addr_rom[ 1854]='h00001cf8;  wr_data_rom[ 1854]='h00001b70;
    rd_cycle[ 1855] = 1'b0;  wr_cycle[ 1855] = 1'b1;  addr_rom[ 1855]='h00001cfc;  wr_data_rom[ 1855]='h00001806;
    rd_cycle[ 1856] = 1'b0;  wr_cycle[ 1856] = 1'b1;  addr_rom[ 1856]='h00001d00;  wr_data_rom[ 1856]='h00000956;
    rd_cycle[ 1857] = 1'b0;  wr_cycle[ 1857] = 1'b1;  addr_rom[ 1857]='h00001d04;  wr_data_rom[ 1857]='h00003488;
    rd_cycle[ 1858] = 1'b0;  wr_cycle[ 1858] = 1'b1;  addr_rom[ 1858]='h00001d08;  wr_data_rom[ 1858]='h00002e64;
    rd_cycle[ 1859] = 1'b0;  wr_cycle[ 1859] = 1'b1;  addr_rom[ 1859]='h00001d0c;  wr_data_rom[ 1859]='h00003fc1;
    rd_cycle[ 1860] = 1'b0;  wr_cycle[ 1860] = 1'b1;  addr_rom[ 1860]='h00001d10;  wr_data_rom[ 1860]='h00002616;
    rd_cycle[ 1861] = 1'b0;  wr_cycle[ 1861] = 1'b1;  addr_rom[ 1861]='h00001d14;  wr_data_rom[ 1861]='h000038de;
    rd_cycle[ 1862] = 1'b0;  wr_cycle[ 1862] = 1'b1;  addr_rom[ 1862]='h00001d18;  wr_data_rom[ 1862]='h00000bf8;
    rd_cycle[ 1863] = 1'b0;  wr_cycle[ 1863] = 1'b1;  addr_rom[ 1863]='h00001d1c;  wr_data_rom[ 1863]='h000013c0;
    rd_cycle[ 1864] = 1'b0;  wr_cycle[ 1864] = 1'b1;  addr_rom[ 1864]='h00001d20;  wr_data_rom[ 1864]='h0000117d;
    rd_cycle[ 1865] = 1'b0;  wr_cycle[ 1865] = 1'b1;  addr_rom[ 1865]='h00001d24;  wr_data_rom[ 1865]='h00000f71;
    rd_cycle[ 1866] = 1'b0;  wr_cycle[ 1866] = 1'b1;  addr_rom[ 1866]='h00001d28;  wr_data_rom[ 1866]='h00003a9e;
    rd_cycle[ 1867] = 1'b0;  wr_cycle[ 1867] = 1'b1;  addr_rom[ 1867]='h00001d2c;  wr_data_rom[ 1867]='h0000356a;
    rd_cycle[ 1868] = 1'b0;  wr_cycle[ 1868] = 1'b1;  addr_rom[ 1868]='h00001d30;  wr_data_rom[ 1868]='h00001464;
    rd_cycle[ 1869] = 1'b0;  wr_cycle[ 1869] = 1'b1;  addr_rom[ 1869]='h00001d34;  wr_data_rom[ 1869]='h00002054;
    rd_cycle[ 1870] = 1'b0;  wr_cycle[ 1870] = 1'b1;  addr_rom[ 1870]='h00001d38;  wr_data_rom[ 1870]='h00003e41;
    rd_cycle[ 1871] = 1'b0;  wr_cycle[ 1871] = 1'b1;  addr_rom[ 1871]='h00001d3c;  wr_data_rom[ 1871]='h00003703;
    rd_cycle[ 1872] = 1'b0;  wr_cycle[ 1872] = 1'b1;  addr_rom[ 1872]='h00001d40;  wr_data_rom[ 1872]='h00000066;
    rd_cycle[ 1873] = 1'b0;  wr_cycle[ 1873] = 1'b1;  addr_rom[ 1873]='h00001d44;  wr_data_rom[ 1873]='h00000e27;
    rd_cycle[ 1874] = 1'b0;  wr_cycle[ 1874] = 1'b1;  addr_rom[ 1874]='h00001d48;  wr_data_rom[ 1874]='h00000220;
    rd_cycle[ 1875] = 1'b0;  wr_cycle[ 1875] = 1'b1;  addr_rom[ 1875]='h00001d4c;  wr_data_rom[ 1875]='h00003f93;
    rd_cycle[ 1876] = 1'b0;  wr_cycle[ 1876] = 1'b1;  addr_rom[ 1876]='h00001d50;  wr_data_rom[ 1876]='h00000037;
    rd_cycle[ 1877] = 1'b0;  wr_cycle[ 1877] = 1'b1;  addr_rom[ 1877]='h00001d54;  wr_data_rom[ 1877]='h00000b11;
    rd_cycle[ 1878] = 1'b0;  wr_cycle[ 1878] = 1'b1;  addr_rom[ 1878]='h00001d58;  wr_data_rom[ 1878]='h00000eb7;
    rd_cycle[ 1879] = 1'b0;  wr_cycle[ 1879] = 1'b1;  addr_rom[ 1879]='h00001d5c;  wr_data_rom[ 1879]='h0000100f;
    rd_cycle[ 1880] = 1'b0;  wr_cycle[ 1880] = 1'b1;  addr_rom[ 1880]='h00001d60;  wr_data_rom[ 1880]='h000006cf;
    rd_cycle[ 1881] = 1'b0;  wr_cycle[ 1881] = 1'b1;  addr_rom[ 1881]='h00001d64;  wr_data_rom[ 1881]='h0000139c;
    rd_cycle[ 1882] = 1'b0;  wr_cycle[ 1882] = 1'b1;  addr_rom[ 1882]='h00001d68;  wr_data_rom[ 1882]='h00003eae;
    rd_cycle[ 1883] = 1'b0;  wr_cycle[ 1883] = 1'b1;  addr_rom[ 1883]='h00001d6c;  wr_data_rom[ 1883]='h00000e40;
    rd_cycle[ 1884] = 1'b0;  wr_cycle[ 1884] = 1'b1;  addr_rom[ 1884]='h00001d70;  wr_data_rom[ 1884]='h00002f6c;
    rd_cycle[ 1885] = 1'b0;  wr_cycle[ 1885] = 1'b1;  addr_rom[ 1885]='h00001d74;  wr_data_rom[ 1885]='h00002c22;
    rd_cycle[ 1886] = 1'b0;  wr_cycle[ 1886] = 1'b1;  addr_rom[ 1886]='h00001d78;  wr_data_rom[ 1886]='h00002955;
    rd_cycle[ 1887] = 1'b0;  wr_cycle[ 1887] = 1'b1;  addr_rom[ 1887]='h00001d7c;  wr_data_rom[ 1887]='h0000208c;
    rd_cycle[ 1888] = 1'b0;  wr_cycle[ 1888] = 1'b1;  addr_rom[ 1888]='h00001d80;  wr_data_rom[ 1888]='h00000767;
    rd_cycle[ 1889] = 1'b0;  wr_cycle[ 1889] = 1'b1;  addr_rom[ 1889]='h00001d84;  wr_data_rom[ 1889]='h000020f9;
    rd_cycle[ 1890] = 1'b0;  wr_cycle[ 1890] = 1'b1;  addr_rom[ 1890]='h00001d88;  wr_data_rom[ 1890]='h000035e5;
    rd_cycle[ 1891] = 1'b0;  wr_cycle[ 1891] = 1'b1;  addr_rom[ 1891]='h00001d8c;  wr_data_rom[ 1891]='h00002166;
    rd_cycle[ 1892] = 1'b0;  wr_cycle[ 1892] = 1'b1;  addr_rom[ 1892]='h00001d90;  wr_data_rom[ 1892]='h00000292;
    rd_cycle[ 1893] = 1'b0;  wr_cycle[ 1893] = 1'b1;  addr_rom[ 1893]='h00001d94;  wr_data_rom[ 1893]='h0000348c;
    rd_cycle[ 1894] = 1'b0;  wr_cycle[ 1894] = 1'b1;  addr_rom[ 1894]='h00001d98;  wr_data_rom[ 1894]='h00000ec9;
    rd_cycle[ 1895] = 1'b0;  wr_cycle[ 1895] = 1'b1;  addr_rom[ 1895]='h00001d9c;  wr_data_rom[ 1895]='h000019ff;
    rd_cycle[ 1896] = 1'b0;  wr_cycle[ 1896] = 1'b1;  addr_rom[ 1896]='h00001da0;  wr_data_rom[ 1896]='h00003e11;
    rd_cycle[ 1897] = 1'b0;  wr_cycle[ 1897] = 1'b1;  addr_rom[ 1897]='h00001da4;  wr_data_rom[ 1897]='h000028c2;
    rd_cycle[ 1898] = 1'b0;  wr_cycle[ 1898] = 1'b1;  addr_rom[ 1898]='h00001da8;  wr_data_rom[ 1898]='h00002051;
    rd_cycle[ 1899] = 1'b0;  wr_cycle[ 1899] = 1'b1;  addr_rom[ 1899]='h00001dac;  wr_data_rom[ 1899]='h00000824;
    rd_cycle[ 1900] = 1'b0;  wr_cycle[ 1900] = 1'b1;  addr_rom[ 1900]='h00001db0;  wr_data_rom[ 1900]='h0000126e;
    rd_cycle[ 1901] = 1'b0;  wr_cycle[ 1901] = 1'b1;  addr_rom[ 1901]='h00001db4;  wr_data_rom[ 1901]='h00003051;
    rd_cycle[ 1902] = 1'b0;  wr_cycle[ 1902] = 1'b1;  addr_rom[ 1902]='h00001db8;  wr_data_rom[ 1902]='h0000349b;
    rd_cycle[ 1903] = 1'b0;  wr_cycle[ 1903] = 1'b1;  addr_rom[ 1903]='h00001dbc;  wr_data_rom[ 1903]='h000002f3;
    rd_cycle[ 1904] = 1'b0;  wr_cycle[ 1904] = 1'b1;  addr_rom[ 1904]='h00001dc0;  wr_data_rom[ 1904]='h000012d2;
    rd_cycle[ 1905] = 1'b0;  wr_cycle[ 1905] = 1'b1;  addr_rom[ 1905]='h00001dc4;  wr_data_rom[ 1905]='h00002656;
    rd_cycle[ 1906] = 1'b0;  wr_cycle[ 1906] = 1'b1;  addr_rom[ 1906]='h00001dc8;  wr_data_rom[ 1906]='h00002616;
    rd_cycle[ 1907] = 1'b0;  wr_cycle[ 1907] = 1'b1;  addr_rom[ 1907]='h00001dcc;  wr_data_rom[ 1907]='h00003b4c;
    rd_cycle[ 1908] = 1'b0;  wr_cycle[ 1908] = 1'b1;  addr_rom[ 1908]='h00001dd0;  wr_data_rom[ 1908]='h00000149;
    rd_cycle[ 1909] = 1'b0;  wr_cycle[ 1909] = 1'b1;  addr_rom[ 1909]='h00001dd4;  wr_data_rom[ 1909]='h0000304a;
    rd_cycle[ 1910] = 1'b0;  wr_cycle[ 1910] = 1'b1;  addr_rom[ 1910]='h00001dd8;  wr_data_rom[ 1910]='h0000381a;
    rd_cycle[ 1911] = 1'b0;  wr_cycle[ 1911] = 1'b1;  addr_rom[ 1911]='h00001ddc;  wr_data_rom[ 1911]='h00000d00;
    rd_cycle[ 1912] = 1'b0;  wr_cycle[ 1912] = 1'b1;  addr_rom[ 1912]='h00001de0;  wr_data_rom[ 1912]='h0000098b;
    rd_cycle[ 1913] = 1'b0;  wr_cycle[ 1913] = 1'b1;  addr_rom[ 1913]='h00001de4;  wr_data_rom[ 1913]='h000026a7;
    rd_cycle[ 1914] = 1'b0;  wr_cycle[ 1914] = 1'b1;  addr_rom[ 1914]='h00001de8;  wr_data_rom[ 1914]='h00001c2a;
    rd_cycle[ 1915] = 1'b0;  wr_cycle[ 1915] = 1'b1;  addr_rom[ 1915]='h00001dec;  wr_data_rom[ 1915]='h00001dc7;
    rd_cycle[ 1916] = 1'b0;  wr_cycle[ 1916] = 1'b1;  addr_rom[ 1916]='h00001df0;  wr_data_rom[ 1916]='h00001625;
    rd_cycle[ 1917] = 1'b0;  wr_cycle[ 1917] = 1'b1;  addr_rom[ 1917]='h00001df4;  wr_data_rom[ 1917]='h00000e2a;
    rd_cycle[ 1918] = 1'b0;  wr_cycle[ 1918] = 1'b1;  addr_rom[ 1918]='h00001df8;  wr_data_rom[ 1918]='h00000841;
    rd_cycle[ 1919] = 1'b0;  wr_cycle[ 1919] = 1'b1;  addr_rom[ 1919]='h00001dfc;  wr_data_rom[ 1919]='h0000032e;
    rd_cycle[ 1920] = 1'b0;  wr_cycle[ 1920] = 1'b1;  addr_rom[ 1920]='h00001e00;  wr_data_rom[ 1920]='h000023bf;
    rd_cycle[ 1921] = 1'b0;  wr_cycle[ 1921] = 1'b1;  addr_rom[ 1921]='h00001e04;  wr_data_rom[ 1921]='h000036e3;
    rd_cycle[ 1922] = 1'b0;  wr_cycle[ 1922] = 1'b1;  addr_rom[ 1922]='h00001e08;  wr_data_rom[ 1922]='h00000791;
    rd_cycle[ 1923] = 1'b0;  wr_cycle[ 1923] = 1'b1;  addr_rom[ 1923]='h00001e0c;  wr_data_rom[ 1923]='h00000327;
    rd_cycle[ 1924] = 1'b0;  wr_cycle[ 1924] = 1'b1;  addr_rom[ 1924]='h00001e10;  wr_data_rom[ 1924]='h00002d65;
    rd_cycle[ 1925] = 1'b0;  wr_cycle[ 1925] = 1'b1;  addr_rom[ 1925]='h00001e14;  wr_data_rom[ 1925]='h000008bd;
    rd_cycle[ 1926] = 1'b0;  wr_cycle[ 1926] = 1'b1;  addr_rom[ 1926]='h00001e18;  wr_data_rom[ 1926]='h00002eae;
    rd_cycle[ 1927] = 1'b0;  wr_cycle[ 1927] = 1'b1;  addr_rom[ 1927]='h00001e1c;  wr_data_rom[ 1927]='h00001cde;
    rd_cycle[ 1928] = 1'b0;  wr_cycle[ 1928] = 1'b1;  addr_rom[ 1928]='h00001e20;  wr_data_rom[ 1928]='h000018fc;
    rd_cycle[ 1929] = 1'b0;  wr_cycle[ 1929] = 1'b1;  addr_rom[ 1929]='h00001e24;  wr_data_rom[ 1929]='h00003f0b;
    rd_cycle[ 1930] = 1'b0;  wr_cycle[ 1930] = 1'b1;  addr_rom[ 1930]='h00001e28;  wr_data_rom[ 1930]='h000021ef;
    rd_cycle[ 1931] = 1'b0;  wr_cycle[ 1931] = 1'b1;  addr_rom[ 1931]='h00001e2c;  wr_data_rom[ 1931]='h0000315a;
    rd_cycle[ 1932] = 1'b0;  wr_cycle[ 1932] = 1'b1;  addr_rom[ 1932]='h00001e30;  wr_data_rom[ 1932]='h00000d37;
    rd_cycle[ 1933] = 1'b0;  wr_cycle[ 1933] = 1'b1;  addr_rom[ 1933]='h00001e34;  wr_data_rom[ 1933]='h00000468;
    rd_cycle[ 1934] = 1'b0;  wr_cycle[ 1934] = 1'b1;  addr_rom[ 1934]='h00001e38;  wr_data_rom[ 1934]='h000036c2;
    rd_cycle[ 1935] = 1'b0;  wr_cycle[ 1935] = 1'b1;  addr_rom[ 1935]='h00001e3c;  wr_data_rom[ 1935]='h00000044;
    rd_cycle[ 1936] = 1'b0;  wr_cycle[ 1936] = 1'b1;  addr_rom[ 1936]='h00001e40;  wr_data_rom[ 1936]='h00001157;
    rd_cycle[ 1937] = 1'b0;  wr_cycle[ 1937] = 1'b1;  addr_rom[ 1937]='h00001e44;  wr_data_rom[ 1937]='h00003452;
    rd_cycle[ 1938] = 1'b0;  wr_cycle[ 1938] = 1'b1;  addr_rom[ 1938]='h00001e48;  wr_data_rom[ 1938]='h00003f8e;
    rd_cycle[ 1939] = 1'b0;  wr_cycle[ 1939] = 1'b1;  addr_rom[ 1939]='h00001e4c;  wr_data_rom[ 1939]='h000018f4;
    rd_cycle[ 1940] = 1'b0;  wr_cycle[ 1940] = 1'b1;  addr_rom[ 1940]='h00001e50;  wr_data_rom[ 1940]='h00003433;
    rd_cycle[ 1941] = 1'b0;  wr_cycle[ 1941] = 1'b1;  addr_rom[ 1941]='h00001e54;  wr_data_rom[ 1941]='h00003507;
    rd_cycle[ 1942] = 1'b0;  wr_cycle[ 1942] = 1'b1;  addr_rom[ 1942]='h00001e58;  wr_data_rom[ 1942]='h00000658;
    rd_cycle[ 1943] = 1'b0;  wr_cycle[ 1943] = 1'b1;  addr_rom[ 1943]='h00001e5c;  wr_data_rom[ 1943]='h0000235a;
    rd_cycle[ 1944] = 1'b0;  wr_cycle[ 1944] = 1'b1;  addr_rom[ 1944]='h00001e60;  wr_data_rom[ 1944]='h00003f42;
    rd_cycle[ 1945] = 1'b0;  wr_cycle[ 1945] = 1'b1;  addr_rom[ 1945]='h00001e64;  wr_data_rom[ 1945]='h00002d32;
    rd_cycle[ 1946] = 1'b0;  wr_cycle[ 1946] = 1'b1;  addr_rom[ 1946]='h00001e68;  wr_data_rom[ 1946]='h0000305c;
    rd_cycle[ 1947] = 1'b0;  wr_cycle[ 1947] = 1'b1;  addr_rom[ 1947]='h00001e6c;  wr_data_rom[ 1947]='h00003a81;
    rd_cycle[ 1948] = 1'b0;  wr_cycle[ 1948] = 1'b1;  addr_rom[ 1948]='h00001e70;  wr_data_rom[ 1948]='h00001d4e;
    rd_cycle[ 1949] = 1'b0;  wr_cycle[ 1949] = 1'b1;  addr_rom[ 1949]='h00001e74;  wr_data_rom[ 1949]='h000033c7;
    rd_cycle[ 1950] = 1'b0;  wr_cycle[ 1950] = 1'b1;  addr_rom[ 1950]='h00001e78;  wr_data_rom[ 1950]='h00000ec0;
    rd_cycle[ 1951] = 1'b0;  wr_cycle[ 1951] = 1'b1;  addr_rom[ 1951]='h00001e7c;  wr_data_rom[ 1951]='h0000241f;
    rd_cycle[ 1952] = 1'b0;  wr_cycle[ 1952] = 1'b1;  addr_rom[ 1952]='h00001e80;  wr_data_rom[ 1952]='h00003c03;
    rd_cycle[ 1953] = 1'b0;  wr_cycle[ 1953] = 1'b1;  addr_rom[ 1953]='h00001e84;  wr_data_rom[ 1953]='h000008f1;
    rd_cycle[ 1954] = 1'b0;  wr_cycle[ 1954] = 1'b1;  addr_rom[ 1954]='h00001e88;  wr_data_rom[ 1954]='h000016e3;
    rd_cycle[ 1955] = 1'b0;  wr_cycle[ 1955] = 1'b1;  addr_rom[ 1955]='h00001e8c;  wr_data_rom[ 1955]='h0000283b;
    rd_cycle[ 1956] = 1'b0;  wr_cycle[ 1956] = 1'b1;  addr_rom[ 1956]='h00001e90;  wr_data_rom[ 1956]='h000021b4;
    rd_cycle[ 1957] = 1'b0;  wr_cycle[ 1957] = 1'b1;  addr_rom[ 1957]='h00001e94;  wr_data_rom[ 1957]='h0000388e;
    rd_cycle[ 1958] = 1'b0;  wr_cycle[ 1958] = 1'b1;  addr_rom[ 1958]='h00001e98;  wr_data_rom[ 1958]='h00001848;
    rd_cycle[ 1959] = 1'b0;  wr_cycle[ 1959] = 1'b1;  addr_rom[ 1959]='h00001e9c;  wr_data_rom[ 1959]='h00000bb9;
    rd_cycle[ 1960] = 1'b0;  wr_cycle[ 1960] = 1'b1;  addr_rom[ 1960]='h00001ea0;  wr_data_rom[ 1960]='h000002dd;
    rd_cycle[ 1961] = 1'b0;  wr_cycle[ 1961] = 1'b1;  addr_rom[ 1961]='h00001ea4;  wr_data_rom[ 1961]='h00003f51;
    rd_cycle[ 1962] = 1'b0;  wr_cycle[ 1962] = 1'b1;  addr_rom[ 1962]='h00001ea8;  wr_data_rom[ 1962]='h00001b97;
    rd_cycle[ 1963] = 1'b0;  wr_cycle[ 1963] = 1'b1;  addr_rom[ 1963]='h00001eac;  wr_data_rom[ 1963]='h00000e0e;
    rd_cycle[ 1964] = 1'b0;  wr_cycle[ 1964] = 1'b1;  addr_rom[ 1964]='h00001eb0;  wr_data_rom[ 1964]='h000006ba;
    rd_cycle[ 1965] = 1'b0;  wr_cycle[ 1965] = 1'b1;  addr_rom[ 1965]='h00001eb4;  wr_data_rom[ 1965]='h000037da;
    rd_cycle[ 1966] = 1'b0;  wr_cycle[ 1966] = 1'b1;  addr_rom[ 1966]='h00001eb8;  wr_data_rom[ 1966]='h00001c5d;
    rd_cycle[ 1967] = 1'b0;  wr_cycle[ 1967] = 1'b1;  addr_rom[ 1967]='h00001ebc;  wr_data_rom[ 1967]='h000032ab;
    rd_cycle[ 1968] = 1'b0;  wr_cycle[ 1968] = 1'b1;  addr_rom[ 1968]='h00001ec0;  wr_data_rom[ 1968]='h000022ea;
    rd_cycle[ 1969] = 1'b0;  wr_cycle[ 1969] = 1'b1;  addr_rom[ 1969]='h00001ec4;  wr_data_rom[ 1969]='h000016c9;
    rd_cycle[ 1970] = 1'b0;  wr_cycle[ 1970] = 1'b1;  addr_rom[ 1970]='h00001ec8;  wr_data_rom[ 1970]='h00002208;
    rd_cycle[ 1971] = 1'b0;  wr_cycle[ 1971] = 1'b1;  addr_rom[ 1971]='h00001ecc;  wr_data_rom[ 1971]='h0000346d;
    rd_cycle[ 1972] = 1'b0;  wr_cycle[ 1972] = 1'b1;  addr_rom[ 1972]='h00001ed0;  wr_data_rom[ 1972]='h000021d8;
    rd_cycle[ 1973] = 1'b0;  wr_cycle[ 1973] = 1'b1;  addr_rom[ 1973]='h00001ed4;  wr_data_rom[ 1973]='h00001893;
    rd_cycle[ 1974] = 1'b0;  wr_cycle[ 1974] = 1'b1;  addr_rom[ 1974]='h00001ed8;  wr_data_rom[ 1974]='h000038ae;
    rd_cycle[ 1975] = 1'b0;  wr_cycle[ 1975] = 1'b1;  addr_rom[ 1975]='h00001edc;  wr_data_rom[ 1975]='h000005d7;
    rd_cycle[ 1976] = 1'b0;  wr_cycle[ 1976] = 1'b1;  addr_rom[ 1976]='h00001ee0;  wr_data_rom[ 1976]='h0000275a;
    rd_cycle[ 1977] = 1'b0;  wr_cycle[ 1977] = 1'b1;  addr_rom[ 1977]='h00001ee4;  wr_data_rom[ 1977]='h0000359a;
    rd_cycle[ 1978] = 1'b0;  wr_cycle[ 1978] = 1'b1;  addr_rom[ 1978]='h00001ee8;  wr_data_rom[ 1978]='h00002e22;
    rd_cycle[ 1979] = 1'b0;  wr_cycle[ 1979] = 1'b1;  addr_rom[ 1979]='h00001eec;  wr_data_rom[ 1979]='h00003665;
    rd_cycle[ 1980] = 1'b0;  wr_cycle[ 1980] = 1'b1;  addr_rom[ 1980]='h00001ef0;  wr_data_rom[ 1980]='h00001e82;
    rd_cycle[ 1981] = 1'b0;  wr_cycle[ 1981] = 1'b1;  addr_rom[ 1981]='h00001ef4;  wr_data_rom[ 1981]='h000009fb;
    rd_cycle[ 1982] = 1'b0;  wr_cycle[ 1982] = 1'b1;  addr_rom[ 1982]='h00001ef8;  wr_data_rom[ 1982]='h00003b74;
    rd_cycle[ 1983] = 1'b0;  wr_cycle[ 1983] = 1'b1;  addr_rom[ 1983]='h00001efc;  wr_data_rom[ 1983]='h00001ed8;
    rd_cycle[ 1984] = 1'b0;  wr_cycle[ 1984] = 1'b1;  addr_rom[ 1984]='h00001f00;  wr_data_rom[ 1984]='h00002358;
    rd_cycle[ 1985] = 1'b0;  wr_cycle[ 1985] = 1'b1;  addr_rom[ 1985]='h00001f04;  wr_data_rom[ 1985]='h000035d2;
    rd_cycle[ 1986] = 1'b0;  wr_cycle[ 1986] = 1'b1;  addr_rom[ 1986]='h00001f08;  wr_data_rom[ 1986]='h00000a12;
    rd_cycle[ 1987] = 1'b0;  wr_cycle[ 1987] = 1'b1;  addr_rom[ 1987]='h00001f0c;  wr_data_rom[ 1987]='h000020b6;
    rd_cycle[ 1988] = 1'b0;  wr_cycle[ 1988] = 1'b1;  addr_rom[ 1988]='h00001f10;  wr_data_rom[ 1988]='h000007b6;
    rd_cycle[ 1989] = 1'b0;  wr_cycle[ 1989] = 1'b1;  addr_rom[ 1989]='h00001f14;  wr_data_rom[ 1989]='h00002a08;
    rd_cycle[ 1990] = 1'b0;  wr_cycle[ 1990] = 1'b1;  addr_rom[ 1990]='h00001f18;  wr_data_rom[ 1990]='h00003252;
    rd_cycle[ 1991] = 1'b0;  wr_cycle[ 1991] = 1'b1;  addr_rom[ 1991]='h00001f1c;  wr_data_rom[ 1991]='h00003207;
    rd_cycle[ 1992] = 1'b0;  wr_cycle[ 1992] = 1'b1;  addr_rom[ 1992]='h00001f20;  wr_data_rom[ 1992]='h00000fe1;
    rd_cycle[ 1993] = 1'b0;  wr_cycle[ 1993] = 1'b1;  addr_rom[ 1993]='h00001f24;  wr_data_rom[ 1993]='h00002852;
    rd_cycle[ 1994] = 1'b0;  wr_cycle[ 1994] = 1'b1;  addr_rom[ 1994]='h00001f28;  wr_data_rom[ 1994]='h00000d12;
    rd_cycle[ 1995] = 1'b0;  wr_cycle[ 1995] = 1'b1;  addr_rom[ 1995]='h00001f2c;  wr_data_rom[ 1995]='h000011a2;
    rd_cycle[ 1996] = 1'b0;  wr_cycle[ 1996] = 1'b1;  addr_rom[ 1996]='h00001f30;  wr_data_rom[ 1996]='h0000127f;
    rd_cycle[ 1997] = 1'b0;  wr_cycle[ 1997] = 1'b1;  addr_rom[ 1997]='h00001f34;  wr_data_rom[ 1997]='h00000f2f;
    rd_cycle[ 1998] = 1'b0;  wr_cycle[ 1998] = 1'b1;  addr_rom[ 1998]='h00001f38;  wr_data_rom[ 1998]='h00000631;
    rd_cycle[ 1999] = 1'b0;  wr_cycle[ 1999] = 1'b1;  addr_rom[ 1999]='h00001f3c;  wr_data_rom[ 1999]='h00001aac;
    rd_cycle[ 2000] = 1'b0;  wr_cycle[ 2000] = 1'b1;  addr_rom[ 2000]='h00001f40;  wr_data_rom[ 2000]='h00003875;
    rd_cycle[ 2001] = 1'b0;  wr_cycle[ 2001] = 1'b1;  addr_rom[ 2001]='h00001f44;  wr_data_rom[ 2001]='h00002968;
    rd_cycle[ 2002] = 1'b0;  wr_cycle[ 2002] = 1'b1;  addr_rom[ 2002]='h00001f48;  wr_data_rom[ 2002]='h00003e45;
    rd_cycle[ 2003] = 1'b0;  wr_cycle[ 2003] = 1'b1;  addr_rom[ 2003]='h00001f4c;  wr_data_rom[ 2003]='h0000254d;
    rd_cycle[ 2004] = 1'b0;  wr_cycle[ 2004] = 1'b1;  addr_rom[ 2004]='h00001f50;  wr_data_rom[ 2004]='h00000710;
    rd_cycle[ 2005] = 1'b0;  wr_cycle[ 2005] = 1'b1;  addr_rom[ 2005]='h00001f54;  wr_data_rom[ 2005]='h00001fb1;
    rd_cycle[ 2006] = 1'b0;  wr_cycle[ 2006] = 1'b1;  addr_rom[ 2006]='h00001f58;  wr_data_rom[ 2006]='h000029d0;
    rd_cycle[ 2007] = 1'b0;  wr_cycle[ 2007] = 1'b1;  addr_rom[ 2007]='h00001f5c;  wr_data_rom[ 2007]='h00001cc6;
    rd_cycle[ 2008] = 1'b0;  wr_cycle[ 2008] = 1'b1;  addr_rom[ 2008]='h00001f60;  wr_data_rom[ 2008]='h00000168;
    rd_cycle[ 2009] = 1'b0;  wr_cycle[ 2009] = 1'b1;  addr_rom[ 2009]='h00001f64;  wr_data_rom[ 2009]='h00003145;
    rd_cycle[ 2010] = 1'b0;  wr_cycle[ 2010] = 1'b1;  addr_rom[ 2010]='h00001f68;  wr_data_rom[ 2010]='h000017f0;
    rd_cycle[ 2011] = 1'b0;  wr_cycle[ 2011] = 1'b1;  addr_rom[ 2011]='h00001f6c;  wr_data_rom[ 2011]='h00001ea2;
    rd_cycle[ 2012] = 1'b0;  wr_cycle[ 2012] = 1'b1;  addr_rom[ 2012]='h00001f70;  wr_data_rom[ 2012]='h00002fdd;
    rd_cycle[ 2013] = 1'b0;  wr_cycle[ 2013] = 1'b1;  addr_rom[ 2013]='h00001f74;  wr_data_rom[ 2013]='h00003e6b;
    rd_cycle[ 2014] = 1'b0;  wr_cycle[ 2014] = 1'b1;  addr_rom[ 2014]='h00001f78;  wr_data_rom[ 2014]='h000024d8;
    rd_cycle[ 2015] = 1'b0;  wr_cycle[ 2015] = 1'b1;  addr_rom[ 2015]='h00001f7c;  wr_data_rom[ 2015]='h00000aef;
    rd_cycle[ 2016] = 1'b0;  wr_cycle[ 2016] = 1'b1;  addr_rom[ 2016]='h00001f80;  wr_data_rom[ 2016]='h000033a9;
    rd_cycle[ 2017] = 1'b0;  wr_cycle[ 2017] = 1'b1;  addr_rom[ 2017]='h00001f84;  wr_data_rom[ 2017]='h000000ab;
    rd_cycle[ 2018] = 1'b0;  wr_cycle[ 2018] = 1'b1;  addr_rom[ 2018]='h00001f88;  wr_data_rom[ 2018]='h00003cbb;
    rd_cycle[ 2019] = 1'b0;  wr_cycle[ 2019] = 1'b1;  addr_rom[ 2019]='h00001f8c;  wr_data_rom[ 2019]='h00003c1a;
    rd_cycle[ 2020] = 1'b0;  wr_cycle[ 2020] = 1'b1;  addr_rom[ 2020]='h00001f90;  wr_data_rom[ 2020]='h00002511;
    rd_cycle[ 2021] = 1'b0;  wr_cycle[ 2021] = 1'b1;  addr_rom[ 2021]='h00001f94;  wr_data_rom[ 2021]='h00000a6f;
    rd_cycle[ 2022] = 1'b0;  wr_cycle[ 2022] = 1'b1;  addr_rom[ 2022]='h00001f98;  wr_data_rom[ 2022]='h00001c8b;
    rd_cycle[ 2023] = 1'b0;  wr_cycle[ 2023] = 1'b1;  addr_rom[ 2023]='h00001f9c;  wr_data_rom[ 2023]='h00002757;
    rd_cycle[ 2024] = 1'b0;  wr_cycle[ 2024] = 1'b1;  addr_rom[ 2024]='h00001fa0;  wr_data_rom[ 2024]='h0000159f;
    rd_cycle[ 2025] = 1'b0;  wr_cycle[ 2025] = 1'b1;  addr_rom[ 2025]='h00001fa4;  wr_data_rom[ 2025]='h00003754;
    rd_cycle[ 2026] = 1'b0;  wr_cycle[ 2026] = 1'b1;  addr_rom[ 2026]='h00001fa8;  wr_data_rom[ 2026]='h00002cbb;
    rd_cycle[ 2027] = 1'b0;  wr_cycle[ 2027] = 1'b1;  addr_rom[ 2027]='h00001fac;  wr_data_rom[ 2027]='h00003828;
    rd_cycle[ 2028] = 1'b0;  wr_cycle[ 2028] = 1'b1;  addr_rom[ 2028]='h00001fb0;  wr_data_rom[ 2028]='h00001503;
    rd_cycle[ 2029] = 1'b0;  wr_cycle[ 2029] = 1'b1;  addr_rom[ 2029]='h00001fb4;  wr_data_rom[ 2029]='h00002bab;
    rd_cycle[ 2030] = 1'b0;  wr_cycle[ 2030] = 1'b1;  addr_rom[ 2030]='h00001fb8;  wr_data_rom[ 2030]='h00003966;
    rd_cycle[ 2031] = 1'b0;  wr_cycle[ 2031] = 1'b1;  addr_rom[ 2031]='h00001fbc;  wr_data_rom[ 2031]='h00000c1d;
    rd_cycle[ 2032] = 1'b0;  wr_cycle[ 2032] = 1'b1;  addr_rom[ 2032]='h00001fc0;  wr_data_rom[ 2032]='h000027c6;
    rd_cycle[ 2033] = 1'b0;  wr_cycle[ 2033] = 1'b1;  addr_rom[ 2033]='h00001fc4;  wr_data_rom[ 2033]='h00001fae;
    rd_cycle[ 2034] = 1'b0;  wr_cycle[ 2034] = 1'b1;  addr_rom[ 2034]='h00001fc8;  wr_data_rom[ 2034]='h000023aa;
    rd_cycle[ 2035] = 1'b0;  wr_cycle[ 2035] = 1'b1;  addr_rom[ 2035]='h00001fcc;  wr_data_rom[ 2035]='h0000314b;
    rd_cycle[ 2036] = 1'b0;  wr_cycle[ 2036] = 1'b1;  addr_rom[ 2036]='h00001fd0;  wr_data_rom[ 2036]='h0000169f;
    rd_cycle[ 2037] = 1'b0;  wr_cycle[ 2037] = 1'b1;  addr_rom[ 2037]='h00001fd4;  wr_data_rom[ 2037]='h00001683;
    rd_cycle[ 2038] = 1'b0;  wr_cycle[ 2038] = 1'b1;  addr_rom[ 2038]='h00001fd8;  wr_data_rom[ 2038]='h00001a9d;
    rd_cycle[ 2039] = 1'b0;  wr_cycle[ 2039] = 1'b1;  addr_rom[ 2039]='h00001fdc;  wr_data_rom[ 2039]='h00003846;
    rd_cycle[ 2040] = 1'b0;  wr_cycle[ 2040] = 1'b1;  addr_rom[ 2040]='h00001fe0;  wr_data_rom[ 2040]='h000004d1;
    rd_cycle[ 2041] = 1'b0;  wr_cycle[ 2041] = 1'b1;  addr_rom[ 2041]='h00001fe4;  wr_data_rom[ 2041]='h00002b23;
    rd_cycle[ 2042] = 1'b0;  wr_cycle[ 2042] = 1'b1;  addr_rom[ 2042]='h00001fe8;  wr_data_rom[ 2042]='h00003442;
    rd_cycle[ 2043] = 1'b0;  wr_cycle[ 2043] = 1'b1;  addr_rom[ 2043]='h00001fec;  wr_data_rom[ 2043]='h0000323c;
    rd_cycle[ 2044] = 1'b0;  wr_cycle[ 2044] = 1'b1;  addr_rom[ 2044]='h00001ff0;  wr_data_rom[ 2044]='h00000d19;
    rd_cycle[ 2045] = 1'b0;  wr_cycle[ 2045] = 1'b1;  addr_rom[ 2045]='h00001ff4;  wr_data_rom[ 2045]='h0000254c;
    rd_cycle[ 2046] = 1'b0;  wr_cycle[ 2046] = 1'b1;  addr_rom[ 2046]='h00001ff8;  wr_data_rom[ 2046]='h0000175b;
    rd_cycle[ 2047] = 1'b0;  wr_cycle[ 2047] = 1'b1;  addr_rom[ 2047]='h00001ffc;  wr_data_rom[ 2047]='h000004dc;
    rd_cycle[ 2048] = 1'b0;  wr_cycle[ 2048] = 1'b1;  addr_rom[ 2048]='h00002000;  wr_data_rom[ 2048]='h00000461;
    rd_cycle[ 2049] = 1'b0;  wr_cycle[ 2049] = 1'b1;  addr_rom[ 2049]='h00002004;  wr_data_rom[ 2049]='h00000cca;
    rd_cycle[ 2050] = 1'b0;  wr_cycle[ 2050] = 1'b1;  addr_rom[ 2050]='h00002008;  wr_data_rom[ 2050]='h0000093a;
    rd_cycle[ 2051] = 1'b0;  wr_cycle[ 2051] = 1'b1;  addr_rom[ 2051]='h0000200c;  wr_data_rom[ 2051]='h00003afc;
    rd_cycle[ 2052] = 1'b0;  wr_cycle[ 2052] = 1'b1;  addr_rom[ 2052]='h00002010;  wr_data_rom[ 2052]='h00000334;
    rd_cycle[ 2053] = 1'b0;  wr_cycle[ 2053] = 1'b1;  addr_rom[ 2053]='h00002014;  wr_data_rom[ 2053]='h00002114;
    rd_cycle[ 2054] = 1'b0;  wr_cycle[ 2054] = 1'b1;  addr_rom[ 2054]='h00002018;  wr_data_rom[ 2054]='h0000273d;
    rd_cycle[ 2055] = 1'b0;  wr_cycle[ 2055] = 1'b1;  addr_rom[ 2055]='h0000201c;  wr_data_rom[ 2055]='h000024f9;
    rd_cycle[ 2056] = 1'b0;  wr_cycle[ 2056] = 1'b1;  addr_rom[ 2056]='h00002020;  wr_data_rom[ 2056]='h00001a31;
    rd_cycle[ 2057] = 1'b0;  wr_cycle[ 2057] = 1'b1;  addr_rom[ 2057]='h00002024;  wr_data_rom[ 2057]='h000030c9;
    rd_cycle[ 2058] = 1'b0;  wr_cycle[ 2058] = 1'b1;  addr_rom[ 2058]='h00002028;  wr_data_rom[ 2058]='h00001f0e;
    rd_cycle[ 2059] = 1'b0;  wr_cycle[ 2059] = 1'b1;  addr_rom[ 2059]='h0000202c;  wr_data_rom[ 2059]='h0000045d;
    rd_cycle[ 2060] = 1'b0;  wr_cycle[ 2060] = 1'b1;  addr_rom[ 2060]='h00002030;  wr_data_rom[ 2060]='h000007ec;
    rd_cycle[ 2061] = 1'b0;  wr_cycle[ 2061] = 1'b1;  addr_rom[ 2061]='h00002034;  wr_data_rom[ 2061]='h00000211;
    rd_cycle[ 2062] = 1'b0;  wr_cycle[ 2062] = 1'b1;  addr_rom[ 2062]='h00002038;  wr_data_rom[ 2062]='h0000021e;
    rd_cycle[ 2063] = 1'b0;  wr_cycle[ 2063] = 1'b1;  addr_rom[ 2063]='h0000203c;  wr_data_rom[ 2063]='h00000af1;
    rd_cycle[ 2064] = 1'b0;  wr_cycle[ 2064] = 1'b1;  addr_rom[ 2064]='h00002040;  wr_data_rom[ 2064]='h00001b62;
    rd_cycle[ 2065] = 1'b0;  wr_cycle[ 2065] = 1'b1;  addr_rom[ 2065]='h00002044;  wr_data_rom[ 2065]='h00003b15;
    rd_cycle[ 2066] = 1'b0;  wr_cycle[ 2066] = 1'b1;  addr_rom[ 2066]='h00002048;  wr_data_rom[ 2066]='h00001547;
    rd_cycle[ 2067] = 1'b0;  wr_cycle[ 2067] = 1'b1;  addr_rom[ 2067]='h0000204c;  wr_data_rom[ 2067]='h0000244a;
    rd_cycle[ 2068] = 1'b0;  wr_cycle[ 2068] = 1'b1;  addr_rom[ 2068]='h00002050;  wr_data_rom[ 2068]='h00001a97;
    rd_cycle[ 2069] = 1'b0;  wr_cycle[ 2069] = 1'b1;  addr_rom[ 2069]='h00002054;  wr_data_rom[ 2069]='h00003ede;
    rd_cycle[ 2070] = 1'b0;  wr_cycle[ 2070] = 1'b1;  addr_rom[ 2070]='h00002058;  wr_data_rom[ 2070]='h0000373b;
    rd_cycle[ 2071] = 1'b0;  wr_cycle[ 2071] = 1'b1;  addr_rom[ 2071]='h0000205c;  wr_data_rom[ 2071]='h000034da;
    rd_cycle[ 2072] = 1'b0;  wr_cycle[ 2072] = 1'b1;  addr_rom[ 2072]='h00002060;  wr_data_rom[ 2072]='h000005ee;
    rd_cycle[ 2073] = 1'b0;  wr_cycle[ 2073] = 1'b1;  addr_rom[ 2073]='h00002064;  wr_data_rom[ 2073]='h00000d1f;
    rd_cycle[ 2074] = 1'b0;  wr_cycle[ 2074] = 1'b1;  addr_rom[ 2074]='h00002068;  wr_data_rom[ 2074]='h000023da;
    rd_cycle[ 2075] = 1'b0;  wr_cycle[ 2075] = 1'b1;  addr_rom[ 2075]='h0000206c;  wr_data_rom[ 2075]='h00003b59;
    rd_cycle[ 2076] = 1'b0;  wr_cycle[ 2076] = 1'b1;  addr_rom[ 2076]='h00002070;  wr_data_rom[ 2076]='h000035ed;
    rd_cycle[ 2077] = 1'b0;  wr_cycle[ 2077] = 1'b1;  addr_rom[ 2077]='h00002074;  wr_data_rom[ 2077]='h00002d7d;
    rd_cycle[ 2078] = 1'b0;  wr_cycle[ 2078] = 1'b1;  addr_rom[ 2078]='h00002078;  wr_data_rom[ 2078]='h00003eff;
    rd_cycle[ 2079] = 1'b0;  wr_cycle[ 2079] = 1'b1;  addr_rom[ 2079]='h0000207c;  wr_data_rom[ 2079]='h00000e11;
    rd_cycle[ 2080] = 1'b0;  wr_cycle[ 2080] = 1'b1;  addr_rom[ 2080]='h00002080;  wr_data_rom[ 2080]='h0000361b;
    rd_cycle[ 2081] = 1'b0;  wr_cycle[ 2081] = 1'b1;  addr_rom[ 2081]='h00002084;  wr_data_rom[ 2081]='h00000e58;
    rd_cycle[ 2082] = 1'b0;  wr_cycle[ 2082] = 1'b1;  addr_rom[ 2082]='h00002088;  wr_data_rom[ 2082]='h00000896;
    rd_cycle[ 2083] = 1'b0;  wr_cycle[ 2083] = 1'b1;  addr_rom[ 2083]='h0000208c;  wr_data_rom[ 2083]='h00002c33;
    rd_cycle[ 2084] = 1'b0;  wr_cycle[ 2084] = 1'b1;  addr_rom[ 2084]='h00002090;  wr_data_rom[ 2084]='h00001bc1;
    rd_cycle[ 2085] = 1'b0;  wr_cycle[ 2085] = 1'b1;  addr_rom[ 2085]='h00002094;  wr_data_rom[ 2085]='h00002879;
    rd_cycle[ 2086] = 1'b0;  wr_cycle[ 2086] = 1'b1;  addr_rom[ 2086]='h00002098;  wr_data_rom[ 2086]='h000028b2;
    rd_cycle[ 2087] = 1'b0;  wr_cycle[ 2087] = 1'b1;  addr_rom[ 2087]='h0000209c;  wr_data_rom[ 2087]='h000038e1;
    rd_cycle[ 2088] = 1'b0;  wr_cycle[ 2088] = 1'b1;  addr_rom[ 2088]='h000020a0;  wr_data_rom[ 2088]='h000038d5;
    rd_cycle[ 2089] = 1'b0;  wr_cycle[ 2089] = 1'b1;  addr_rom[ 2089]='h000020a4;  wr_data_rom[ 2089]='h000038e1;
    rd_cycle[ 2090] = 1'b0;  wr_cycle[ 2090] = 1'b1;  addr_rom[ 2090]='h000020a8;  wr_data_rom[ 2090]='h00002c9f;
    rd_cycle[ 2091] = 1'b0;  wr_cycle[ 2091] = 1'b1;  addr_rom[ 2091]='h000020ac;  wr_data_rom[ 2091]='h00003fbc;
    rd_cycle[ 2092] = 1'b0;  wr_cycle[ 2092] = 1'b1;  addr_rom[ 2092]='h000020b0;  wr_data_rom[ 2092]='h00002eaf;
    rd_cycle[ 2093] = 1'b0;  wr_cycle[ 2093] = 1'b1;  addr_rom[ 2093]='h000020b4;  wr_data_rom[ 2093]='h00001226;
    rd_cycle[ 2094] = 1'b0;  wr_cycle[ 2094] = 1'b1;  addr_rom[ 2094]='h000020b8;  wr_data_rom[ 2094]='h00000067;
    rd_cycle[ 2095] = 1'b0;  wr_cycle[ 2095] = 1'b1;  addr_rom[ 2095]='h000020bc;  wr_data_rom[ 2095]='h00000e33;
    rd_cycle[ 2096] = 1'b0;  wr_cycle[ 2096] = 1'b1;  addr_rom[ 2096]='h000020c0;  wr_data_rom[ 2096]='h0000371e;
    rd_cycle[ 2097] = 1'b0;  wr_cycle[ 2097] = 1'b1;  addr_rom[ 2097]='h000020c4;  wr_data_rom[ 2097]='h00003c62;
    rd_cycle[ 2098] = 1'b0;  wr_cycle[ 2098] = 1'b1;  addr_rom[ 2098]='h000020c8;  wr_data_rom[ 2098]='h000005a4;
    rd_cycle[ 2099] = 1'b0;  wr_cycle[ 2099] = 1'b1;  addr_rom[ 2099]='h000020cc;  wr_data_rom[ 2099]='h00003f42;
    rd_cycle[ 2100] = 1'b0;  wr_cycle[ 2100] = 1'b1;  addr_rom[ 2100]='h000020d0;  wr_data_rom[ 2100]='h00000c21;
    rd_cycle[ 2101] = 1'b0;  wr_cycle[ 2101] = 1'b1;  addr_rom[ 2101]='h000020d4;  wr_data_rom[ 2101]='h00002c53;
    rd_cycle[ 2102] = 1'b0;  wr_cycle[ 2102] = 1'b1;  addr_rom[ 2102]='h000020d8;  wr_data_rom[ 2102]='h00003a18;
    rd_cycle[ 2103] = 1'b0;  wr_cycle[ 2103] = 1'b1;  addr_rom[ 2103]='h000020dc;  wr_data_rom[ 2103]='h00000602;
    rd_cycle[ 2104] = 1'b0;  wr_cycle[ 2104] = 1'b1;  addr_rom[ 2104]='h000020e0;  wr_data_rom[ 2104]='h00000dce;
    rd_cycle[ 2105] = 1'b0;  wr_cycle[ 2105] = 1'b1;  addr_rom[ 2105]='h000020e4;  wr_data_rom[ 2105]='h000039ef;
    rd_cycle[ 2106] = 1'b0;  wr_cycle[ 2106] = 1'b1;  addr_rom[ 2106]='h000020e8;  wr_data_rom[ 2106]='h00003a3d;
    rd_cycle[ 2107] = 1'b0;  wr_cycle[ 2107] = 1'b1;  addr_rom[ 2107]='h000020ec;  wr_data_rom[ 2107]='h00003fb8;
    rd_cycle[ 2108] = 1'b0;  wr_cycle[ 2108] = 1'b1;  addr_rom[ 2108]='h000020f0;  wr_data_rom[ 2108]='h000023b2;
    rd_cycle[ 2109] = 1'b0;  wr_cycle[ 2109] = 1'b1;  addr_rom[ 2109]='h000020f4;  wr_data_rom[ 2109]='h00000bee;
    rd_cycle[ 2110] = 1'b0;  wr_cycle[ 2110] = 1'b1;  addr_rom[ 2110]='h000020f8;  wr_data_rom[ 2110]='h000017dc;
    rd_cycle[ 2111] = 1'b0;  wr_cycle[ 2111] = 1'b1;  addr_rom[ 2111]='h000020fc;  wr_data_rom[ 2111]='h00001892;
    rd_cycle[ 2112] = 1'b0;  wr_cycle[ 2112] = 1'b1;  addr_rom[ 2112]='h00002100;  wr_data_rom[ 2112]='h00001552;
    rd_cycle[ 2113] = 1'b0;  wr_cycle[ 2113] = 1'b1;  addr_rom[ 2113]='h00002104;  wr_data_rom[ 2113]='h00003bb0;
    rd_cycle[ 2114] = 1'b0;  wr_cycle[ 2114] = 1'b1;  addr_rom[ 2114]='h00002108;  wr_data_rom[ 2114]='h0000397b;
    rd_cycle[ 2115] = 1'b0;  wr_cycle[ 2115] = 1'b1;  addr_rom[ 2115]='h0000210c;  wr_data_rom[ 2115]='h000033f8;
    rd_cycle[ 2116] = 1'b0;  wr_cycle[ 2116] = 1'b1;  addr_rom[ 2116]='h00002110;  wr_data_rom[ 2116]='h00003aa9;
    rd_cycle[ 2117] = 1'b0;  wr_cycle[ 2117] = 1'b1;  addr_rom[ 2117]='h00002114;  wr_data_rom[ 2117]='h00000f2a;
    rd_cycle[ 2118] = 1'b0;  wr_cycle[ 2118] = 1'b1;  addr_rom[ 2118]='h00002118;  wr_data_rom[ 2118]='h000036c0;
    rd_cycle[ 2119] = 1'b0;  wr_cycle[ 2119] = 1'b1;  addr_rom[ 2119]='h0000211c;  wr_data_rom[ 2119]='h000009b2;
    rd_cycle[ 2120] = 1'b0;  wr_cycle[ 2120] = 1'b1;  addr_rom[ 2120]='h00002120;  wr_data_rom[ 2120]='h0000076a;
    rd_cycle[ 2121] = 1'b0;  wr_cycle[ 2121] = 1'b1;  addr_rom[ 2121]='h00002124;  wr_data_rom[ 2121]='h000006b6;
    rd_cycle[ 2122] = 1'b0;  wr_cycle[ 2122] = 1'b1;  addr_rom[ 2122]='h00002128;  wr_data_rom[ 2122]='h00002d62;
    rd_cycle[ 2123] = 1'b0;  wr_cycle[ 2123] = 1'b1;  addr_rom[ 2123]='h0000212c;  wr_data_rom[ 2123]='h000036ac;
    rd_cycle[ 2124] = 1'b0;  wr_cycle[ 2124] = 1'b1;  addr_rom[ 2124]='h00002130;  wr_data_rom[ 2124]='h00003d37;
    rd_cycle[ 2125] = 1'b0;  wr_cycle[ 2125] = 1'b1;  addr_rom[ 2125]='h00002134;  wr_data_rom[ 2125]='h00002755;
    rd_cycle[ 2126] = 1'b0;  wr_cycle[ 2126] = 1'b1;  addr_rom[ 2126]='h00002138;  wr_data_rom[ 2126]='h00001535;
    rd_cycle[ 2127] = 1'b0;  wr_cycle[ 2127] = 1'b1;  addr_rom[ 2127]='h0000213c;  wr_data_rom[ 2127]='h0000326d;
    rd_cycle[ 2128] = 1'b0;  wr_cycle[ 2128] = 1'b1;  addr_rom[ 2128]='h00002140;  wr_data_rom[ 2128]='h00002abe;
    rd_cycle[ 2129] = 1'b0;  wr_cycle[ 2129] = 1'b1;  addr_rom[ 2129]='h00002144;  wr_data_rom[ 2129]='h00000377;
    rd_cycle[ 2130] = 1'b0;  wr_cycle[ 2130] = 1'b1;  addr_rom[ 2130]='h00002148;  wr_data_rom[ 2130]='h00002da8;
    rd_cycle[ 2131] = 1'b0;  wr_cycle[ 2131] = 1'b1;  addr_rom[ 2131]='h0000214c;  wr_data_rom[ 2131]='h000038e7;
    rd_cycle[ 2132] = 1'b0;  wr_cycle[ 2132] = 1'b1;  addr_rom[ 2132]='h00002150;  wr_data_rom[ 2132]='h00003f42;
    rd_cycle[ 2133] = 1'b0;  wr_cycle[ 2133] = 1'b1;  addr_rom[ 2133]='h00002154;  wr_data_rom[ 2133]='h00002098;
    rd_cycle[ 2134] = 1'b0;  wr_cycle[ 2134] = 1'b1;  addr_rom[ 2134]='h00002158;  wr_data_rom[ 2134]='h000033c5;
    rd_cycle[ 2135] = 1'b0;  wr_cycle[ 2135] = 1'b1;  addr_rom[ 2135]='h0000215c;  wr_data_rom[ 2135]='h00000876;
    rd_cycle[ 2136] = 1'b0;  wr_cycle[ 2136] = 1'b1;  addr_rom[ 2136]='h00002160;  wr_data_rom[ 2136]='h0000012e;
    rd_cycle[ 2137] = 1'b0;  wr_cycle[ 2137] = 1'b1;  addr_rom[ 2137]='h00002164;  wr_data_rom[ 2137]='h00001a07;
    rd_cycle[ 2138] = 1'b0;  wr_cycle[ 2138] = 1'b1;  addr_rom[ 2138]='h00002168;  wr_data_rom[ 2138]='h000019ee;
    rd_cycle[ 2139] = 1'b0;  wr_cycle[ 2139] = 1'b1;  addr_rom[ 2139]='h0000216c;  wr_data_rom[ 2139]='h000014c0;
    rd_cycle[ 2140] = 1'b0;  wr_cycle[ 2140] = 1'b1;  addr_rom[ 2140]='h00002170;  wr_data_rom[ 2140]='h00001ca2;
    rd_cycle[ 2141] = 1'b0;  wr_cycle[ 2141] = 1'b1;  addr_rom[ 2141]='h00002174;  wr_data_rom[ 2141]='h000038f7;
    rd_cycle[ 2142] = 1'b0;  wr_cycle[ 2142] = 1'b1;  addr_rom[ 2142]='h00002178;  wr_data_rom[ 2142]='h000027de;
    rd_cycle[ 2143] = 1'b0;  wr_cycle[ 2143] = 1'b1;  addr_rom[ 2143]='h0000217c;  wr_data_rom[ 2143]='h00001d87;
    rd_cycle[ 2144] = 1'b0;  wr_cycle[ 2144] = 1'b1;  addr_rom[ 2144]='h00002180;  wr_data_rom[ 2144]='h00000a62;
    rd_cycle[ 2145] = 1'b0;  wr_cycle[ 2145] = 1'b1;  addr_rom[ 2145]='h00002184;  wr_data_rom[ 2145]='h00001ce0;
    rd_cycle[ 2146] = 1'b0;  wr_cycle[ 2146] = 1'b1;  addr_rom[ 2146]='h00002188;  wr_data_rom[ 2146]='h0000335d;
    rd_cycle[ 2147] = 1'b0;  wr_cycle[ 2147] = 1'b1;  addr_rom[ 2147]='h0000218c;  wr_data_rom[ 2147]='h00001cb1;
    rd_cycle[ 2148] = 1'b0;  wr_cycle[ 2148] = 1'b1;  addr_rom[ 2148]='h00002190;  wr_data_rom[ 2148]='h000021b2;
    rd_cycle[ 2149] = 1'b0;  wr_cycle[ 2149] = 1'b1;  addr_rom[ 2149]='h00002194;  wr_data_rom[ 2149]='h0000332a;
    rd_cycle[ 2150] = 1'b0;  wr_cycle[ 2150] = 1'b1;  addr_rom[ 2150]='h00002198;  wr_data_rom[ 2150]='h00000be1;
    rd_cycle[ 2151] = 1'b0;  wr_cycle[ 2151] = 1'b1;  addr_rom[ 2151]='h0000219c;  wr_data_rom[ 2151]='h00003e2a;
    rd_cycle[ 2152] = 1'b0;  wr_cycle[ 2152] = 1'b1;  addr_rom[ 2152]='h000021a0;  wr_data_rom[ 2152]='h00001f35;
    rd_cycle[ 2153] = 1'b0;  wr_cycle[ 2153] = 1'b1;  addr_rom[ 2153]='h000021a4;  wr_data_rom[ 2153]='h000033a2;
    rd_cycle[ 2154] = 1'b0;  wr_cycle[ 2154] = 1'b1;  addr_rom[ 2154]='h000021a8;  wr_data_rom[ 2154]='h000017e7;
    rd_cycle[ 2155] = 1'b0;  wr_cycle[ 2155] = 1'b1;  addr_rom[ 2155]='h000021ac;  wr_data_rom[ 2155]='h00000daf;
    rd_cycle[ 2156] = 1'b0;  wr_cycle[ 2156] = 1'b1;  addr_rom[ 2156]='h000021b0;  wr_data_rom[ 2156]='h00002e76;
    rd_cycle[ 2157] = 1'b0;  wr_cycle[ 2157] = 1'b1;  addr_rom[ 2157]='h000021b4;  wr_data_rom[ 2157]='h00001bd9;
    rd_cycle[ 2158] = 1'b0;  wr_cycle[ 2158] = 1'b1;  addr_rom[ 2158]='h000021b8;  wr_data_rom[ 2158]='h0000228d;
    rd_cycle[ 2159] = 1'b0;  wr_cycle[ 2159] = 1'b1;  addr_rom[ 2159]='h000021bc;  wr_data_rom[ 2159]='h00002d20;
    rd_cycle[ 2160] = 1'b0;  wr_cycle[ 2160] = 1'b1;  addr_rom[ 2160]='h000021c0;  wr_data_rom[ 2160]='h00001fec;
    rd_cycle[ 2161] = 1'b0;  wr_cycle[ 2161] = 1'b1;  addr_rom[ 2161]='h000021c4;  wr_data_rom[ 2161]='h0000076a;
    rd_cycle[ 2162] = 1'b0;  wr_cycle[ 2162] = 1'b1;  addr_rom[ 2162]='h000021c8;  wr_data_rom[ 2162]='h000012c6;
    rd_cycle[ 2163] = 1'b0;  wr_cycle[ 2163] = 1'b1;  addr_rom[ 2163]='h000021cc;  wr_data_rom[ 2163]='h000034d8;
    rd_cycle[ 2164] = 1'b0;  wr_cycle[ 2164] = 1'b1;  addr_rom[ 2164]='h000021d0;  wr_data_rom[ 2164]='h00002d34;
    rd_cycle[ 2165] = 1'b0;  wr_cycle[ 2165] = 1'b1;  addr_rom[ 2165]='h000021d4;  wr_data_rom[ 2165]='h000008ae;
    rd_cycle[ 2166] = 1'b0;  wr_cycle[ 2166] = 1'b1;  addr_rom[ 2166]='h000021d8;  wr_data_rom[ 2166]='h00001561;
    rd_cycle[ 2167] = 1'b0;  wr_cycle[ 2167] = 1'b1;  addr_rom[ 2167]='h000021dc;  wr_data_rom[ 2167]='h00000bee;
    rd_cycle[ 2168] = 1'b0;  wr_cycle[ 2168] = 1'b1;  addr_rom[ 2168]='h000021e0;  wr_data_rom[ 2168]='h00001aa9;
    rd_cycle[ 2169] = 1'b0;  wr_cycle[ 2169] = 1'b1;  addr_rom[ 2169]='h000021e4;  wr_data_rom[ 2169]='h00001552;
    rd_cycle[ 2170] = 1'b0;  wr_cycle[ 2170] = 1'b1;  addr_rom[ 2170]='h000021e8;  wr_data_rom[ 2170]='h0000351f;
    rd_cycle[ 2171] = 1'b0;  wr_cycle[ 2171] = 1'b1;  addr_rom[ 2171]='h000021ec;  wr_data_rom[ 2171]='h00000023;
    rd_cycle[ 2172] = 1'b0;  wr_cycle[ 2172] = 1'b1;  addr_rom[ 2172]='h000021f0;  wr_data_rom[ 2172]='h00000347;
    rd_cycle[ 2173] = 1'b0;  wr_cycle[ 2173] = 1'b1;  addr_rom[ 2173]='h000021f4;  wr_data_rom[ 2173]='h00002180;
    rd_cycle[ 2174] = 1'b0;  wr_cycle[ 2174] = 1'b1;  addr_rom[ 2174]='h000021f8;  wr_data_rom[ 2174]='h00000e3b;
    rd_cycle[ 2175] = 1'b0;  wr_cycle[ 2175] = 1'b1;  addr_rom[ 2175]='h000021fc;  wr_data_rom[ 2175]='h00002319;
    rd_cycle[ 2176] = 1'b0;  wr_cycle[ 2176] = 1'b1;  addr_rom[ 2176]='h00002200;  wr_data_rom[ 2176]='h000029dc;
    rd_cycle[ 2177] = 1'b0;  wr_cycle[ 2177] = 1'b1;  addr_rom[ 2177]='h00002204;  wr_data_rom[ 2177]='h00001da3;
    rd_cycle[ 2178] = 1'b0;  wr_cycle[ 2178] = 1'b1;  addr_rom[ 2178]='h00002208;  wr_data_rom[ 2178]='h00000a98;
    rd_cycle[ 2179] = 1'b0;  wr_cycle[ 2179] = 1'b1;  addr_rom[ 2179]='h0000220c;  wr_data_rom[ 2179]='h00002bfe;
    rd_cycle[ 2180] = 1'b0;  wr_cycle[ 2180] = 1'b1;  addr_rom[ 2180]='h00002210;  wr_data_rom[ 2180]='h0000037a;
    rd_cycle[ 2181] = 1'b0;  wr_cycle[ 2181] = 1'b1;  addr_rom[ 2181]='h00002214;  wr_data_rom[ 2181]='h00000fb5;
    rd_cycle[ 2182] = 1'b0;  wr_cycle[ 2182] = 1'b1;  addr_rom[ 2182]='h00002218;  wr_data_rom[ 2182]='h00002d58;
    rd_cycle[ 2183] = 1'b0;  wr_cycle[ 2183] = 1'b1;  addr_rom[ 2183]='h0000221c;  wr_data_rom[ 2183]='h00002ae0;
    rd_cycle[ 2184] = 1'b0;  wr_cycle[ 2184] = 1'b1;  addr_rom[ 2184]='h00002220;  wr_data_rom[ 2184]='h00001e85;
    rd_cycle[ 2185] = 1'b0;  wr_cycle[ 2185] = 1'b1;  addr_rom[ 2185]='h00002224;  wr_data_rom[ 2185]='h00001c4f;
    rd_cycle[ 2186] = 1'b0;  wr_cycle[ 2186] = 1'b1;  addr_rom[ 2186]='h00002228;  wr_data_rom[ 2186]='h0000225e;
    rd_cycle[ 2187] = 1'b0;  wr_cycle[ 2187] = 1'b1;  addr_rom[ 2187]='h0000222c;  wr_data_rom[ 2187]='h000026ba;
    rd_cycle[ 2188] = 1'b0;  wr_cycle[ 2188] = 1'b1;  addr_rom[ 2188]='h00002230;  wr_data_rom[ 2188]='h00000c91;
    rd_cycle[ 2189] = 1'b0;  wr_cycle[ 2189] = 1'b1;  addr_rom[ 2189]='h00002234;  wr_data_rom[ 2189]='h000038bf;
    rd_cycle[ 2190] = 1'b0;  wr_cycle[ 2190] = 1'b1;  addr_rom[ 2190]='h00002238;  wr_data_rom[ 2190]='h000015e4;
    rd_cycle[ 2191] = 1'b0;  wr_cycle[ 2191] = 1'b1;  addr_rom[ 2191]='h0000223c;  wr_data_rom[ 2191]='h00002e17;
    rd_cycle[ 2192] = 1'b0;  wr_cycle[ 2192] = 1'b1;  addr_rom[ 2192]='h00002240;  wr_data_rom[ 2192]='h000009fb;
    rd_cycle[ 2193] = 1'b0;  wr_cycle[ 2193] = 1'b1;  addr_rom[ 2193]='h00002244;  wr_data_rom[ 2193]='h00003d84;
    rd_cycle[ 2194] = 1'b0;  wr_cycle[ 2194] = 1'b1;  addr_rom[ 2194]='h00002248;  wr_data_rom[ 2194]='h00001aa3;
    rd_cycle[ 2195] = 1'b0;  wr_cycle[ 2195] = 1'b1;  addr_rom[ 2195]='h0000224c;  wr_data_rom[ 2195]='h000019ad;
    rd_cycle[ 2196] = 1'b0;  wr_cycle[ 2196] = 1'b1;  addr_rom[ 2196]='h00002250;  wr_data_rom[ 2196]='h00003883;
    rd_cycle[ 2197] = 1'b0;  wr_cycle[ 2197] = 1'b1;  addr_rom[ 2197]='h00002254;  wr_data_rom[ 2197]='h00000159;
    rd_cycle[ 2198] = 1'b0;  wr_cycle[ 2198] = 1'b1;  addr_rom[ 2198]='h00002258;  wr_data_rom[ 2198]='h000014f1;
    rd_cycle[ 2199] = 1'b0;  wr_cycle[ 2199] = 1'b1;  addr_rom[ 2199]='h0000225c;  wr_data_rom[ 2199]='h00003cab;
    rd_cycle[ 2200] = 1'b0;  wr_cycle[ 2200] = 1'b1;  addr_rom[ 2200]='h00002260;  wr_data_rom[ 2200]='h000022d2;
    rd_cycle[ 2201] = 1'b0;  wr_cycle[ 2201] = 1'b1;  addr_rom[ 2201]='h00002264;  wr_data_rom[ 2201]='h00002660;
    rd_cycle[ 2202] = 1'b0;  wr_cycle[ 2202] = 1'b1;  addr_rom[ 2202]='h00002268;  wr_data_rom[ 2202]='h00000485;
    rd_cycle[ 2203] = 1'b0;  wr_cycle[ 2203] = 1'b1;  addr_rom[ 2203]='h0000226c;  wr_data_rom[ 2203]='h00001859;
    rd_cycle[ 2204] = 1'b0;  wr_cycle[ 2204] = 1'b1;  addr_rom[ 2204]='h00002270;  wr_data_rom[ 2204]='h00000163;
    rd_cycle[ 2205] = 1'b0;  wr_cycle[ 2205] = 1'b1;  addr_rom[ 2205]='h00002274;  wr_data_rom[ 2205]='h000017e5;
    rd_cycle[ 2206] = 1'b0;  wr_cycle[ 2206] = 1'b1;  addr_rom[ 2206]='h00002278;  wr_data_rom[ 2206]='h0000224b;
    rd_cycle[ 2207] = 1'b0;  wr_cycle[ 2207] = 1'b1;  addr_rom[ 2207]='h0000227c;  wr_data_rom[ 2207]='h0000091e;
    rd_cycle[ 2208] = 1'b0;  wr_cycle[ 2208] = 1'b1;  addr_rom[ 2208]='h00002280;  wr_data_rom[ 2208]='h0000179b;
    rd_cycle[ 2209] = 1'b0;  wr_cycle[ 2209] = 1'b1;  addr_rom[ 2209]='h00002284;  wr_data_rom[ 2209]='h00002e8d;
    rd_cycle[ 2210] = 1'b0;  wr_cycle[ 2210] = 1'b1;  addr_rom[ 2210]='h00002288;  wr_data_rom[ 2210]='h00003977;
    rd_cycle[ 2211] = 1'b0;  wr_cycle[ 2211] = 1'b1;  addr_rom[ 2211]='h0000228c;  wr_data_rom[ 2211]='h00002667;
    rd_cycle[ 2212] = 1'b0;  wr_cycle[ 2212] = 1'b1;  addr_rom[ 2212]='h00002290;  wr_data_rom[ 2212]='h0000393a;
    rd_cycle[ 2213] = 1'b0;  wr_cycle[ 2213] = 1'b1;  addr_rom[ 2213]='h00002294;  wr_data_rom[ 2213]='h00000a36;
    rd_cycle[ 2214] = 1'b0;  wr_cycle[ 2214] = 1'b1;  addr_rom[ 2214]='h00002298;  wr_data_rom[ 2214]='h00000dea;
    rd_cycle[ 2215] = 1'b0;  wr_cycle[ 2215] = 1'b1;  addr_rom[ 2215]='h0000229c;  wr_data_rom[ 2215]='h00000261;
    rd_cycle[ 2216] = 1'b0;  wr_cycle[ 2216] = 1'b1;  addr_rom[ 2216]='h000022a0;  wr_data_rom[ 2216]='h000017b1;
    rd_cycle[ 2217] = 1'b0;  wr_cycle[ 2217] = 1'b1;  addr_rom[ 2217]='h000022a4;  wr_data_rom[ 2217]='h00000e92;
    rd_cycle[ 2218] = 1'b0;  wr_cycle[ 2218] = 1'b1;  addr_rom[ 2218]='h000022a8;  wr_data_rom[ 2218]='h00002754;
    rd_cycle[ 2219] = 1'b0;  wr_cycle[ 2219] = 1'b1;  addr_rom[ 2219]='h000022ac;  wr_data_rom[ 2219]='h00003302;
    rd_cycle[ 2220] = 1'b0;  wr_cycle[ 2220] = 1'b1;  addr_rom[ 2220]='h000022b0;  wr_data_rom[ 2220]='h0000278e;
    rd_cycle[ 2221] = 1'b0;  wr_cycle[ 2221] = 1'b1;  addr_rom[ 2221]='h000022b4;  wr_data_rom[ 2221]='h00003304;
    rd_cycle[ 2222] = 1'b0;  wr_cycle[ 2222] = 1'b1;  addr_rom[ 2222]='h000022b8;  wr_data_rom[ 2222]='h00003b9c;
    rd_cycle[ 2223] = 1'b0;  wr_cycle[ 2223] = 1'b1;  addr_rom[ 2223]='h000022bc;  wr_data_rom[ 2223]='h0000083b;
    rd_cycle[ 2224] = 1'b0;  wr_cycle[ 2224] = 1'b1;  addr_rom[ 2224]='h000022c0;  wr_data_rom[ 2224]='h00001525;
    rd_cycle[ 2225] = 1'b0;  wr_cycle[ 2225] = 1'b1;  addr_rom[ 2225]='h000022c4;  wr_data_rom[ 2225]='h00001fd0;
    rd_cycle[ 2226] = 1'b0;  wr_cycle[ 2226] = 1'b1;  addr_rom[ 2226]='h000022c8;  wr_data_rom[ 2226]='h00003589;
    rd_cycle[ 2227] = 1'b0;  wr_cycle[ 2227] = 1'b1;  addr_rom[ 2227]='h000022cc;  wr_data_rom[ 2227]='h0000361c;
    rd_cycle[ 2228] = 1'b0;  wr_cycle[ 2228] = 1'b1;  addr_rom[ 2228]='h000022d0;  wr_data_rom[ 2228]='h00003cec;
    rd_cycle[ 2229] = 1'b0;  wr_cycle[ 2229] = 1'b1;  addr_rom[ 2229]='h000022d4;  wr_data_rom[ 2229]='h00001fcf;
    rd_cycle[ 2230] = 1'b0;  wr_cycle[ 2230] = 1'b1;  addr_rom[ 2230]='h000022d8;  wr_data_rom[ 2230]='h00001d23;
    rd_cycle[ 2231] = 1'b0;  wr_cycle[ 2231] = 1'b1;  addr_rom[ 2231]='h000022dc;  wr_data_rom[ 2231]='h00000db7;
    rd_cycle[ 2232] = 1'b0;  wr_cycle[ 2232] = 1'b1;  addr_rom[ 2232]='h000022e0;  wr_data_rom[ 2232]='h00001d2e;
    rd_cycle[ 2233] = 1'b0;  wr_cycle[ 2233] = 1'b1;  addr_rom[ 2233]='h000022e4;  wr_data_rom[ 2233]='h00001a94;
    rd_cycle[ 2234] = 1'b0;  wr_cycle[ 2234] = 1'b1;  addr_rom[ 2234]='h000022e8;  wr_data_rom[ 2234]='h0000304a;
    rd_cycle[ 2235] = 1'b0;  wr_cycle[ 2235] = 1'b1;  addr_rom[ 2235]='h000022ec;  wr_data_rom[ 2235]='h00003d62;
    rd_cycle[ 2236] = 1'b0;  wr_cycle[ 2236] = 1'b1;  addr_rom[ 2236]='h000022f0;  wr_data_rom[ 2236]='h000002b4;
    rd_cycle[ 2237] = 1'b0;  wr_cycle[ 2237] = 1'b1;  addr_rom[ 2237]='h000022f4;  wr_data_rom[ 2237]='h00000db3;
    rd_cycle[ 2238] = 1'b0;  wr_cycle[ 2238] = 1'b1;  addr_rom[ 2238]='h000022f8;  wr_data_rom[ 2238]='h00001c89;
    rd_cycle[ 2239] = 1'b0;  wr_cycle[ 2239] = 1'b1;  addr_rom[ 2239]='h000022fc;  wr_data_rom[ 2239]='h00000e85;
    rd_cycle[ 2240] = 1'b0;  wr_cycle[ 2240] = 1'b1;  addr_rom[ 2240]='h00002300;  wr_data_rom[ 2240]='h00001284;
    rd_cycle[ 2241] = 1'b0;  wr_cycle[ 2241] = 1'b1;  addr_rom[ 2241]='h00002304;  wr_data_rom[ 2241]='h00000e4c;
    rd_cycle[ 2242] = 1'b0;  wr_cycle[ 2242] = 1'b1;  addr_rom[ 2242]='h00002308;  wr_data_rom[ 2242]='h00002af2;
    rd_cycle[ 2243] = 1'b0;  wr_cycle[ 2243] = 1'b1;  addr_rom[ 2243]='h0000230c;  wr_data_rom[ 2243]='h00002cbd;
    rd_cycle[ 2244] = 1'b0;  wr_cycle[ 2244] = 1'b1;  addr_rom[ 2244]='h00002310;  wr_data_rom[ 2244]='h00003333;
    rd_cycle[ 2245] = 1'b0;  wr_cycle[ 2245] = 1'b1;  addr_rom[ 2245]='h00002314;  wr_data_rom[ 2245]='h00002d64;
    rd_cycle[ 2246] = 1'b0;  wr_cycle[ 2246] = 1'b1;  addr_rom[ 2246]='h00002318;  wr_data_rom[ 2246]='h00002194;
    rd_cycle[ 2247] = 1'b0;  wr_cycle[ 2247] = 1'b1;  addr_rom[ 2247]='h0000231c;  wr_data_rom[ 2247]='h00001882;
    rd_cycle[ 2248] = 1'b0;  wr_cycle[ 2248] = 1'b1;  addr_rom[ 2248]='h00002320;  wr_data_rom[ 2248]='h0000297c;
    rd_cycle[ 2249] = 1'b0;  wr_cycle[ 2249] = 1'b1;  addr_rom[ 2249]='h00002324;  wr_data_rom[ 2249]='h0000383f;
    rd_cycle[ 2250] = 1'b0;  wr_cycle[ 2250] = 1'b1;  addr_rom[ 2250]='h00002328;  wr_data_rom[ 2250]='h00003423;
    rd_cycle[ 2251] = 1'b0;  wr_cycle[ 2251] = 1'b1;  addr_rom[ 2251]='h0000232c;  wr_data_rom[ 2251]='h00003604;
    rd_cycle[ 2252] = 1'b0;  wr_cycle[ 2252] = 1'b1;  addr_rom[ 2252]='h00002330;  wr_data_rom[ 2252]='h00003d92;
    rd_cycle[ 2253] = 1'b0;  wr_cycle[ 2253] = 1'b1;  addr_rom[ 2253]='h00002334;  wr_data_rom[ 2253]='h000031a3;
    rd_cycle[ 2254] = 1'b0;  wr_cycle[ 2254] = 1'b1;  addr_rom[ 2254]='h00002338;  wr_data_rom[ 2254]='h00001dda;
    rd_cycle[ 2255] = 1'b0;  wr_cycle[ 2255] = 1'b1;  addr_rom[ 2255]='h0000233c;  wr_data_rom[ 2255]='h000023b0;
    rd_cycle[ 2256] = 1'b0;  wr_cycle[ 2256] = 1'b1;  addr_rom[ 2256]='h00002340;  wr_data_rom[ 2256]='h00002361;
    rd_cycle[ 2257] = 1'b0;  wr_cycle[ 2257] = 1'b1;  addr_rom[ 2257]='h00002344;  wr_data_rom[ 2257]='h00000ca7;
    rd_cycle[ 2258] = 1'b0;  wr_cycle[ 2258] = 1'b1;  addr_rom[ 2258]='h00002348;  wr_data_rom[ 2258]='h00001d86;
    rd_cycle[ 2259] = 1'b0;  wr_cycle[ 2259] = 1'b1;  addr_rom[ 2259]='h0000234c;  wr_data_rom[ 2259]='h00003800;
    rd_cycle[ 2260] = 1'b0;  wr_cycle[ 2260] = 1'b1;  addr_rom[ 2260]='h00002350;  wr_data_rom[ 2260]='h000000a9;
    rd_cycle[ 2261] = 1'b0;  wr_cycle[ 2261] = 1'b1;  addr_rom[ 2261]='h00002354;  wr_data_rom[ 2261]='h00001c5f;
    rd_cycle[ 2262] = 1'b0;  wr_cycle[ 2262] = 1'b1;  addr_rom[ 2262]='h00002358;  wr_data_rom[ 2262]='h00002a46;
    rd_cycle[ 2263] = 1'b0;  wr_cycle[ 2263] = 1'b1;  addr_rom[ 2263]='h0000235c;  wr_data_rom[ 2263]='h0000023a;
    rd_cycle[ 2264] = 1'b0;  wr_cycle[ 2264] = 1'b1;  addr_rom[ 2264]='h00002360;  wr_data_rom[ 2264]='h00003574;
    rd_cycle[ 2265] = 1'b0;  wr_cycle[ 2265] = 1'b1;  addr_rom[ 2265]='h00002364;  wr_data_rom[ 2265]='h00002ff0;
    rd_cycle[ 2266] = 1'b0;  wr_cycle[ 2266] = 1'b1;  addr_rom[ 2266]='h00002368;  wr_data_rom[ 2266]='h00003312;
    rd_cycle[ 2267] = 1'b0;  wr_cycle[ 2267] = 1'b1;  addr_rom[ 2267]='h0000236c;  wr_data_rom[ 2267]='h00003cf9;
    rd_cycle[ 2268] = 1'b0;  wr_cycle[ 2268] = 1'b1;  addr_rom[ 2268]='h00002370;  wr_data_rom[ 2268]='h00000464;
    rd_cycle[ 2269] = 1'b0;  wr_cycle[ 2269] = 1'b1;  addr_rom[ 2269]='h00002374;  wr_data_rom[ 2269]='h00002c4a;
    rd_cycle[ 2270] = 1'b0;  wr_cycle[ 2270] = 1'b1;  addr_rom[ 2270]='h00002378;  wr_data_rom[ 2270]='h00002de4;
    rd_cycle[ 2271] = 1'b0;  wr_cycle[ 2271] = 1'b1;  addr_rom[ 2271]='h0000237c;  wr_data_rom[ 2271]='h0000260d;
    rd_cycle[ 2272] = 1'b0;  wr_cycle[ 2272] = 1'b1;  addr_rom[ 2272]='h00002380;  wr_data_rom[ 2272]='h00000805;
    rd_cycle[ 2273] = 1'b0;  wr_cycle[ 2273] = 1'b1;  addr_rom[ 2273]='h00002384;  wr_data_rom[ 2273]='h00002cbe;
    rd_cycle[ 2274] = 1'b0;  wr_cycle[ 2274] = 1'b1;  addr_rom[ 2274]='h00002388;  wr_data_rom[ 2274]='h00002fd6;
    rd_cycle[ 2275] = 1'b0;  wr_cycle[ 2275] = 1'b1;  addr_rom[ 2275]='h0000238c;  wr_data_rom[ 2275]='h000000ac;
    rd_cycle[ 2276] = 1'b0;  wr_cycle[ 2276] = 1'b1;  addr_rom[ 2276]='h00002390;  wr_data_rom[ 2276]='h00000060;
    rd_cycle[ 2277] = 1'b0;  wr_cycle[ 2277] = 1'b1;  addr_rom[ 2277]='h00002394;  wr_data_rom[ 2277]='h000030f7;
    rd_cycle[ 2278] = 1'b0;  wr_cycle[ 2278] = 1'b1;  addr_rom[ 2278]='h00002398;  wr_data_rom[ 2278]='h00001f4c;
    rd_cycle[ 2279] = 1'b0;  wr_cycle[ 2279] = 1'b1;  addr_rom[ 2279]='h0000239c;  wr_data_rom[ 2279]='h00002b79;
    rd_cycle[ 2280] = 1'b0;  wr_cycle[ 2280] = 1'b1;  addr_rom[ 2280]='h000023a0;  wr_data_rom[ 2280]='h0000232f;
    rd_cycle[ 2281] = 1'b0;  wr_cycle[ 2281] = 1'b1;  addr_rom[ 2281]='h000023a4;  wr_data_rom[ 2281]='h000018e9;
    rd_cycle[ 2282] = 1'b0;  wr_cycle[ 2282] = 1'b1;  addr_rom[ 2282]='h000023a8;  wr_data_rom[ 2282]='h00001dd2;
    rd_cycle[ 2283] = 1'b0;  wr_cycle[ 2283] = 1'b1;  addr_rom[ 2283]='h000023ac;  wr_data_rom[ 2283]='h00002bca;
    rd_cycle[ 2284] = 1'b0;  wr_cycle[ 2284] = 1'b1;  addr_rom[ 2284]='h000023b0;  wr_data_rom[ 2284]='h00002626;
    rd_cycle[ 2285] = 1'b0;  wr_cycle[ 2285] = 1'b1;  addr_rom[ 2285]='h000023b4;  wr_data_rom[ 2285]='h00000e5d;
    rd_cycle[ 2286] = 1'b0;  wr_cycle[ 2286] = 1'b1;  addr_rom[ 2286]='h000023b8;  wr_data_rom[ 2286]='h000035ee;
    rd_cycle[ 2287] = 1'b0;  wr_cycle[ 2287] = 1'b1;  addr_rom[ 2287]='h000023bc;  wr_data_rom[ 2287]='h00002663;
    rd_cycle[ 2288] = 1'b0;  wr_cycle[ 2288] = 1'b1;  addr_rom[ 2288]='h000023c0;  wr_data_rom[ 2288]='h00001706;
    rd_cycle[ 2289] = 1'b0;  wr_cycle[ 2289] = 1'b1;  addr_rom[ 2289]='h000023c4;  wr_data_rom[ 2289]='h000005cd;
    rd_cycle[ 2290] = 1'b0;  wr_cycle[ 2290] = 1'b1;  addr_rom[ 2290]='h000023c8;  wr_data_rom[ 2290]='h00001c2b;
    rd_cycle[ 2291] = 1'b0;  wr_cycle[ 2291] = 1'b1;  addr_rom[ 2291]='h000023cc;  wr_data_rom[ 2291]='h00001dc7;
    rd_cycle[ 2292] = 1'b0;  wr_cycle[ 2292] = 1'b1;  addr_rom[ 2292]='h000023d0;  wr_data_rom[ 2292]='h00002488;
    rd_cycle[ 2293] = 1'b0;  wr_cycle[ 2293] = 1'b1;  addr_rom[ 2293]='h000023d4;  wr_data_rom[ 2293]='h00002422;
    rd_cycle[ 2294] = 1'b0;  wr_cycle[ 2294] = 1'b1;  addr_rom[ 2294]='h000023d8;  wr_data_rom[ 2294]='h00001933;
    rd_cycle[ 2295] = 1'b0;  wr_cycle[ 2295] = 1'b1;  addr_rom[ 2295]='h000023dc;  wr_data_rom[ 2295]='h00000d50;
    rd_cycle[ 2296] = 1'b0;  wr_cycle[ 2296] = 1'b1;  addr_rom[ 2296]='h000023e0;  wr_data_rom[ 2296]='h00003d93;
    rd_cycle[ 2297] = 1'b0;  wr_cycle[ 2297] = 1'b1;  addr_rom[ 2297]='h000023e4;  wr_data_rom[ 2297]='h000012d5;
    rd_cycle[ 2298] = 1'b0;  wr_cycle[ 2298] = 1'b1;  addr_rom[ 2298]='h000023e8;  wr_data_rom[ 2298]='h00001fef;
    rd_cycle[ 2299] = 1'b0;  wr_cycle[ 2299] = 1'b1;  addr_rom[ 2299]='h000023ec;  wr_data_rom[ 2299]='h0000166f;
    rd_cycle[ 2300] = 1'b0;  wr_cycle[ 2300] = 1'b1;  addr_rom[ 2300]='h000023f0;  wr_data_rom[ 2300]='h00001e57;
    rd_cycle[ 2301] = 1'b0;  wr_cycle[ 2301] = 1'b1;  addr_rom[ 2301]='h000023f4;  wr_data_rom[ 2301]='h00000568;
    rd_cycle[ 2302] = 1'b0;  wr_cycle[ 2302] = 1'b1;  addr_rom[ 2302]='h000023f8;  wr_data_rom[ 2302]='h000012d5;
    rd_cycle[ 2303] = 1'b0;  wr_cycle[ 2303] = 1'b1;  addr_rom[ 2303]='h000023fc;  wr_data_rom[ 2303]='h00000176;
    rd_cycle[ 2304] = 1'b0;  wr_cycle[ 2304] = 1'b1;  addr_rom[ 2304]='h00002400;  wr_data_rom[ 2304]='h00001a83;
    rd_cycle[ 2305] = 1'b0;  wr_cycle[ 2305] = 1'b1;  addr_rom[ 2305]='h00002404;  wr_data_rom[ 2305]='h00001367;
    rd_cycle[ 2306] = 1'b0;  wr_cycle[ 2306] = 1'b1;  addr_rom[ 2306]='h00002408;  wr_data_rom[ 2306]='h000017e9;
    rd_cycle[ 2307] = 1'b0;  wr_cycle[ 2307] = 1'b1;  addr_rom[ 2307]='h0000240c;  wr_data_rom[ 2307]='h0000277a;
    rd_cycle[ 2308] = 1'b0;  wr_cycle[ 2308] = 1'b1;  addr_rom[ 2308]='h00002410;  wr_data_rom[ 2308]='h000015f0;
    rd_cycle[ 2309] = 1'b0;  wr_cycle[ 2309] = 1'b1;  addr_rom[ 2309]='h00002414;  wr_data_rom[ 2309]='h000004c5;
    rd_cycle[ 2310] = 1'b0;  wr_cycle[ 2310] = 1'b1;  addr_rom[ 2310]='h00002418;  wr_data_rom[ 2310]='h00003164;
    rd_cycle[ 2311] = 1'b0;  wr_cycle[ 2311] = 1'b1;  addr_rom[ 2311]='h0000241c;  wr_data_rom[ 2311]='h000005a8;
    rd_cycle[ 2312] = 1'b0;  wr_cycle[ 2312] = 1'b1;  addr_rom[ 2312]='h00002420;  wr_data_rom[ 2312]='h00003bc2;
    rd_cycle[ 2313] = 1'b0;  wr_cycle[ 2313] = 1'b1;  addr_rom[ 2313]='h00002424;  wr_data_rom[ 2313]='h00000f2f;
    rd_cycle[ 2314] = 1'b0;  wr_cycle[ 2314] = 1'b1;  addr_rom[ 2314]='h00002428;  wr_data_rom[ 2314]='h00001cf0;
    rd_cycle[ 2315] = 1'b0;  wr_cycle[ 2315] = 1'b1;  addr_rom[ 2315]='h0000242c;  wr_data_rom[ 2315]='h00002bc2;
    rd_cycle[ 2316] = 1'b0;  wr_cycle[ 2316] = 1'b1;  addr_rom[ 2316]='h00002430;  wr_data_rom[ 2316]='h000031d3;
    rd_cycle[ 2317] = 1'b0;  wr_cycle[ 2317] = 1'b1;  addr_rom[ 2317]='h00002434;  wr_data_rom[ 2317]='h00000fc8;
    rd_cycle[ 2318] = 1'b0;  wr_cycle[ 2318] = 1'b1;  addr_rom[ 2318]='h00002438;  wr_data_rom[ 2318]='h00001059;
    rd_cycle[ 2319] = 1'b0;  wr_cycle[ 2319] = 1'b1;  addr_rom[ 2319]='h0000243c;  wr_data_rom[ 2319]='h00003f2e;
    rd_cycle[ 2320] = 1'b0;  wr_cycle[ 2320] = 1'b1;  addr_rom[ 2320]='h00002440;  wr_data_rom[ 2320]='h00000fc4;
    rd_cycle[ 2321] = 1'b0;  wr_cycle[ 2321] = 1'b1;  addr_rom[ 2321]='h00002444;  wr_data_rom[ 2321]='h00001e1b;
    rd_cycle[ 2322] = 1'b0;  wr_cycle[ 2322] = 1'b1;  addr_rom[ 2322]='h00002448;  wr_data_rom[ 2322]='h0000157a;
    rd_cycle[ 2323] = 1'b0;  wr_cycle[ 2323] = 1'b1;  addr_rom[ 2323]='h0000244c;  wr_data_rom[ 2323]='h00003a65;
    rd_cycle[ 2324] = 1'b0;  wr_cycle[ 2324] = 1'b1;  addr_rom[ 2324]='h00002450;  wr_data_rom[ 2324]='h000013ae;
    rd_cycle[ 2325] = 1'b0;  wr_cycle[ 2325] = 1'b1;  addr_rom[ 2325]='h00002454;  wr_data_rom[ 2325]='h0000395a;
    rd_cycle[ 2326] = 1'b0;  wr_cycle[ 2326] = 1'b1;  addr_rom[ 2326]='h00002458;  wr_data_rom[ 2326]='h00002726;
    rd_cycle[ 2327] = 1'b0;  wr_cycle[ 2327] = 1'b1;  addr_rom[ 2327]='h0000245c;  wr_data_rom[ 2327]='h00000a7e;
    rd_cycle[ 2328] = 1'b0;  wr_cycle[ 2328] = 1'b1;  addr_rom[ 2328]='h00002460;  wr_data_rom[ 2328]='h00002cd2;
    rd_cycle[ 2329] = 1'b0;  wr_cycle[ 2329] = 1'b1;  addr_rom[ 2329]='h00002464;  wr_data_rom[ 2329]='h00002b66;
    rd_cycle[ 2330] = 1'b0;  wr_cycle[ 2330] = 1'b1;  addr_rom[ 2330]='h00002468;  wr_data_rom[ 2330]='h00003ea3;
    rd_cycle[ 2331] = 1'b0;  wr_cycle[ 2331] = 1'b1;  addr_rom[ 2331]='h0000246c;  wr_data_rom[ 2331]='h00000822;
    rd_cycle[ 2332] = 1'b0;  wr_cycle[ 2332] = 1'b1;  addr_rom[ 2332]='h00002470;  wr_data_rom[ 2332]='h0000340b;
    rd_cycle[ 2333] = 1'b0;  wr_cycle[ 2333] = 1'b1;  addr_rom[ 2333]='h00002474;  wr_data_rom[ 2333]='h0000148b;
    rd_cycle[ 2334] = 1'b0;  wr_cycle[ 2334] = 1'b1;  addr_rom[ 2334]='h00002478;  wr_data_rom[ 2334]='h000015fd;
    rd_cycle[ 2335] = 1'b0;  wr_cycle[ 2335] = 1'b1;  addr_rom[ 2335]='h0000247c;  wr_data_rom[ 2335]='h00003156;
    rd_cycle[ 2336] = 1'b0;  wr_cycle[ 2336] = 1'b1;  addr_rom[ 2336]='h00002480;  wr_data_rom[ 2336]='h00000083;
    rd_cycle[ 2337] = 1'b0;  wr_cycle[ 2337] = 1'b1;  addr_rom[ 2337]='h00002484;  wr_data_rom[ 2337]='h00002b0b;
    rd_cycle[ 2338] = 1'b0;  wr_cycle[ 2338] = 1'b1;  addr_rom[ 2338]='h00002488;  wr_data_rom[ 2338]='h00000485;
    rd_cycle[ 2339] = 1'b0;  wr_cycle[ 2339] = 1'b1;  addr_rom[ 2339]='h0000248c;  wr_data_rom[ 2339]='h00002da1;
    rd_cycle[ 2340] = 1'b0;  wr_cycle[ 2340] = 1'b1;  addr_rom[ 2340]='h00002490;  wr_data_rom[ 2340]='h00000796;
    rd_cycle[ 2341] = 1'b0;  wr_cycle[ 2341] = 1'b1;  addr_rom[ 2341]='h00002494;  wr_data_rom[ 2341]='h00003473;
    rd_cycle[ 2342] = 1'b0;  wr_cycle[ 2342] = 1'b1;  addr_rom[ 2342]='h00002498;  wr_data_rom[ 2342]='h00003e80;
    rd_cycle[ 2343] = 1'b0;  wr_cycle[ 2343] = 1'b1;  addr_rom[ 2343]='h0000249c;  wr_data_rom[ 2343]='h000030df;
    rd_cycle[ 2344] = 1'b0;  wr_cycle[ 2344] = 1'b1;  addr_rom[ 2344]='h000024a0;  wr_data_rom[ 2344]='h0000036d;
    rd_cycle[ 2345] = 1'b0;  wr_cycle[ 2345] = 1'b1;  addr_rom[ 2345]='h000024a4;  wr_data_rom[ 2345]='h0000223e;
    rd_cycle[ 2346] = 1'b0;  wr_cycle[ 2346] = 1'b1;  addr_rom[ 2346]='h000024a8;  wr_data_rom[ 2346]='h0000162a;
    rd_cycle[ 2347] = 1'b0;  wr_cycle[ 2347] = 1'b1;  addr_rom[ 2347]='h000024ac;  wr_data_rom[ 2347]='h00002b21;
    rd_cycle[ 2348] = 1'b0;  wr_cycle[ 2348] = 1'b1;  addr_rom[ 2348]='h000024b0;  wr_data_rom[ 2348]='h000005f4;
    rd_cycle[ 2349] = 1'b0;  wr_cycle[ 2349] = 1'b1;  addr_rom[ 2349]='h000024b4;  wr_data_rom[ 2349]='h00001d8e;
    rd_cycle[ 2350] = 1'b0;  wr_cycle[ 2350] = 1'b1;  addr_rom[ 2350]='h000024b8;  wr_data_rom[ 2350]='h00000c0f;
    rd_cycle[ 2351] = 1'b0;  wr_cycle[ 2351] = 1'b1;  addr_rom[ 2351]='h000024bc;  wr_data_rom[ 2351]='h0000076a;
    rd_cycle[ 2352] = 1'b0;  wr_cycle[ 2352] = 1'b1;  addr_rom[ 2352]='h000024c0;  wr_data_rom[ 2352]='h000039f8;
    rd_cycle[ 2353] = 1'b0;  wr_cycle[ 2353] = 1'b1;  addr_rom[ 2353]='h000024c4;  wr_data_rom[ 2353]='h00000ec0;
    rd_cycle[ 2354] = 1'b0;  wr_cycle[ 2354] = 1'b1;  addr_rom[ 2354]='h000024c8;  wr_data_rom[ 2354]='h00003550;
    rd_cycle[ 2355] = 1'b0;  wr_cycle[ 2355] = 1'b1;  addr_rom[ 2355]='h000024cc;  wr_data_rom[ 2355]='h0000006d;
    rd_cycle[ 2356] = 1'b0;  wr_cycle[ 2356] = 1'b1;  addr_rom[ 2356]='h000024d0;  wr_data_rom[ 2356]='h00000cd6;
    rd_cycle[ 2357] = 1'b0;  wr_cycle[ 2357] = 1'b1;  addr_rom[ 2357]='h000024d4;  wr_data_rom[ 2357]='h000009c8;
    rd_cycle[ 2358] = 1'b0;  wr_cycle[ 2358] = 1'b1;  addr_rom[ 2358]='h000024d8;  wr_data_rom[ 2358]='h00000df2;
    rd_cycle[ 2359] = 1'b0;  wr_cycle[ 2359] = 1'b1;  addr_rom[ 2359]='h000024dc;  wr_data_rom[ 2359]='h0000196f;
    rd_cycle[ 2360] = 1'b0;  wr_cycle[ 2360] = 1'b1;  addr_rom[ 2360]='h000024e0;  wr_data_rom[ 2360]='h00001260;
    rd_cycle[ 2361] = 1'b0;  wr_cycle[ 2361] = 1'b1;  addr_rom[ 2361]='h000024e4;  wr_data_rom[ 2361]='h0000252a;
    rd_cycle[ 2362] = 1'b0;  wr_cycle[ 2362] = 1'b1;  addr_rom[ 2362]='h000024e8;  wr_data_rom[ 2362]='h000029fa;
    rd_cycle[ 2363] = 1'b0;  wr_cycle[ 2363] = 1'b1;  addr_rom[ 2363]='h000024ec;  wr_data_rom[ 2363]='h00001c4a;
    rd_cycle[ 2364] = 1'b0;  wr_cycle[ 2364] = 1'b1;  addr_rom[ 2364]='h000024f0;  wr_data_rom[ 2364]='h00003e4f;
    rd_cycle[ 2365] = 1'b0;  wr_cycle[ 2365] = 1'b1;  addr_rom[ 2365]='h000024f4;  wr_data_rom[ 2365]='h0000062b;
    rd_cycle[ 2366] = 1'b0;  wr_cycle[ 2366] = 1'b1;  addr_rom[ 2366]='h000024f8;  wr_data_rom[ 2366]='h00002968;
    rd_cycle[ 2367] = 1'b0;  wr_cycle[ 2367] = 1'b1;  addr_rom[ 2367]='h000024fc;  wr_data_rom[ 2367]='h00000c84;
    rd_cycle[ 2368] = 1'b0;  wr_cycle[ 2368] = 1'b1;  addr_rom[ 2368]='h00002500;  wr_data_rom[ 2368]='h00000f36;
    rd_cycle[ 2369] = 1'b0;  wr_cycle[ 2369] = 1'b1;  addr_rom[ 2369]='h00002504;  wr_data_rom[ 2369]='h00003d7d;
    rd_cycle[ 2370] = 1'b0;  wr_cycle[ 2370] = 1'b1;  addr_rom[ 2370]='h00002508;  wr_data_rom[ 2370]='h00000d42;
    rd_cycle[ 2371] = 1'b0;  wr_cycle[ 2371] = 1'b1;  addr_rom[ 2371]='h0000250c;  wr_data_rom[ 2371]='h00002b34;
    rd_cycle[ 2372] = 1'b0;  wr_cycle[ 2372] = 1'b1;  addr_rom[ 2372]='h00002510;  wr_data_rom[ 2372]='h00002bc2;
    rd_cycle[ 2373] = 1'b0;  wr_cycle[ 2373] = 1'b1;  addr_rom[ 2373]='h00002514;  wr_data_rom[ 2373]='h00001454;
    rd_cycle[ 2374] = 1'b0;  wr_cycle[ 2374] = 1'b1;  addr_rom[ 2374]='h00002518;  wr_data_rom[ 2374]='h000017eb;
    rd_cycle[ 2375] = 1'b0;  wr_cycle[ 2375] = 1'b1;  addr_rom[ 2375]='h0000251c;  wr_data_rom[ 2375]='h00002558;
    rd_cycle[ 2376] = 1'b0;  wr_cycle[ 2376] = 1'b1;  addr_rom[ 2376]='h00002520;  wr_data_rom[ 2376]='h00001ccc;
    rd_cycle[ 2377] = 1'b0;  wr_cycle[ 2377] = 1'b1;  addr_rom[ 2377]='h00002524;  wr_data_rom[ 2377]='h00001737;
    rd_cycle[ 2378] = 1'b0;  wr_cycle[ 2378] = 1'b1;  addr_rom[ 2378]='h00002528;  wr_data_rom[ 2378]='h00001412;
    rd_cycle[ 2379] = 1'b0;  wr_cycle[ 2379] = 1'b1;  addr_rom[ 2379]='h0000252c;  wr_data_rom[ 2379]='h00001e4e;
    rd_cycle[ 2380] = 1'b0;  wr_cycle[ 2380] = 1'b1;  addr_rom[ 2380]='h00002530;  wr_data_rom[ 2380]='h00000805;
    rd_cycle[ 2381] = 1'b0;  wr_cycle[ 2381] = 1'b1;  addr_rom[ 2381]='h00002534;  wr_data_rom[ 2381]='h000013a1;
    rd_cycle[ 2382] = 1'b0;  wr_cycle[ 2382] = 1'b1;  addr_rom[ 2382]='h00002538;  wr_data_rom[ 2382]='h00003efb;
    rd_cycle[ 2383] = 1'b0;  wr_cycle[ 2383] = 1'b1;  addr_rom[ 2383]='h0000253c;  wr_data_rom[ 2383]='h00001d21;
    rd_cycle[ 2384] = 1'b0;  wr_cycle[ 2384] = 1'b1;  addr_rom[ 2384]='h00002540;  wr_data_rom[ 2384]='h000019ee;
    rd_cycle[ 2385] = 1'b0;  wr_cycle[ 2385] = 1'b1;  addr_rom[ 2385]='h00002544;  wr_data_rom[ 2385]='h000005e5;
    rd_cycle[ 2386] = 1'b0;  wr_cycle[ 2386] = 1'b1;  addr_rom[ 2386]='h00002548;  wr_data_rom[ 2386]='h00002d8f;
    rd_cycle[ 2387] = 1'b0;  wr_cycle[ 2387] = 1'b1;  addr_rom[ 2387]='h0000254c;  wr_data_rom[ 2387]='h000038c5;
    rd_cycle[ 2388] = 1'b0;  wr_cycle[ 2388] = 1'b1;  addr_rom[ 2388]='h00002550;  wr_data_rom[ 2388]='h000003d9;
    rd_cycle[ 2389] = 1'b0;  wr_cycle[ 2389] = 1'b1;  addr_rom[ 2389]='h00002554;  wr_data_rom[ 2389]='h000021e4;
    rd_cycle[ 2390] = 1'b0;  wr_cycle[ 2390] = 1'b1;  addr_rom[ 2390]='h00002558;  wr_data_rom[ 2390]='h0000291a;
    rd_cycle[ 2391] = 1'b0;  wr_cycle[ 2391] = 1'b1;  addr_rom[ 2391]='h0000255c;  wr_data_rom[ 2391]='h00001969;
    rd_cycle[ 2392] = 1'b0;  wr_cycle[ 2392] = 1'b1;  addr_rom[ 2392]='h00002560;  wr_data_rom[ 2392]='h00001536;
    rd_cycle[ 2393] = 1'b0;  wr_cycle[ 2393] = 1'b1;  addr_rom[ 2393]='h00002564;  wr_data_rom[ 2393]='h0000233f;
    rd_cycle[ 2394] = 1'b0;  wr_cycle[ 2394] = 1'b1;  addr_rom[ 2394]='h00002568;  wr_data_rom[ 2394]='h00003045;
    rd_cycle[ 2395] = 1'b0;  wr_cycle[ 2395] = 1'b1;  addr_rom[ 2395]='h0000256c;  wr_data_rom[ 2395]='h0000394f;
    rd_cycle[ 2396] = 1'b0;  wr_cycle[ 2396] = 1'b1;  addr_rom[ 2396]='h00002570;  wr_data_rom[ 2396]='h00002c59;
    rd_cycle[ 2397] = 1'b0;  wr_cycle[ 2397] = 1'b1;  addr_rom[ 2397]='h00002574;  wr_data_rom[ 2397]='h00001276;
    rd_cycle[ 2398] = 1'b0;  wr_cycle[ 2398] = 1'b1;  addr_rom[ 2398]='h00002578;  wr_data_rom[ 2398]='h00000681;
    rd_cycle[ 2399] = 1'b0;  wr_cycle[ 2399] = 1'b1;  addr_rom[ 2399]='h0000257c;  wr_data_rom[ 2399]='h00002902;
    rd_cycle[ 2400] = 1'b0;  wr_cycle[ 2400] = 1'b1;  addr_rom[ 2400]='h00002580;  wr_data_rom[ 2400]='h00003426;
    rd_cycle[ 2401] = 1'b0;  wr_cycle[ 2401] = 1'b1;  addr_rom[ 2401]='h00002584;  wr_data_rom[ 2401]='h000005fd;
    rd_cycle[ 2402] = 1'b0;  wr_cycle[ 2402] = 1'b1;  addr_rom[ 2402]='h00002588;  wr_data_rom[ 2402]='h000018b4;
    rd_cycle[ 2403] = 1'b0;  wr_cycle[ 2403] = 1'b1;  addr_rom[ 2403]='h0000258c;  wr_data_rom[ 2403]='h00003971;
    rd_cycle[ 2404] = 1'b0;  wr_cycle[ 2404] = 1'b1;  addr_rom[ 2404]='h00002590;  wr_data_rom[ 2404]='h000024b7;
    rd_cycle[ 2405] = 1'b0;  wr_cycle[ 2405] = 1'b1;  addr_rom[ 2405]='h00002594;  wr_data_rom[ 2405]='h00001579;
    rd_cycle[ 2406] = 1'b0;  wr_cycle[ 2406] = 1'b1;  addr_rom[ 2406]='h00002598;  wr_data_rom[ 2406]='h00001d1d;
    rd_cycle[ 2407] = 1'b0;  wr_cycle[ 2407] = 1'b1;  addr_rom[ 2407]='h0000259c;  wr_data_rom[ 2407]='h00001187;
    rd_cycle[ 2408] = 1'b0;  wr_cycle[ 2408] = 1'b1;  addr_rom[ 2408]='h000025a0;  wr_data_rom[ 2408]='h00003bfc;
    rd_cycle[ 2409] = 1'b0;  wr_cycle[ 2409] = 1'b1;  addr_rom[ 2409]='h000025a4;  wr_data_rom[ 2409]='h0000130f;
    rd_cycle[ 2410] = 1'b0;  wr_cycle[ 2410] = 1'b1;  addr_rom[ 2410]='h000025a8;  wr_data_rom[ 2410]='h000005fa;
    rd_cycle[ 2411] = 1'b0;  wr_cycle[ 2411] = 1'b1;  addr_rom[ 2411]='h000025ac;  wr_data_rom[ 2411]='h00001a57;
    rd_cycle[ 2412] = 1'b0;  wr_cycle[ 2412] = 1'b1;  addr_rom[ 2412]='h000025b0;  wr_data_rom[ 2412]='h00001f80;
    rd_cycle[ 2413] = 1'b0;  wr_cycle[ 2413] = 1'b1;  addr_rom[ 2413]='h000025b4;  wr_data_rom[ 2413]='h00002357;
    rd_cycle[ 2414] = 1'b0;  wr_cycle[ 2414] = 1'b1;  addr_rom[ 2414]='h000025b8;  wr_data_rom[ 2414]='h00002f76;
    rd_cycle[ 2415] = 1'b0;  wr_cycle[ 2415] = 1'b1;  addr_rom[ 2415]='h000025bc;  wr_data_rom[ 2415]='h00001bea;
    rd_cycle[ 2416] = 1'b0;  wr_cycle[ 2416] = 1'b1;  addr_rom[ 2416]='h000025c0;  wr_data_rom[ 2416]='h0000187c;
    rd_cycle[ 2417] = 1'b0;  wr_cycle[ 2417] = 1'b1;  addr_rom[ 2417]='h000025c4;  wr_data_rom[ 2417]='h00003bc7;
    rd_cycle[ 2418] = 1'b0;  wr_cycle[ 2418] = 1'b1;  addr_rom[ 2418]='h000025c8;  wr_data_rom[ 2418]='h0000202e;
    rd_cycle[ 2419] = 1'b0;  wr_cycle[ 2419] = 1'b1;  addr_rom[ 2419]='h000025cc;  wr_data_rom[ 2419]='h00003507;
    rd_cycle[ 2420] = 1'b0;  wr_cycle[ 2420] = 1'b1;  addr_rom[ 2420]='h000025d0;  wr_data_rom[ 2420]='h00002420;
    rd_cycle[ 2421] = 1'b0;  wr_cycle[ 2421] = 1'b1;  addr_rom[ 2421]='h000025d4;  wr_data_rom[ 2421]='h00002595;
    rd_cycle[ 2422] = 1'b0;  wr_cycle[ 2422] = 1'b1;  addr_rom[ 2422]='h000025d8;  wr_data_rom[ 2422]='h000022fe;
    rd_cycle[ 2423] = 1'b0;  wr_cycle[ 2423] = 1'b1;  addr_rom[ 2423]='h000025dc;  wr_data_rom[ 2423]='h00001d98;
    rd_cycle[ 2424] = 1'b0;  wr_cycle[ 2424] = 1'b1;  addr_rom[ 2424]='h000025e0;  wr_data_rom[ 2424]='h00001374;
    rd_cycle[ 2425] = 1'b0;  wr_cycle[ 2425] = 1'b1;  addr_rom[ 2425]='h000025e4;  wr_data_rom[ 2425]='h00002db8;
    rd_cycle[ 2426] = 1'b0;  wr_cycle[ 2426] = 1'b1;  addr_rom[ 2426]='h000025e8;  wr_data_rom[ 2426]='h0000166a;
    rd_cycle[ 2427] = 1'b0;  wr_cycle[ 2427] = 1'b1;  addr_rom[ 2427]='h000025ec;  wr_data_rom[ 2427]='h000006ac;
    rd_cycle[ 2428] = 1'b0;  wr_cycle[ 2428] = 1'b1;  addr_rom[ 2428]='h000025f0;  wr_data_rom[ 2428]='h00003a9f;
    rd_cycle[ 2429] = 1'b0;  wr_cycle[ 2429] = 1'b1;  addr_rom[ 2429]='h000025f4;  wr_data_rom[ 2429]='h000035d0;
    rd_cycle[ 2430] = 1'b0;  wr_cycle[ 2430] = 1'b1;  addr_rom[ 2430]='h000025f8;  wr_data_rom[ 2430]='h000023b5;
    rd_cycle[ 2431] = 1'b0;  wr_cycle[ 2431] = 1'b1;  addr_rom[ 2431]='h000025fc;  wr_data_rom[ 2431]='h0000170e;
    rd_cycle[ 2432] = 1'b0;  wr_cycle[ 2432] = 1'b1;  addr_rom[ 2432]='h00002600;  wr_data_rom[ 2432]='h0000354b;
    rd_cycle[ 2433] = 1'b0;  wr_cycle[ 2433] = 1'b1;  addr_rom[ 2433]='h00002604;  wr_data_rom[ 2433]='h00001b21;
    rd_cycle[ 2434] = 1'b0;  wr_cycle[ 2434] = 1'b1;  addr_rom[ 2434]='h00002608;  wr_data_rom[ 2434]='h00000f41;
    rd_cycle[ 2435] = 1'b0;  wr_cycle[ 2435] = 1'b1;  addr_rom[ 2435]='h0000260c;  wr_data_rom[ 2435]='h000016a5;
    rd_cycle[ 2436] = 1'b0;  wr_cycle[ 2436] = 1'b1;  addr_rom[ 2436]='h00002610;  wr_data_rom[ 2436]='h00000c02;
    rd_cycle[ 2437] = 1'b0;  wr_cycle[ 2437] = 1'b1;  addr_rom[ 2437]='h00002614;  wr_data_rom[ 2437]='h00003895;
    rd_cycle[ 2438] = 1'b0;  wr_cycle[ 2438] = 1'b1;  addr_rom[ 2438]='h00002618;  wr_data_rom[ 2438]='h00003b22;
    rd_cycle[ 2439] = 1'b0;  wr_cycle[ 2439] = 1'b1;  addr_rom[ 2439]='h0000261c;  wr_data_rom[ 2439]='h00001a07;
    rd_cycle[ 2440] = 1'b0;  wr_cycle[ 2440] = 1'b1;  addr_rom[ 2440]='h00002620;  wr_data_rom[ 2440]='h0000115a;
    rd_cycle[ 2441] = 1'b0;  wr_cycle[ 2441] = 1'b1;  addr_rom[ 2441]='h00002624;  wr_data_rom[ 2441]='h00003060;
    rd_cycle[ 2442] = 1'b0;  wr_cycle[ 2442] = 1'b1;  addr_rom[ 2442]='h00002628;  wr_data_rom[ 2442]='h000022e5;
    rd_cycle[ 2443] = 1'b0;  wr_cycle[ 2443] = 1'b1;  addr_rom[ 2443]='h0000262c;  wr_data_rom[ 2443]='h00003465;
    rd_cycle[ 2444] = 1'b0;  wr_cycle[ 2444] = 1'b1;  addr_rom[ 2444]='h00002630;  wr_data_rom[ 2444]='h00002142;
    rd_cycle[ 2445] = 1'b0;  wr_cycle[ 2445] = 1'b1;  addr_rom[ 2445]='h00002634;  wr_data_rom[ 2445]='h000009d5;
    rd_cycle[ 2446] = 1'b0;  wr_cycle[ 2446] = 1'b1;  addr_rom[ 2446]='h00002638;  wr_data_rom[ 2446]='h00002ef2;
    rd_cycle[ 2447] = 1'b0;  wr_cycle[ 2447] = 1'b1;  addr_rom[ 2447]='h0000263c;  wr_data_rom[ 2447]='h00002a5b;
    rd_cycle[ 2448] = 1'b0;  wr_cycle[ 2448] = 1'b1;  addr_rom[ 2448]='h00002640;  wr_data_rom[ 2448]='h000010f9;
    rd_cycle[ 2449] = 1'b0;  wr_cycle[ 2449] = 1'b1;  addr_rom[ 2449]='h00002644;  wr_data_rom[ 2449]='h00002d9e;
    rd_cycle[ 2450] = 1'b0;  wr_cycle[ 2450] = 1'b1;  addr_rom[ 2450]='h00002648;  wr_data_rom[ 2450]='h000038f8;
    rd_cycle[ 2451] = 1'b0;  wr_cycle[ 2451] = 1'b1;  addr_rom[ 2451]='h0000264c;  wr_data_rom[ 2451]='h00003b5a;
    rd_cycle[ 2452] = 1'b0;  wr_cycle[ 2452] = 1'b1;  addr_rom[ 2452]='h00002650;  wr_data_rom[ 2452]='h00001b38;
    rd_cycle[ 2453] = 1'b0;  wr_cycle[ 2453] = 1'b1;  addr_rom[ 2453]='h00002654;  wr_data_rom[ 2453]='h00001a13;
    rd_cycle[ 2454] = 1'b0;  wr_cycle[ 2454] = 1'b1;  addr_rom[ 2454]='h00002658;  wr_data_rom[ 2454]='h000027ca;
    rd_cycle[ 2455] = 1'b0;  wr_cycle[ 2455] = 1'b1;  addr_rom[ 2455]='h0000265c;  wr_data_rom[ 2455]='h00002a5a;
    rd_cycle[ 2456] = 1'b0;  wr_cycle[ 2456] = 1'b1;  addr_rom[ 2456]='h00002660;  wr_data_rom[ 2456]='h0000057a;
    rd_cycle[ 2457] = 1'b0;  wr_cycle[ 2457] = 1'b1;  addr_rom[ 2457]='h00002664;  wr_data_rom[ 2457]='h00001b9b;
    rd_cycle[ 2458] = 1'b0;  wr_cycle[ 2458] = 1'b1;  addr_rom[ 2458]='h00002668;  wr_data_rom[ 2458]='h00000dc3;
    rd_cycle[ 2459] = 1'b0;  wr_cycle[ 2459] = 1'b1;  addr_rom[ 2459]='h0000266c;  wr_data_rom[ 2459]='h000030c8;
    rd_cycle[ 2460] = 1'b0;  wr_cycle[ 2460] = 1'b1;  addr_rom[ 2460]='h00002670;  wr_data_rom[ 2460]='h00003d06;
    rd_cycle[ 2461] = 1'b0;  wr_cycle[ 2461] = 1'b1;  addr_rom[ 2461]='h00002674;  wr_data_rom[ 2461]='h0000030b;
    rd_cycle[ 2462] = 1'b0;  wr_cycle[ 2462] = 1'b1;  addr_rom[ 2462]='h00002678;  wr_data_rom[ 2462]='h00002b6a;
    rd_cycle[ 2463] = 1'b0;  wr_cycle[ 2463] = 1'b1;  addr_rom[ 2463]='h0000267c;  wr_data_rom[ 2463]='h00002720;
    rd_cycle[ 2464] = 1'b0;  wr_cycle[ 2464] = 1'b1;  addr_rom[ 2464]='h00002680;  wr_data_rom[ 2464]='h00003215;
    rd_cycle[ 2465] = 1'b0;  wr_cycle[ 2465] = 1'b1;  addr_rom[ 2465]='h00002684;  wr_data_rom[ 2465]='h00001aed;
    rd_cycle[ 2466] = 1'b0;  wr_cycle[ 2466] = 1'b1;  addr_rom[ 2466]='h00002688;  wr_data_rom[ 2466]='h000038b7;
    rd_cycle[ 2467] = 1'b0;  wr_cycle[ 2467] = 1'b1;  addr_rom[ 2467]='h0000268c;  wr_data_rom[ 2467]='h000001be;
    rd_cycle[ 2468] = 1'b0;  wr_cycle[ 2468] = 1'b1;  addr_rom[ 2468]='h00002690;  wr_data_rom[ 2468]='h0000111b;
    rd_cycle[ 2469] = 1'b0;  wr_cycle[ 2469] = 1'b1;  addr_rom[ 2469]='h00002694;  wr_data_rom[ 2469]='h00003efb;
    rd_cycle[ 2470] = 1'b0;  wr_cycle[ 2470] = 1'b1;  addr_rom[ 2470]='h00002698;  wr_data_rom[ 2470]='h000010c5;
    rd_cycle[ 2471] = 1'b0;  wr_cycle[ 2471] = 1'b1;  addr_rom[ 2471]='h0000269c;  wr_data_rom[ 2471]='h00001b1b;
    rd_cycle[ 2472] = 1'b0;  wr_cycle[ 2472] = 1'b1;  addr_rom[ 2472]='h000026a0;  wr_data_rom[ 2472]='h00001c95;
    rd_cycle[ 2473] = 1'b0;  wr_cycle[ 2473] = 1'b1;  addr_rom[ 2473]='h000026a4;  wr_data_rom[ 2473]='h0000280f;
    rd_cycle[ 2474] = 1'b0;  wr_cycle[ 2474] = 1'b1;  addr_rom[ 2474]='h000026a8;  wr_data_rom[ 2474]='h00001ee6;
    rd_cycle[ 2475] = 1'b0;  wr_cycle[ 2475] = 1'b1;  addr_rom[ 2475]='h000026ac;  wr_data_rom[ 2475]='h00001074;
    rd_cycle[ 2476] = 1'b0;  wr_cycle[ 2476] = 1'b1;  addr_rom[ 2476]='h000026b0;  wr_data_rom[ 2476]='h0000018b;
    rd_cycle[ 2477] = 1'b0;  wr_cycle[ 2477] = 1'b1;  addr_rom[ 2477]='h000026b4;  wr_data_rom[ 2477]='h000027dc;
    rd_cycle[ 2478] = 1'b0;  wr_cycle[ 2478] = 1'b1;  addr_rom[ 2478]='h000026b8;  wr_data_rom[ 2478]='h00003bdd;
    rd_cycle[ 2479] = 1'b0;  wr_cycle[ 2479] = 1'b1;  addr_rom[ 2479]='h000026bc;  wr_data_rom[ 2479]='h00002abb;
    rd_cycle[ 2480] = 1'b0;  wr_cycle[ 2480] = 1'b1;  addr_rom[ 2480]='h000026c0;  wr_data_rom[ 2480]='h00000d40;
    rd_cycle[ 2481] = 1'b0;  wr_cycle[ 2481] = 1'b1;  addr_rom[ 2481]='h000026c4;  wr_data_rom[ 2481]='h00003199;
    rd_cycle[ 2482] = 1'b0;  wr_cycle[ 2482] = 1'b1;  addr_rom[ 2482]='h000026c8;  wr_data_rom[ 2482]='h000006dc;
    rd_cycle[ 2483] = 1'b0;  wr_cycle[ 2483] = 1'b1;  addr_rom[ 2483]='h000026cc;  wr_data_rom[ 2483]='h000023ff;
    rd_cycle[ 2484] = 1'b0;  wr_cycle[ 2484] = 1'b1;  addr_rom[ 2484]='h000026d0;  wr_data_rom[ 2484]='h000032ae;
    rd_cycle[ 2485] = 1'b0;  wr_cycle[ 2485] = 1'b1;  addr_rom[ 2485]='h000026d4;  wr_data_rom[ 2485]='h000003f8;
    rd_cycle[ 2486] = 1'b0;  wr_cycle[ 2486] = 1'b1;  addr_rom[ 2486]='h000026d8;  wr_data_rom[ 2486]='h000030eb;
    rd_cycle[ 2487] = 1'b0;  wr_cycle[ 2487] = 1'b1;  addr_rom[ 2487]='h000026dc;  wr_data_rom[ 2487]='h000014b6;
    rd_cycle[ 2488] = 1'b0;  wr_cycle[ 2488] = 1'b1;  addr_rom[ 2488]='h000026e0;  wr_data_rom[ 2488]='h00003516;
    rd_cycle[ 2489] = 1'b0;  wr_cycle[ 2489] = 1'b1;  addr_rom[ 2489]='h000026e4;  wr_data_rom[ 2489]='h00002560;
    rd_cycle[ 2490] = 1'b0;  wr_cycle[ 2490] = 1'b1;  addr_rom[ 2490]='h000026e8;  wr_data_rom[ 2490]='h00003fc1;
    rd_cycle[ 2491] = 1'b0;  wr_cycle[ 2491] = 1'b1;  addr_rom[ 2491]='h000026ec;  wr_data_rom[ 2491]='h000019f9;
    rd_cycle[ 2492] = 1'b0;  wr_cycle[ 2492] = 1'b1;  addr_rom[ 2492]='h000026f0;  wr_data_rom[ 2492]='h00001d49;
    rd_cycle[ 2493] = 1'b0;  wr_cycle[ 2493] = 1'b1;  addr_rom[ 2493]='h000026f4;  wr_data_rom[ 2493]='h00003bf9;
    rd_cycle[ 2494] = 1'b0;  wr_cycle[ 2494] = 1'b1;  addr_rom[ 2494]='h000026f8;  wr_data_rom[ 2494]='h00000c0a;
    rd_cycle[ 2495] = 1'b0;  wr_cycle[ 2495] = 1'b1;  addr_rom[ 2495]='h000026fc;  wr_data_rom[ 2495]='h00003193;
    rd_cycle[ 2496] = 1'b0;  wr_cycle[ 2496] = 1'b1;  addr_rom[ 2496]='h00002700;  wr_data_rom[ 2496]='h00003f9a;
    rd_cycle[ 2497] = 1'b0;  wr_cycle[ 2497] = 1'b1;  addr_rom[ 2497]='h00002704;  wr_data_rom[ 2497]='h00002e15;
    rd_cycle[ 2498] = 1'b0;  wr_cycle[ 2498] = 1'b1;  addr_rom[ 2498]='h00002708;  wr_data_rom[ 2498]='h00001e42;
    rd_cycle[ 2499] = 1'b0;  wr_cycle[ 2499] = 1'b1;  addr_rom[ 2499]='h0000270c;  wr_data_rom[ 2499]='h00000167;
    rd_cycle[ 2500] = 1'b0;  wr_cycle[ 2500] = 1'b1;  addr_rom[ 2500]='h00002710;  wr_data_rom[ 2500]='h000039bf;
    rd_cycle[ 2501] = 1'b0;  wr_cycle[ 2501] = 1'b1;  addr_rom[ 2501]='h00002714;  wr_data_rom[ 2501]='h00000ab4;
    rd_cycle[ 2502] = 1'b0;  wr_cycle[ 2502] = 1'b1;  addr_rom[ 2502]='h00002718;  wr_data_rom[ 2502]='h000032f7;
    rd_cycle[ 2503] = 1'b0;  wr_cycle[ 2503] = 1'b1;  addr_rom[ 2503]='h0000271c;  wr_data_rom[ 2503]='h00000005;
    rd_cycle[ 2504] = 1'b0;  wr_cycle[ 2504] = 1'b1;  addr_rom[ 2504]='h00002720;  wr_data_rom[ 2504]='h00002f0d;
    rd_cycle[ 2505] = 1'b0;  wr_cycle[ 2505] = 1'b1;  addr_rom[ 2505]='h00002724;  wr_data_rom[ 2505]='h00003a0f;
    rd_cycle[ 2506] = 1'b0;  wr_cycle[ 2506] = 1'b1;  addr_rom[ 2506]='h00002728;  wr_data_rom[ 2506]='h00000130;
    rd_cycle[ 2507] = 1'b0;  wr_cycle[ 2507] = 1'b1;  addr_rom[ 2507]='h0000272c;  wr_data_rom[ 2507]='h000035b4;
    rd_cycle[ 2508] = 1'b0;  wr_cycle[ 2508] = 1'b1;  addr_rom[ 2508]='h00002730;  wr_data_rom[ 2508]='h00001862;
    rd_cycle[ 2509] = 1'b0;  wr_cycle[ 2509] = 1'b1;  addr_rom[ 2509]='h00002734;  wr_data_rom[ 2509]='h00003874;
    rd_cycle[ 2510] = 1'b0;  wr_cycle[ 2510] = 1'b1;  addr_rom[ 2510]='h00002738;  wr_data_rom[ 2510]='h0000064c;
    rd_cycle[ 2511] = 1'b0;  wr_cycle[ 2511] = 1'b1;  addr_rom[ 2511]='h0000273c;  wr_data_rom[ 2511]='h000037b0;
    rd_cycle[ 2512] = 1'b0;  wr_cycle[ 2512] = 1'b1;  addr_rom[ 2512]='h00002740;  wr_data_rom[ 2512]='h00002488;
    rd_cycle[ 2513] = 1'b0;  wr_cycle[ 2513] = 1'b1;  addr_rom[ 2513]='h00002744;  wr_data_rom[ 2513]='h000028cb;
    rd_cycle[ 2514] = 1'b0;  wr_cycle[ 2514] = 1'b1;  addr_rom[ 2514]='h00002748;  wr_data_rom[ 2514]='h00001419;
    rd_cycle[ 2515] = 1'b0;  wr_cycle[ 2515] = 1'b1;  addr_rom[ 2515]='h0000274c;  wr_data_rom[ 2515]='h000016eb;
    rd_cycle[ 2516] = 1'b0;  wr_cycle[ 2516] = 1'b1;  addr_rom[ 2516]='h00002750;  wr_data_rom[ 2516]='h0000356c;
    rd_cycle[ 2517] = 1'b0;  wr_cycle[ 2517] = 1'b1;  addr_rom[ 2517]='h00002754;  wr_data_rom[ 2517]='h0000360e;
    rd_cycle[ 2518] = 1'b0;  wr_cycle[ 2518] = 1'b1;  addr_rom[ 2518]='h00002758;  wr_data_rom[ 2518]='h00001294;
    rd_cycle[ 2519] = 1'b0;  wr_cycle[ 2519] = 1'b1;  addr_rom[ 2519]='h0000275c;  wr_data_rom[ 2519]='h00003c8e;
    rd_cycle[ 2520] = 1'b0;  wr_cycle[ 2520] = 1'b1;  addr_rom[ 2520]='h00002760;  wr_data_rom[ 2520]='h000008b3;
    rd_cycle[ 2521] = 1'b0;  wr_cycle[ 2521] = 1'b1;  addr_rom[ 2521]='h00002764;  wr_data_rom[ 2521]='h00002ec0;
    rd_cycle[ 2522] = 1'b0;  wr_cycle[ 2522] = 1'b1;  addr_rom[ 2522]='h00002768;  wr_data_rom[ 2522]='h000009d8;
    rd_cycle[ 2523] = 1'b0;  wr_cycle[ 2523] = 1'b1;  addr_rom[ 2523]='h0000276c;  wr_data_rom[ 2523]='h000034d6;
    rd_cycle[ 2524] = 1'b0;  wr_cycle[ 2524] = 1'b1;  addr_rom[ 2524]='h00002770;  wr_data_rom[ 2524]='h00003216;
    rd_cycle[ 2525] = 1'b0;  wr_cycle[ 2525] = 1'b1;  addr_rom[ 2525]='h00002774;  wr_data_rom[ 2525]='h00002e60;
    rd_cycle[ 2526] = 1'b0;  wr_cycle[ 2526] = 1'b1;  addr_rom[ 2526]='h00002778;  wr_data_rom[ 2526]='h0000053a;
    rd_cycle[ 2527] = 1'b0;  wr_cycle[ 2527] = 1'b1;  addr_rom[ 2527]='h0000277c;  wr_data_rom[ 2527]='h00002e9f;
    rd_cycle[ 2528] = 1'b0;  wr_cycle[ 2528] = 1'b1;  addr_rom[ 2528]='h00002780;  wr_data_rom[ 2528]='h00001a39;
    rd_cycle[ 2529] = 1'b0;  wr_cycle[ 2529] = 1'b1;  addr_rom[ 2529]='h00002784;  wr_data_rom[ 2529]='h00003118;
    rd_cycle[ 2530] = 1'b0;  wr_cycle[ 2530] = 1'b1;  addr_rom[ 2530]='h00002788;  wr_data_rom[ 2530]='h00003fb3;
    rd_cycle[ 2531] = 1'b0;  wr_cycle[ 2531] = 1'b1;  addr_rom[ 2531]='h0000278c;  wr_data_rom[ 2531]='h0000191d;
    rd_cycle[ 2532] = 1'b0;  wr_cycle[ 2532] = 1'b1;  addr_rom[ 2532]='h00002790;  wr_data_rom[ 2532]='h00001483;
    rd_cycle[ 2533] = 1'b0;  wr_cycle[ 2533] = 1'b1;  addr_rom[ 2533]='h00002794;  wr_data_rom[ 2533]='h000022e9;
    rd_cycle[ 2534] = 1'b0;  wr_cycle[ 2534] = 1'b1;  addr_rom[ 2534]='h00002798;  wr_data_rom[ 2534]='h00000a4d;
    rd_cycle[ 2535] = 1'b0;  wr_cycle[ 2535] = 1'b1;  addr_rom[ 2535]='h0000279c;  wr_data_rom[ 2535]='h00000cfa;
    rd_cycle[ 2536] = 1'b0;  wr_cycle[ 2536] = 1'b1;  addr_rom[ 2536]='h000027a0;  wr_data_rom[ 2536]='h000033fa;
    rd_cycle[ 2537] = 1'b0;  wr_cycle[ 2537] = 1'b1;  addr_rom[ 2537]='h000027a4;  wr_data_rom[ 2537]='h00003b8c;
    rd_cycle[ 2538] = 1'b0;  wr_cycle[ 2538] = 1'b1;  addr_rom[ 2538]='h000027a8;  wr_data_rom[ 2538]='h0000234c;
    rd_cycle[ 2539] = 1'b0;  wr_cycle[ 2539] = 1'b1;  addr_rom[ 2539]='h000027ac;  wr_data_rom[ 2539]='h000010ca;
    rd_cycle[ 2540] = 1'b0;  wr_cycle[ 2540] = 1'b1;  addr_rom[ 2540]='h000027b0;  wr_data_rom[ 2540]='h00001919;
    rd_cycle[ 2541] = 1'b0;  wr_cycle[ 2541] = 1'b1;  addr_rom[ 2541]='h000027b4;  wr_data_rom[ 2541]='h000037c8;
    rd_cycle[ 2542] = 1'b0;  wr_cycle[ 2542] = 1'b1;  addr_rom[ 2542]='h000027b8;  wr_data_rom[ 2542]='h00000b63;
    rd_cycle[ 2543] = 1'b0;  wr_cycle[ 2543] = 1'b1;  addr_rom[ 2543]='h000027bc;  wr_data_rom[ 2543]='h00001647;
    rd_cycle[ 2544] = 1'b0;  wr_cycle[ 2544] = 1'b1;  addr_rom[ 2544]='h000027c0;  wr_data_rom[ 2544]='h00003c64;
    rd_cycle[ 2545] = 1'b0;  wr_cycle[ 2545] = 1'b1;  addr_rom[ 2545]='h000027c4;  wr_data_rom[ 2545]='h00001756;
    rd_cycle[ 2546] = 1'b0;  wr_cycle[ 2546] = 1'b1;  addr_rom[ 2546]='h000027c8;  wr_data_rom[ 2546]='h00003cee;
    rd_cycle[ 2547] = 1'b0;  wr_cycle[ 2547] = 1'b1;  addr_rom[ 2547]='h000027cc;  wr_data_rom[ 2547]='h00001f52;
    rd_cycle[ 2548] = 1'b0;  wr_cycle[ 2548] = 1'b1;  addr_rom[ 2548]='h000027d0;  wr_data_rom[ 2548]='h000028b8;
    rd_cycle[ 2549] = 1'b0;  wr_cycle[ 2549] = 1'b1;  addr_rom[ 2549]='h000027d4;  wr_data_rom[ 2549]='h00002657;
    rd_cycle[ 2550] = 1'b0;  wr_cycle[ 2550] = 1'b1;  addr_rom[ 2550]='h000027d8;  wr_data_rom[ 2550]='h00000754;
    rd_cycle[ 2551] = 1'b0;  wr_cycle[ 2551] = 1'b1;  addr_rom[ 2551]='h000027dc;  wr_data_rom[ 2551]='h00002d58;
    rd_cycle[ 2552] = 1'b0;  wr_cycle[ 2552] = 1'b1;  addr_rom[ 2552]='h000027e0;  wr_data_rom[ 2552]='h000020c6;
    rd_cycle[ 2553] = 1'b0;  wr_cycle[ 2553] = 1'b1;  addr_rom[ 2553]='h000027e4;  wr_data_rom[ 2553]='h0000059d;
    rd_cycle[ 2554] = 1'b0;  wr_cycle[ 2554] = 1'b1;  addr_rom[ 2554]='h000027e8;  wr_data_rom[ 2554]='h00002762;
    rd_cycle[ 2555] = 1'b0;  wr_cycle[ 2555] = 1'b1;  addr_rom[ 2555]='h000027ec;  wr_data_rom[ 2555]='h000038cf;
    rd_cycle[ 2556] = 1'b0;  wr_cycle[ 2556] = 1'b1;  addr_rom[ 2556]='h000027f0;  wr_data_rom[ 2556]='h00001a85;
    rd_cycle[ 2557] = 1'b0;  wr_cycle[ 2557] = 1'b1;  addr_rom[ 2557]='h000027f4;  wr_data_rom[ 2557]='h00003fec;
    rd_cycle[ 2558] = 1'b0;  wr_cycle[ 2558] = 1'b1;  addr_rom[ 2558]='h000027f8;  wr_data_rom[ 2558]='h0000037a;
    rd_cycle[ 2559] = 1'b0;  wr_cycle[ 2559] = 1'b1;  addr_rom[ 2559]='h000027fc;  wr_data_rom[ 2559]='h00002ffa;
    rd_cycle[ 2560] = 1'b0;  wr_cycle[ 2560] = 1'b1;  addr_rom[ 2560]='h00002800;  wr_data_rom[ 2560]='h000012bd;
    rd_cycle[ 2561] = 1'b0;  wr_cycle[ 2561] = 1'b1;  addr_rom[ 2561]='h00002804;  wr_data_rom[ 2561]='h000012c5;
    rd_cycle[ 2562] = 1'b0;  wr_cycle[ 2562] = 1'b1;  addr_rom[ 2562]='h00002808;  wr_data_rom[ 2562]='h00003545;
    rd_cycle[ 2563] = 1'b0;  wr_cycle[ 2563] = 1'b1;  addr_rom[ 2563]='h0000280c;  wr_data_rom[ 2563]='h000020d1;
    rd_cycle[ 2564] = 1'b0;  wr_cycle[ 2564] = 1'b1;  addr_rom[ 2564]='h00002810;  wr_data_rom[ 2564]='h0000269a;
    rd_cycle[ 2565] = 1'b0;  wr_cycle[ 2565] = 1'b1;  addr_rom[ 2565]='h00002814;  wr_data_rom[ 2565]='h00001503;
    rd_cycle[ 2566] = 1'b0;  wr_cycle[ 2566] = 1'b1;  addr_rom[ 2566]='h00002818;  wr_data_rom[ 2566]='h00003587;
    rd_cycle[ 2567] = 1'b0;  wr_cycle[ 2567] = 1'b1;  addr_rom[ 2567]='h0000281c;  wr_data_rom[ 2567]='h00002f9e;
    rd_cycle[ 2568] = 1'b0;  wr_cycle[ 2568] = 1'b1;  addr_rom[ 2568]='h00002820;  wr_data_rom[ 2568]='h00003ec3;
    rd_cycle[ 2569] = 1'b0;  wr_cycle[ 2569] = 1'b1;  addr_rom[ 2569]='h00002824;  wr_data_rom[ 2569]='h000032ca;
    rd_cycle[ 2570] = 1'b0;  wr_cycle[ 2570] = 1'b1;  addr_rom[ 2570]='h00002828;  wr_data_rom[ 2570]='h00002fbc;
    rd_cycle[ 2571] = 1'b0;  wr_cycle[ 2571] = 1'b1;  addr_rom[ 2571]='h0000282c;  wr_data_rom[ 2571]='h00002172;
    rd_cycle[ 2572] = 1'b0;  wr_cycle[ 2572] = 1'b1;  addr_rom[ 2572]='h00002830;  wr_data_rom[ 2572]='h00000905;
    rd_cycle[ 2573] = 1'b0;  wr_cycle[ 2573] = 1'b1;  addr_rom[ 2573]='h00002834;  wr_data_rom[ 2573]='h00000e55;
    rd_cycle[ 2574] = 1'b0;  wr_cycle[ 2574] = 1'b1;  addr_rom[ 2574]='h00002838;  wr_data_rom[ 2574]='h00002b34;
    rd_cycle[ 2575] = 1'b0;  wr_cycle[ 2575] = 1'b1;  addr_rom[ 2575]='h0000283c;  wr_data_rom[ 2575]='h000000b6;
    rd_cycle[ 2576] = 1'b0;  wr_cycle[ 2576] = 1'b1;  addr_rom[ 2576]='h00002840;  wr_data_rom[ 2576]='h00001056;
    rd_cycle[ 2577] = 1'b0;  wr_cycle[ 2577] = 1'b1;  addr_rom[ 2577]='h00002844;  wr_data_rom[ 2577]='h0000051b;
    rd_cycle[ 2578] = 1'b0;  wr_cycle[ 2578] = 1'b1;  addr_rom[ 2578]='h00002848;  wr_data_rom[ 2578]='h00000e2f;
    rd_cycle[ 2579] = 1'b0;  wr_cycle[ 2579] = 1'b1;  addr_rom[ 2579]='h0000284c;  wr_data_rom[ 2579]='h000002bc;
    rd_cycle[ 2580] = 1'b0;  wr_cycle[ 2580] = 1'b1;  addr_rom[ 2580]='h00002850;  wr_data_rom[ 2580]='h00003546;
    rd_cycle[ 2581] = 1'b0;  wr_cycle[ 2581] = 1'b1;  addr_rom[ 2581]='h00002854;  wr_data_rom[ 2581]='h000003a3;
    rd_cycle[ 2582] = 1'b0;  wr_cycle[ 2582] = 1'b1;  addr_rom[ 2582]='h00002858;  wr_data_rom[ 2582]='h00001868;
    rd_cycle[ 2583] = 1'b0;  wr_cycle[ 2583] = 1'b1;  addr_rom[ 2583]='h0000285c;  wr_data_rom[ 2583]='h000030e3;
    rd_cycle[ 2584] = 1'b0;  wr_cycle[ 2584] = 1'b1;  addr_rom[ 2584]='h00002860;  wr_data_rom[ 2584]='h00002f00;
    rd_cycle[ 2585] = 1'b0;  wr_cycle[ 2585] = 1'b1;  addr_rom[ 2585]='h00002864;  wr_data_rom[ 2585]='h00002df9;
    rd_cycle[ 2586] = 1'b0;  wr_cycle[ 2586] = 1'b1;  addr_rom[ 2586]='h00002868;  wr_data_rom[ 2586]='h0000163c;
    rd_cycle[ 2587] = 1'b0;  wr_cycle[ 2587] = 1'b1;  addr_rom[ 2587]='h0000286c;  wr_data_rom[ 2587]='h000010d6;
    rd_cycle[ 2588] = 1'b0;  wr_cycle[ 2588] = 1'b1;  addr_rom[ 2588]='h00002870;  wr_data_rom[ 2588]='h00002f24;
    rd_cycle[ 2589] = 1'b0;  wr_cycle[ 2589] = 1'b1;  addr_rom[ 2589]='h00002874;  wr_data_rom[ 2589]='h000018c4;
    rd_cycle[ 2590] = 1'b0;  wr_cycle[ 2590] = 1'b1;  addr_rom[ 2590]='h00002878;  wr_data_rom[ 2590]='h00000ded;
    rd_cycle[ 2591] = 1'b0;  wr_cycle[ 2591] = 1'b1;  addr_rom[ 2591]='h0000287c;  wr_data_rom[ 2591]='h000027a3;
    rd_cycle[ 2592] = 1'b0;  wr_cycle[ 2592] = 1'b1;  addr_rom[ 2592]='h00002880;  wr_data_rom[ 2592]='h000008f2;
    rd_cycle[ 2593] = 1'b0;  wr_cycle[ 2593] = 1'b1;  addr_rom[ 2593]='h00002884;  wr_data_rom[ 2593]='h00003034;
    rd_cycle[ 2594] = 1'b0;  wr_cycle[ 2594] = 1'b1;  addr_rom[ 2594]='h00002888;  wr_data_rom[ 2594]='h00003613;
    rd_cycle[ 2595] = 1'b0;  wr_cycle[ 2595] = 1'b1;  addr_rom[ 2595]='h0000288c;  wr_data_rom[ 2595]='h00000d72;
    rd_cycle[ 2596] = 1'b0;  wr_cycle[ 2596] = 1'b1;  addr_rom[ 2596]='h00002890;  wr_data_rom[ 2596]='h000023d8;
    rd_cycle[ 2597] = 1'b0;  wr_cycle[ 2597] = 1'b1;  addr_rom[ 2597]='h00002894;  wr_data_rom[ 2597]='h00001bf2;
    rd_cycle[ 2598] = 1'b0;  wr_cycle[ 2598] = 1'b1;  addr_rom[ 2598]='h00002898;  wr_data_rom[ 2598]='h000023cf;
    rd_cycle[ 2599] = 1'b0;  wr_cycle[ 2599] = 1'b1;  addr_rom[ 2599]='h0000289c;  wr_data_rom[ 2599]='h00001a4a;
    rd_cycle[ 2600] = 1'b0;  wr_cycle[ 2600] = 1'b1;  addr_rom[ 2600]='h000028a0;  wr_data_rom[ 2600]='h0000284b;
    rd_cycle[ 2601] = 1'b0;  wr_cycle[ 2601] = 1'b1;  addr_rom[ 2601]='h000028a4;  wr_data_rom[ 2601]='h000013fd;
    rd_cycle[ 2602] = 1'b0;  wr_cycle[ 2602] = 1'b1;  addr_rom[ 2602]='h000028a8;  wr_data_rom[ 2602]='h00000e72;
    rd_cycle[ 2603] = 1'b0;  wr_cycle[ 2603] = 1'b1;  addr_rom[ 2603]='h000028ac;  wr_data_rom[ 2603]='h00003e31;
    rd_cycle[ 2604] = 1'b0;  wr_cycle[ 2604] = 1'b1;  addr_rom[ 2604]='h000028b0;  wr_data_rom[ 2604]='h0000138d;
    rd_cycle[ 2605] = 1'b0;  wr_cycle[ 2605] = 1'b1;  addr_rom[ 2605]='h000028b4;  wr_data_rom[ 2605]='h000026c4;
    rd_cycle[ 2606] = 1'b0;  wr_cycle[ 2606] = 1'b1;  addr_rom[ 2606]='h000028b8;  wr_data_rom[ 2606]='h00003b13;
    rd_cycle[ 2607] = 1'b0;  wr_cycle[ 2607] = 1'b1;  addr_rom[ 2607]='h000028bc;  wr_data_rom[ 2607]='h00003b3c;
    rd_cycle[ 2608] = 1'b0;  wr_cycle[ 2608] = 1'b1;  addr_rom[ 2608]='h000028c0;  wr_data_rom[ 2608]='h00002aae;
    rd_cycle[ 2609] = 1'b0;  wr_cycle[ 2609] = 1'b1;  addr_rom[ 2609]='h000028c4;  wr_data_rom[ 2609]='h00003793;
    rd_cycle[ 2610] = 1'b0;  wr_cycle[ 2610] = 1'b1;  addr_rom[ 2610]='h000028c8;  wr_data_rom[ 2610]='h00001d26;
    rd_cycle[ 2611] = 1'b0;  wr_cycle[ 2611] = 1'b1;  addr_rom[ 2611]='h000028cc;  wr_data_rom[ 2611]='h000007f4;
    rd_cycle[ 2612] = 1'b0;  wr_cycle[ 2612] = 1'b1;  addr_rom[ 2612]='h000028d0;  wr_data_rom[ 2612]='h00000fe2;
    rd_cycle[ 2613] = 1'b0;  wr_cycle[ 2613] = 1'b1;  addr_rom[ 2613]='h000028d4;  wr_data_rom[ 2613]='h00003d9b;
    rd_cycle[ 2614] = 1'b0;  wr_cycle[ 2614] = 1'b1;  addr_rom[ 2614]='h000028d8;  wr_data_rom[ 2614]='h000038b7;
    rd_cycle[ 2615] = 1'b0;  wr_cycle[ 2615] = 1'b1;  addr_rom[ 2615]='h000028dc;  wr_data_rom[ 2615]='h000039fb;
    rd_cycle[ 2616] = 1'b0;  wr_cycle[ 2616] = 1'b1;  addr_rom[ 2616]='h000028e0;  wr_data_rom[ 2616]='h00002d1d;
    rd_cycle[ 2617] = 1'b0;  wr_cycle[ 2617] = 1'b1;  addr_rom[ 2617]='h000028e4;  wr_data_rom[ 2617]='h000026dc;
    rd_cycle[ 2618] = 1'b0;  wr_cycle[ 2618] = 1'b1;  addr_rom[ 2618]='h000028e8;  wr_data_rom[ 2618]='h00003a31;
    rd_cycle[ 2619] = 1'b0;  wr_cycle[ 2619] = 1'b1;  addr_rom[ 2619]='h000028ec;  wr_data_rom[ 2619]='h00003eb3;
    rd_cycle[ 2620] = 1'b0;  wr_cycle[ 2620] = 1'b1;  addr_rom[ 2620]='h000028f0;  wr_data_rom[ 2620]='h00002eaf;
    rd_cycle[ 2621] = 1'b0;  wr_cycle[ 2621] = 1'b1;  addr_rom[ 2621]='h000028f4;  wr_data_rom[ 2621]='h00000c94;
    rd_cycle[ 2622] = 1'b0;  wr_cycle[ 2622] = 1'b1;  addr_rom[ 2622]='h000028f8;  wr_data_rom[ 2622]='h00003e86;
    rd_cycle[ 2623] = 1'b0;  wr_cycle[ 2623] = 1'b1;  addr_rom[ 2623]='h000028fc;  wr_data_rom[ 2623]='h000039e9;
    rd_cycle[ 2624] = 1'b0;  wr_cycle[ 2624] = 1'b1;  addr_rom[ 2624]='h00002900;  wr_data_rom[ 2624]='h000029ec;
    rd_cycle[ 2625] = 1'b0;  wr_cycle[ 2625] = 1'b1;  addr_rom[ 2625]='h00002904;  wr_data_rom[ 2625]='h0000317a;
    rd_cycle[ 2626] = 1'b0;  wr_cycle[ 2626] = 1'b1;  addr_rom[ 2626]='h00002908;  wr_data_rom[ 2626]='h00002da6;
    rd_cycle[ 2627] = 1'b0;  wr_cycle[ 2627] = 1'b1;  addr_rom[ 2627]='h0000290c;  wr_data_rom[ 2627]='h00001872;
    rd_cycle[ 2628] = 1'b0;  wr_cycle[ 2628] = 1'b1;  addr_rom[ 2628]='h00002910;  wr_data_rom[ 2628]='h000026a8;
    rd_cycle[ 2629] = 1'b0;  wr_cycle[ 2629] = 1'b1;  addr_rom[ 2629]='h00002914;  wr_data_rom[ 2629]='h00002f91;
    rd_cycle[ 2630] = 1'b0;  wr_cycle[ 2630] = 1'b1;  addr_rom[ 2630]='h00002918;  wr_data_rom[ 2630]='h00003a25;
    rd_cycle[ 2631] = 1'b0;  wr_cycle[ 2631] = 1'b1;  addr_rom[ 2631]='h0000291c;  wr_data_rom[ 2631]='h00001cbf;
    rd_cycle[ 2632] = 1'b0;  wr_cycle[ 2632] = 1'b1;  addr_rom[ 2632]='h00002920;  wr_data_rom[ 2632]='h00000350;
    rd_cycle[ 2633] = 1'b0;  wr_cycle[ 2633] = 1'b1;  addr_rom[ 2633]='h00002924;  wr_data_rom[ 2633]='h000029cf;
    rd_cycle[ 2634] = 1'b0;  wr_cycle[ 2634] = 1'b1;  addr_rom[ 2634]='h00002928;  wr_data_rom[ 2634]='h00000f9d;
    rd_cycle[ 2635] = 1'b0;  wr_cycle[ 2635] = 1'b1;  addr_rom[ 2635]='h0000292c;  wr_data_rom[ 2635]='h0000266c;
    rd_cycle[ 2636] = 1'b0;  wr_cycle[ 2636] = 1'b1;  addr_rom[ 2636]='h00002930;  wr_data_rom[ 2636]='h00002715;
    rd_cycle[ 2637] = 1'b0;  wr_cycle[ 2637] = 1'b1;  addr_rom[ 2637]='h00002934;  wr_data_rom[ 2637]='h000015a7;
    rd_cycle[ 2638] = 1'b0;  wr_cycle[ 2638] = 1'b1;  addr_rom[ 2638]='h00002938;  wr_data_rom[ 2638]='h00003047;
    rd_cycle[ 2639] = 1'b0;  wr_cycle[ 2639] = 1'b1;  addr_rom[ 2639]='h0000293c;  wr_data_rom[ 2639]='h00002aa6;
    rd_cycle[ 2640] = 1'b0;  wr_cycle[ 2640] = 1'b1;  addr_rom[ 2640]='h00002940;  wr_data_rom[ 2640]='h000015bd;
    rd_cycle[ 2641] = 1'b0;  wr_cycle[ 2641] = 1'b1;  addr_rom[ 2641]='h00002944;  wr_data_rom[ 2641]='h0000011a;
    rd_cycle[ 2642] = 1'b0;  wr_cycle[ 2642] = 1'b1;  addr_rom[ 2642]='h00002948;  wr_data_rom[ 2642]='h000032c0;
    rd_cycle[ 2643] = 1'b0;  wr_cycle[ 2643] = 1'b1;  addr_rom[ 2643]='h0000294c;  wr_data_rom[ 2643]='h00002f70;
    rd_cycle[ 2644] = 1'b0;  wr_cycle[ 2644] = 1'b1;  addr_rom[ 2644]='h00002950;  wr_data_rom[ 2644]='h00000425;
    rd_cycle[ 2645] = 1'b0;  wr_cycle[ 2645] = 1'b1;  addr_rom[ 2645]='h00002954;  wr_data_rom[ 2645]='h00000524;
    rd_cycle[ 2646] = 1'b0;  wr_cycle[ 2646] = 1'b1;  addr_rom[ 2646]='h00002958;  wr_data_rom[ 2646]='h00001159;
    rd_cycle[ 2647] = 1'b0;  wr_cycle[ 2647] = 1'b1;  addr_rom[ 2647]='h0000295c;  wr_data_rom[ 2647]='h000007f2;
    rd_cycle[ 2648] = 1'b0;  wr_cycle[ 2648] = 1'b1;  addr_rom[ 2648]='h00002960;  wr_data_rom[ 2648]='h00003480;
    rd_cycle[ 2649] = 1'b0;  wr_cycle[ 2649] = 1'b1;  addr_rom[ 2649]='h00002964;  wr_data_rom[ 2649]='h00000454;
    rd_cycle[ 2650] = 1'b0;  wr_cycle[ 2650] = 1'b1;  addr_rom[ 2650]='h00002968;  wr_data_rom[ 2650]='h00002d5a;
    rd_cycle[ 2651] = 1'b0;  wr_cycle[ 2651] = 1'b1;  addr_rom[ 2651]='h0000296c;  wr_data_rom[ 2651]='h00001b3d;
    rd_cycle[ 2652] = 1'b0;  wr_cycle[ 2652] = 1'b1;  addr_rom[ 2652]='h00002970;  wr_data_rom[ 2652]='h00003b79;
    rd_cycle[ 2653] = 1'b0;  wr_cycle[ 2653] = 1'b1;  addr_rom[ 2653]='h00002974;  wr_data_rom[ 2653]='h000033de;
    rd_cycle[ 2654] = 1'b0;  wr_cycle[ 2654] = 1'b1;  addr_rom[ 2654]='h00002978;  wr_data_rom[ 2654]='h00000d27;
    rd_cycle[ 2655] = 1'b0;  wr_cycle[ 2655] = 1'b1;  addr_rom[ 2655]='h0000297c;  wr_data_rom[ 2655]='h00001cff;
    rd_cycle[ 2656] = 1'b0;  wr_cycle[ 2656] = 1'b1;  addr_rom[ 2656]='h00002980;  wr_data_rom[ 2656]='h00002769;
    rd_cycle[ 2657] = 1'b0;  wr_cycle[ 2657] = 1'b1;  addr_rom[ 2657]='h00002984;  wr_data_rom[ 2657]='h000018e7;
    rd_cycle[ 2658] = 1'b0;  wr_cycle[ 2658] = 1'b1;  addr_rom[ 2658]='h00002988;  wr_data_rom[ 2658]='h00003c9d;
    rd_cycle[ 2659] = 1'b0;  wr_cycle[ 2659] = 1'b1;  addr_rom[ 2659]='h0000298c;  wr_data_rom[ 2659]='h00002860;
    rd_cycle[ 2660] = 1'b0;  wr_cycle[ 2660] = 1'b1;  addr_rom[ 2660]='h00002990;  wr_data_rom[ 2660]='h00000bba;
    rd_cycle[ 2661] = 1'b0;  wr_cycle[ 2661] = 1'b1;  addr_rom[ 2661]='h00002994;  wr_data_rom[ 2661]='h0000317c;
    rd_cycle[ 2662] = 1'b0;  wr_cycle[ 2662] = 1'b1;  addr_rom[ 2662]='h00002998;  wr_data_rom[ 2662]='h00002771;
    rd_cycle[ 2663] = 1'b0;  wr_cycle[ 2663] = 1'b1;  addr_rom[ 2663]='h0000299c;  wr_data_rom[ 2663]='h0000173e;
    rd_cycle[ 2664] = 1'b0;  wr_cycle[ 2664] = 1'b1;  addr_rom[ 2664]='h000029a0;  wr_data_rom[ 2664]='h00003973;
    rd_cycle[ 2665] = 1'b0;  wr_cycle[ 2665] = 1'b1;  addr_rom[ 2665]='h000029a4;  wr_data_rom[ 2665]='h000026ff;
    rd_cycle[ 2666] = 1'b0;  wr_cycle[ 2666] = 1'b1;  addr_rom[ 2666]='h000029a8;  wr_data_rom[ 2666]='h000006fa;
    rd_cycle[ 2667] = 1'b0;  wr_cycle[ 2667] = 1'b1;  addr_rom[ 2667]='h000029ac;  wr_data_rom[ 2667]='h00001bae;
    rd_cycle[ 2668] = 1'b0;  wr_cycle[ 2668] = 1'b1;  addr_rom[ 2668]='h000029b0;  wr_data_rom[ 2668]='h00003ac2;
    rd_cycle[ 2669] = 1'b0;  wr_cycle[ 2669] = 1'b1;  addr_rom[ 2669]='h000029b4;  wr_data_rom[ 2669]='h000039b8;
    rd_cycle[ 2670] = 1'b0;  wr_cycle[ 2670] = 1'b1;  addr_rom[ 2670]='h000029b8;  wr_data_rom[ 2670]='h00003ae9;
    rd_cycle[ 2671] = 1'b0;  wr_cycle[ 2671] = 1'b1;  addr_rom[ 2671]='h000029bc;  wr_data_rom[ 2671]='h0000306b;
    rd_cycle[ 2672] = 1'b0;  wr_cycle[ 2672] = 1'b1;  addr_rom[ 2672]='h000029c0;  wr_data_rom[ 2672]='h00003984;
    rd_cycle[ 2673] = 1'b0;  wr_cycle[ 2673] = 1'b1;  addr_rom[ 2673]='h000029c4;  wr_data_rom[ 2673]='h00003b68;
    rd_cycle[ 2674] = 1'b0;  wr_cycle[ 2674] = 1'b1;  addr_rom[ 2674]='h000029c8;  wr_data_rom[ 2674]='h00003389;
    rd_cycle[ 2675] = 1'b0;  wr_cycle[ 2675] = 1'b1;  addr_rom[ 2675]='h000029cc;  wr_data_rom[ 2675]='h0000071f;
    rd_cycle[ 2676] = 1'b0;  wr_cycle[ 2676] = 1'b1;  addr_rom[ 2676]='h000029d0;  wr_data_rom[ 2676]='h00000566;
    rd_cycle[ 2677] = 1'b0;  wr_cycle[ 2677] = 1'b1;  addr_rom[ 2677]='h000029d4;  wr_data_rom[ 2677]='h00001fff;
    rd_cycle[ 2678] = 1'b0;  wr_cycle[ 2678] = 1'b1;  addr_rom[ 2678]='h000029d8;  wr_data_rom[ 2678]='h000030fc;
    rd_cycle[ 2679] = 1'b0;  wr_cycle[ 2679] = 1'b1;  addr_rom[ 2679]='h000029dc;  wr_data_rom[ 2679]='h00000f8a;
    rd_cycle[ 2680] = 1'b0;  wr_cycle[ 2680] = 1'b1;  addr_rom[ 2680]='h000029e0;  wr_data_rom[ 2680]='h00001268;
    rd_cycle[ 2681] = 1'b0;  wr_cycle[ 2681] = 1'b1;  addr_rom[ 2681]='h000029e4;  wr_data_rom[ 2681]='h00003c6c;
    rd_cycle[ 2682] = 1'b0;  wr_cycle[ 2682] = 1'b1;  addr_rom[ 2682]='h000029e8;  wr_data_rom[ 2682]='h00003da8;
    rd_cycle[ 2683] = 1'b0;  wr_cycle[ 2683] = 1'b1;  addr_rom[ 2683]='h000029ec;  wr_data_rom[ 2683]='h00003fe2;
    rd_cycle[ 2684] = 1'b0;  wr_cycle[ 2684] = 1'b1;  addr_rom[ 2684]='h000029f0;  wr_data_rom[ 2684]='h00002a3a;
    rd_cycle[ 2685] = 1'b0;  wr_cycle[ 2685] = 1'b1;  addr_rom[ 2685]='h000029f4;  wr_data_rom[ 2685]='h000039bd;
    rd_cycle[ 2686] = 1'b0;  wr_cycle[ 2686] = 1'b1;  addr_rom[ 2686]='h000029f8;  wr_data_rom[ 2686]='h00000fe1;
    rd_cycle[ 2687] = 1'b0;  wr_cycle[ 2687] = 1'b1;  addr_rom[ 2687]='h000029fc;  wr_data_rom[ 2687]='h00001745;
    rd_cycle[ 2688] = 1'b0;  wr_cycle[ 2688] = 1'b1;  addr_rom[ 2688]='h00002a00;  wr_data_rom[ 2688]='h000014c7;
    rd_cycle[ 2689] = 1'b0;  wr_cycle[ 2689] = 1'b1;  addr_rom[ 2689]='h00002a04;  wr_data_rom[ 2689]='h000013a1;
    rd_cycle[ 2690] = 1'b0;  wr_cycle[ 2690] = 1'b1;  addr_rom[ 2690]='h00002a08;  wr_data_rom[ 2690]='h000038dd;
    rd_cycle[ 2691] = 1'b0;  wr_cycle[ 2691] = 1'b1;  addr_rom[ 2691]='h00002a0c;  wr_data_rom[ 2691]='h0000195a;
    rd_cycle[ 2692] = 1'b0;  wr_cycle[ 2692] = 1'b1;  addr_rom[ 2692]='h00002a10;  wr_data_rom[ 2692]='h000015dc;
    rd_cycle[ 2693] = 1'b0;  wr_cycle[ 2693] = 1'b1;  addr_rom[ 2693]='h00002a14;  wr_data_rom[ 2693]='h00002e59;
    rd_cycle[ 2694] = 1'b0;  wr_cycle[ 2694] = 1'b1;  addr_rom[ 2694]='h00002a18;  wr_data_rom[ 2694]='h00002aab;
    rd_cycle[ 2695] = 1'b0;  wr_cycle[ 2695] = 1'b1;  addr_rom[ 2695]='h00002a1c;  wr_data_rom[ 2695]='h000009b6;
    rd_cycle[ 2696] = 1'b0;  wr_cycle[ 2696] = 1'b1;  addr_rom[ 2696]='h00002a20;  wr_data_rom[ 2696]='h000020d8;
    rd_cycle[ 2697] = 1'b0;  wr_cycle[ 2697] = 1'b1;  addr_rom[ 2697]='h00002a24;  wr_data_rom[ 2697]='h000006da;
    rd_cycle[ 2698] = 1'b0;  wr_cycle[ 2698] = 1'b1;  addr_rom[ 2698]='h00002a28;  wr_data_rom[ 2698]='h0000164e;
    rd_cycle[ 2699] = 1'b0;  wr_cycle[ 2699] = 1'b1;  addr_rom[ 2699]='h00002a2c;  wr_data_rom[ 2699]='h000009d9;
    rd_cycle[ 2700] = 1'b0;  wr_cycle[ 2700] = 1'b1;  addr_rom[ 2700]='h00002a30;  wr_data_rom[ 2700]='h000012c6;
    rd_cycle[ 2701] = 1'b0;  wr_cycle[ 2701] = 1'b1;  addr_rom[ 2701]='h00002a34;  wr_data_rom[ 2701]='h00000fb3;
    rd_cycle[ 2702] = 1'b0;  wr_cycle[ 2702] = 1'b1;  addr_rom[ 2702]='h00002a38;  wr_data_rom[ 2702]='h00001082;
    rd_cycle[ 2703] = 1'b0;  wr_cycle[ 2703] = 1'b1;  addr_rom[ 2703]='h00002a3c;  wr_data_rom[ 2703]='h000018e2;
    rd_cycle[ 2704] = 1'b0;  wr_cycle[ 2704] = 1'b1;  addr_rom[ 2704]='h00002a40;  wr_data_rom[ 2704]='h000001e9;
    rd_cycle[ 2705] = 1'b0;  wr_cycle[ 2705] = 1'b1;  addr_rom[ 2705]='h00002a44;  wr_data_rom[ 2705]='h00003b5a;
    rd_cycle[ 2706] = 1'b0;  wr_cycle[ 2706] = 1'b1;  addr_rom[ 2706]='h00002a48;  wr_data_rom[ 2706]='h00002493;
    rd_cycle[ 2707] = 1'b0;  wr_cycle[ 2707] = 1'b1;  addr_rom[ 2707]='h00002a4c;  wr_data_rom[ 2707]='h000025fa;
    rd_cycle[ 2708] = 1'b0;  wr_cycle[ 2708] = 1'b1;  addr_rom[ 2708]='h00002a50;  wr_data_rom[ 2708]='h00001e62;
    rd_cycle[ 2709] = 1'b0;  wr_cycle[ 2709] = 1'b1;  addr_rom[ 2709]='h00002a54;  wr_data_rom[ 2709]='h0000034f;
    rd_cycle[ 2710] = 1'b0;  wr_cycle[ 2710] = 1'b1;  addr_rom[ 2710]='h00002a58;  wr_data_rom[ 2710]='h0000319c;
    rd_cycle[ 2711] = 1'b0;  wr_cycle[ 2711] = 1'b1;  addr_rom[ 2711]='h00002a5c;  wr_data_rom[ 2711]='h000010e9;
    rd_cycle[ 2712] = 1'b0;  wr_cycle[ 2712] = 1'b1;  addr_rom[ 2712]='h00002a60;  wr_data_rom[ 2712]='h000030cb;
    rd_cycle[ 2713] = 1'b0;  wr_cycle[ 2713] = 1'b1;  addr_rom[ 2713]='h00002a64;  wr_data_rom[ 2713]='h0000005b;
    rd_cycle[ 2714] = 1'b0;  wr_cycle[ 2714] = 1'b1;  addr_rom[ 2714]='h00002a68;  wr_data_rom[ 2714]='h000001ae;
    rd_cycle[ 2715] = 1'b0;  wr_cycle[ 2715] = 1'b1;  addr_rom[ 2715]='h00002a6c;  wr_data_rom[ 2715]='h00000c04;
    rd_cycle[ 2716] = 1'b0;  wr_cycle[ 2716] = 1'b1;  addr_rom[ 2716]='h00002a70;  wr_data_rom[ 2716]='h000026d5;
    rd_cycle[ 2717] = 1'b0;  wr_cycle[ 2717] = 1'b1;  addr_rom[ 2717]='h00002a74;  wr_data_rom[ 2717]='h000013e9;
    rd_cycle[ 2718] = 1'b0;  wr_cycle[ 2718] = 1'b1;  addr_rom[ 2718]='h00002a78;  wr_data_rom[ 2718]='h00001b1c;
    rd_cycle[ 2719] = 1'b0;  wr_cycle[ 2719] = 1'b1;  addr_rom[ 2719]='h00002a7c;  wr_data_rom[ 2719]='h0000383b;
    rd_cycle[ 2720] = 1'b0;  wr_cycle[ 2720] = 1'b1;  addr_rom[ 2720]='h00002a80;  wr_data_rom[ 2720]='h00002a0c;
    rd_cycle[ 2721] = 1'b0;  wr_cycle[ 2721] = 1'b1;  addr_rom[ 2721]='h00002a84;  wr_data_rom[ 2721]='h0000126b;
    rd_cycle[ 2722] = 1'b0;  wr_cycle[ 2722] = 1'b1;  addr_rom[ 2722]='h00002a88;  wr_data_rom[ 2722]='h00000a9e;
    rd_cycle[ 2723] = 1'b0;  wr_cycle[ 2723] = 1'b1;  addr_rom[ 2723]='h00002a8c;  wr_data_rom[ 2723]='h000020c1;
    rd_cycle[ 2724] = 1'b0;  wr_cycle[ 2724] = 1'b1;  addr_rom[ 2724]='h00002a90;  wr_data_rom[ 2724]='h00003a43;
    rd_cycle[ 2725] = 1'b0;  wr_cycle[ 2725] = 1'b1;  addr_rom[ 2725]='h00002a94;  wr_data_rom[ 2725]='h000005c4;
    rd_cycle[ 2726] = 1'b0;  wr_cycle[ 2726] = 1'b1;  addr_rom[ 2726]='h00002a98;  wr_data_rom[ 2726]='h00001073;
    rd_cycle[ 2727] = 1'b0;  wr_cycle[ 2727] = 1'b1;  addr_rom[ 2727]='h00002a9c;  wr_data_rom[ 2727]='h000025c5;
    rd_cycle[ 2728] = 1'b0;  wr_cycle[ 2728] = 1'b1;  addr_rom[ 2728]='h00002aa0;  wr_data_rom[ 2728]='h00002116;
    rd_cycle[ 2729] = 1'b0;  wr_cycle[ 2729] = 1'b1;  addr_rom[ 2729]='h00002aa4;  wr_data_rom[ 2729]='h00002df8;
    rd_cycle[ 2730] = 1'b0;  wr_cycle[ 2730] = 1'b1;  addr_rom[ 2730]='h00002aa8;  wr_data_rom[ 2730]='h000038b3;
    rd_cycle[ 2731] = 1'b0;  wr_cycle[ 2731] = 1'b1;  addr_rom[ 2731]='h00002aac;  wr_data_rom[ 2731]='h00002636;
    rd_cycle[ 2732] = 1'b0;  wr_cycle[ 2732] = 1'b1;  addr_rom[ 2732]='h00002ab0;  wr_data_rom[ 2732]='h00000cc3;
    rd_cycle[ 2733] = 1'b0;  wr_cycle[ 2733] = 1'b1;  addr_rom[ 2733]='h00002ab4;  wr_data_rom[ 2733]='h000032e8;
    rd_cycle[ 2734] = 1'b0;  wr_cycle[ 2734] = 1'b1;  addr_rom[ 2734]='h00002ab8;  wr_data_rom[ 2734]='h000000f6;
    rd_cycle[ 2735] = 1'b0;  wr_cycle[ 2735] = 1'b1;  addr_rom[ 2735]='h00002abc;  wr_data_rom[ 2735]='h00001266;
    rd_cycle[ 2736] = 1'b0;  wr_cycle[ 2736] = 1'b1;  addr_rom[ 2736]='h00002ac0;  wr_data_rom[ 2736]='h000024ad;
    rd_cycle[ 2737] = 1'b0;  wr_cycle[ 2737] = 1'b1;  addr_rom[ 2737]='h00002ac4;  wr_data_rom[ 2737]='h000036fb;
    rd_cycle[ 2738] = 1'b0;  wr_cycle[ 2738] = 1'b1;  addr_rom[ 2738]='h00002ac8;  wr_data_rom[ 2738]='h000011f5;
    rd_cycle[ 2739] = 1'b0;  wr_cycle[ 2739] = 1'b1;  addr_rom[ 2739]='h00002acc;  wr_data_rom[ 2739]='h0000022e;
    rd_cycle[ 2740] = 1'b0;  wr_cycle[ 2740] = 1'b1;  addr_rom[ 2740]='h00002ad0;  wr_data_rom[ 2740]='h0000101b;
    rd_cycle[ 2741] = 1'b0;  wr_cycle[ 2741] = 1'b1;  addr_rom[ 2741]='h00002ad4;  wr_data_rom[ 2741]='h00001099;
    rd_cycle[ 2742] = 1'b0;  wr_cycle[ 2742] = 1'b1;  addr_rom[ 2742]='h00002ad8;  wr_data_rom[ 2742]='h00003ba8;
    rd_cycle[ 2743] = 1'b0;  wr_cycle[ 2743] = 1'b1;  addr_rom[ 2743]='h00002adc;  wr_data_rom[ 2743]='h0000350d;
    rd_cycle[ 2744] = 1'b0;  wr_cycle[ 2744] = 1'b1;  addr_rom[ 2744]='h00002ae0;  wr_data_rom[ 2744]='h0000195a;
    rd_cycle[ 2745] = 1'b0;  wr_cycle[ 2745] = 1'b1;  addr_rom[ 2745]='h00002ae4;  wr_data_rom[ 2745]='h000019b5;
    rd_cycle[ 2746] = 1'b0;  wr_cycle[ 2746] = 1'b1;  addr_rom[ 2746]='h00002ae8;  wr_data_rom[ 2746]='h00000c2b;
    rd_cycle[ 2747] = 1'b0;  wr_cycle[ 2747] = 1'b1;  addr_rom[ 2747]='h00002aec;  wr_data_rom[ 2747]='h00000e02;
    rd_cycle[ 2748] = 1'b0;  wr_cycle[ 2748] = 1'b1;  addr_rom[ 2748]='h00002af0;  wr_data_rom[ 2748]='h00000dd9;
    rd_cycle[ 2749] = 1'b0;  wr_cycle[ 2749] = 1'b1;  addr_rom[ 2749]='h00002af4;  wr_data_rom[ 2749]='h00000551;
    rd_cycle[ 2750] = 1'b0;  wr_cycle[ 2750] = 1'b1;  addr_rom[ 2750]='h00002af8;  wr_data_rom[ 2750]='h00002374;
    rd_cycle[ 2751] = 1'b0;  wr_cycle[ 2751] = 1'b1;  addr_rom[ 2751]='h00002afc;  wr_data_rom[ 2751]='h00002447;
    rd_cycle[ 2752] = 1'b0;  wr_cycle[ 2752] = 1'b1;  addr_rom[ 2752]='h00002b00;  wr_data_rom[ 2752]='h0000264f;
    rd_cycle[ 2753] = 1'b0;  wr_cycle[ 2753] = 1'b1;  addr_rom[ 2753]='h00002b04;  wr_data_rom[ 2753]='h00001e43;
    rd_cycle[ 2754] = 1'b0;  wr_cycle[ 2754] = 1'b1;  addr_rom[ 2754]='h00002b08;  wr_data_rom[ 2754]='h00000e5a;
    rd_cycle[ 2755] = 1'b0;  wr_cycle[ 2755] = 1'b1;  addr_rom[ 2755]='h00002b0c;  wr_data_rom[ 2755]='h00001950;
    rd_cycle[ 2756] = 1'b0;  wr_cycle[ 2756] = 1'b1;  addr_rom[ 2756]='h00002b10;  wr_data_rom[ 2756]='h00001ce3;
    rd_cycle[ 2757] = 1'b0;  wr_cycle[ 2757] = 1'b1;  addr_rom[ 2757]='h00002b14;  wr_data_rom[ 2757]='h000027c2;
    rd_cycle[ 2758] = 1'b0;  wr_cycle[ 2758] = 1'b1;  addr_rom[ 2758]='h00002b18;  wr_data_rom[ 2758]='h00001d7d;
    rd_cycle[ 2759] = 1'b0;  wr_cycle[ 2759] = 1'b1;  addr_rom[ 2759]='h00002b1c;  wr_data_rom[ 2759]='h000011b0;
    rd_cycle[ 2760] = 1'b0;  wr_cycle[ 2760] = 1'b1;  addr_rom[ 2760]='h00002b20;  wr_data_rom[ 2760]='h0000247f;
    rd_cycle[ 2761] = 1'b0;  wr_cycle[ 2761] = 1'b1;  addr_rom[ 2761]='h00002b24;  wr_data_rom[ 2761]='h00001bdf;
    rd_cycle[ 2762] = 1'b0;  wr_cycle[ 2762] = 1'b1;  addr_rom[ 2762]='h00002b28;  wr_data_rom[ 2762]='h00002e0c;
    rd_cycle[ 2763] = 1'b0;  wr_cycle[ 2763] = 1'b1;  addr_rom[ 2763]='h00002b2c;  wr_data_rom[ 2763]='h00000856;
    rd_cycle[ 2764] = 1'b0;  wr_cycle[ 2764] = 1'b1;  addr_rom[ 2764]='h00002b30;  wr_data_rom[ 2764]='h00003f37;
    rd_cycle[ 2765] = 1'b0;  wr_cycle[ 2765] = 1'b1;  addr_rom[ 2765]='h00002b34;  wr_data_rom[ 2765]='h00003b27;
    rd_cycle[ 2766] = 1'b0;  wr_cycle[ 2766] = 1'b1;  addr_rom[ 2766]='h00002b38;  wr_data_rom[ 2766]='h0000055d;
    rd_cycle[ 2767] = 1'b0;  wr_cycle[ 2767] = 1'b1;  addr_rom[ 2767]='h00002b3c;  wr_data_rom[ 2767]='h000011f0;
    rd_cycle[ 2768] = 1'b0;  wr_cycle[ 2768] = 1'b1;  addr_rom[ 2768]='h00002b40;  wr_data_rom[ 2768]='h00003249;
    rd_cycle[ 2769] = 1'b0;  wr_cycle[ 2769] = 1'b1;  addr_rom[ 2769]='h00002b44;  wr_data_rom[ 2769]='h00000d72;
    rd_cycle[ 2770] = 1'b0;  wr_cycle[ 2770] = 1'b1;  addr_rom[ 2770]='h00002b48;  wr_data_rom[ 2770]='h00002d9d;
    rd_cycle[ 2771] = 1'b0;  wr_cycle[ 2771] = 1'b1;  addr_rom[ 2771]='h00002b4c;  wr_data_rom[ 2771]='h00003e6a;
    rd_cycle[ 2772] = 1'b0;  wr_cycle[ 2772] = 1'b1;  addr_rom[ 2772]='h00002b50;  wr_data_rom[ 2772]='h00002a8b;
    rd_cycle[ 2773] = 1'b0;  wr_cycle[ 2773] = 1'b1;  addr_rom[ 2773]='h00002b54;  wr_data_rom[ 2773]='h00002196;
    rd_cycle[ 2774] = 1'b0;  wr_cycle[ 2774] = 1'b1;  addr_rom[ 2774]='h00002b58;  wr_data_rom[ 2774]='h00002b98;
    rd_cycle[ 2775] = 1'b0;  wr_cycle[ 2775] = 1'b1;  addr_rom[ 2775]='h00002b5c;  wr_data_rom[ 2775]='h000031c3;
    rd_cycle[ 2776] = 1'b0;  wr_cycle[ 2776] = 1'b1;  addr_rom[ 2776]='h00002b60;  wr_data_rom[ 2776]='h000005c1;
    rd_cycle[ 2777] = 1'b0;  wr_cycle[ 2777] = 1'b1;  addr_rom[ 2777]='h00002b64;  wr_data_rom[ 2777]='h000007d4;
    rd_cycle[ 2778] = 1'b0;  wr_cycle[ 2778] = 1'b1;  addr_rom[ 2778]='h00002b68;  wr_data_rom[ 2778]='h000035f4;
    rd_cycle[ 2779] = 1'b0;  wr_cycle[ 2779] = 1'b1;  addr_rom[ 2779]='h00002b6c;  wr_data_rom[ 2779]='h000004a2;
    rd_cycle[ 2780] = 1'b0;  wr_cycle[ 2780] = 1'b1;  addr_rom[ 2780]='h00002b70;  wr_data_rom[ 2780]='h0000276c;
    rd_cycle[ 2781] = 1'b0;  wr_cycle[ 2781] = 1'b1;  addr_rom[ 2781]='h00002b74;  wr_data_rom[ 2781]='h000023b6;
    rd_cycle[ 2782] = 1'b0;  wr_cycle[ 2782] = 1'b1;  addr_rom[ 2782]='h00002b78;  wr_data_rom[ 2782]='h00001375;
    rd_cycle[ 2783] = 1'b0;  wr_cycle[ 2783] = 1'b1;  addr_rom[ 2783]='h00002b7c;  wr_data_rom[ 2783]='h000038e7;
    rd_cycle[ 2784] = 1'b0;  wr_cycle[ 2784] = 1'b1;  addr_rom[ 2784]='h00002b80;  wr_data_rom[ 2784]='h00001bfe;
    rd_cycle[ 2785] = 1'b0;  wr_cycle[ 2785] = 1'b1;  addr_rom[ 2785]='h00002b84;  wr_data_rom[ 2785]='h000027bb;
    rd_cycle[ 2786] = 1'b0;  wr_cycle[ 2786] = 1'b1;  addr_rom[ 2786]='h00002b88;  wr_data_rom[ 2786]='h000015d9;
    rd_cycle[ 2787] = 1'b0;  wr_cycle[ 2787] = 1'b1;  addr_rom[ 2787]='h00002b8c;  wr_data_rom[ 2787]='h00001dbc;
    rd_cycle[ 2788] = 1'b0;  wr_cycle[ 2788] = 1'b1;  addr_rom[ 2788]='h00002b90;  wr_data_rom[ 2788]='h00002d0c;
    rd_cycle[ 2789] = 1'b0;  wr_cycle[ 2789] = 1'b1;  addr_rom[ 2789]='h00002b94;  wr_data_rom[ 2789]='h00002817;
    rd_cycle[ 2790] = 1'b0;  wr_cycle[ 2790] = 1'b1;  addr_rom[ 2790]='h00002b98;  wr_data_rom[ 2790]='h00000d8a;
    rd_cycle[ 2791] = 1'b0;  wr_cycle[ 2791] = 1'b1;  addr_rom[ 2791]='h00002b9c;  wr_data_rom[ 2791]='h00001e84;
    rd_cycle[ 2792] = 1'b0;  wr_cycle[ 2792] = 1'b1;  addr_rom[ 2792]='h00002ba0;  wr_data_rom[ 2792]='h0000054f;
    rd_cycle[ 2793] = 1'b0;  wr_cycle[ 2793] = 1'b1;  addr_rom[ 2793]='h00002ba4;  wr_data_rom[ 2793]='h000016ad;
    rd_cycle[ 2794] = 1'b0;  wr_cycle[ 2794] = 1'b1;  addr_rom[ 2794]='h00002ba8;  wr_data_rom[ 2794]='h0000219c;
    rd_cycle[ 2795] = 1'b0;  wr_cycle[ 2795] = 1'b1;  addr_rom[ 2795]='h00002bac;  wr_data_rom[ 2795]='h00000c41;
    rd_cycle[ 2796] = 1'b0;  wr_cycle[ 2796] = 1'b1;  addr_rom[ 2796]='h00002bb0;  wr_data_rom[ 2796]='h00001985;
    rd_cycle[ 2797] = 1'b0;  wr_cycle[ 2797] = 1'b1;  addr_rom[ 2797]='h00002bb4;  wr_data_rom[ 2797]='h000018c9;
    rd_cycle[ 2798] = 1'b0;  wr_cycle[ 2798] = 1'b1;  addr_rom[ 2798]='h00002bb8;  wr_data_rom[ 2798]='h0000365c;
    rd_cycle[ 2799] = 1'b0;  wr_cycle[ 2799] = 1'b1;  addr_rom[ 2799]='h00002bbc;  wr_data_rom[ 2799]='h00000c8e;
    rd_cycle[ 2800] = 1'b0;  wr_cycle[ 2800] = 1'b1;  addr_rom[ 2800]='h00002bc0;  wr_data_rom[ 2800]='h00000c66;
    rd_cycle[ 2801] = 1'b0;  wr_cycle[ 2801] = 1'b1;  addr_rom[ 2801]='h00002bc4;  wr_data_rom[ 2801]='h00002095;
    rd_cycle[ 2802] = 1'b0;  wr_cycle[ 2802] = 1'b1;  addr_rom[ 2802]='h00002bc8;  wr_data_rom[ 2802]='h000004ff;
    rd_cycle[ 2803] = 1'b0;  wr_cycle[ 2803] = 1'b1;  addr_rom[ 2803]='h00002bcc;  wr_data_rom[ 2803]='h00001668;
    rd_cycle[ 2804] = 1'b0;  wr_cycle[ 2804] = 1'b1;  addr_rom[ 2804]='h00002bd0;  wr_data_rom[ 2804]='h0000322e;
    rd_cycle[ 2805] = 1'b0;  wr_cycle[ 2805] = 1'b1;  addr_rom[ 2805]='h00002bd4;  wr_data_rom[ 2805]='h000000ac;
    rd_cycle[ 2806] = 1'b0;  wr_cycle[ 2806] = 1'b1;  addr_rom[ 2806]='h00002bd8;  wr_data_rom[ 2806]='h00000b66;
    rd_cycle[ 2807] = 1'b0;  wr_cycle[ 2807] = 1'b1;  addr_rom[ 2807]='h00002bdc;  wr_data_rom[ 2807]='h00002cb9;
    rd_cycle[ 2808] = 1'b0;  wr_cycle[ 2808] = 1'b1;  addr_rom[ 2808]='h00002be0;  wr_data_rom[ 2808]='h000002f6;
    rd_cycle[ 2809] = 1'b0;  wr_cycle[ 2809] = 1'b1;  addr_rom[ 2809]='h00002be4;  wr_data_rom[ 2809]='h00001884;
    rd_cycle[ 2810] = 1'b0;  wr_cycle[ 2810] = 1'b1;  addr_rom[ 2810]='h00002be8;  wr_data_rom[ 2810]='h000018db;
    rd_cycle[ 2811] = 1'b0;  wr_cycle[ 2811] = 1'b1;  addr_rom[ 2811]='h00002bec;  wr_data_rom[ 2811]='h00002fd3;
    rd_cycle[ 2812] = 1'b0;  wr_cycle[ 2812] = 1'b1;  addr_rom[ 2812]='h00002bf0;  wr_data_rom[ 2812]='h00003a47;
    rd_cycle[ 2813] = 1'b0;  wr_cycle[ 2813] = 1'b1;  addr_rom[ 2813]='h00002bf4;  wr_data_rom[ 2813]='h00002d04;
    rd_cycle[ 2814] = 1'b0;  wr_cycle[ 2814] = 1'b1;  addr_rom[ 2814]='h00002bf8;  wr_data_rom[ 2814]='h00001eb1;
    rd_cycle[ 2815] = 1'b0;  wr_cycle[ 2815] = 1'b1;  addr_rom[ 2815]='h00002bfc;  wr_data_rom[ 2815]='h00002f32;
    rd_cycle[ 2816] = 1'b0;  wr_cycle[ 2816] = 1'b1;  addr_rom[ 2816]='h00002c00;  wr_data_rom[ 2816]='h00000f14;
    rd_cycle[ 2817] = 1'b0;  wr_cycle[ 2817] = 1'b1;  addr_rom[ 2817]='h00002c04;  wr_data_rom[ 2817]='h0000337a;
    rd_cycle[ 2818] = 1'b0;  wr_cycle[ 2818] = 1'b1;  addr_rom[ 2818]='h00002c08;  wr_data_rom[ 2818]='h00000a55;
    rd_cycle[ 2819] = 1'b0;  wr_cycle[ 2819] = 1'b1;  addr_rom[ 2819]='h00002c0c;  wr_data_rom[ 2819]='h00001903;
    rd_cycle[ 2820] = 1'b0;  wr_cycle[ 2820] = 1'b1;  addr_rom[ 2820]='h00002c10;  wr_data_rom[ 2820]='h0000150f;
    rd_cycle[ 2821] = 1'b0;  wr_cycle[ 2821] = 1'b1;  addr_rom[ 2821]='h00002c14;  wr_data_rom[ 2821]='h0000118b;
    rd_cycle[ 2822] = 1'b0;  wr_cycle[ 2822] = 1'b1;  addr_rom[ 2822]='h00002c18;  wr_data_rom[ 2822]='h00003532;
    rd_cycle[ 2823] = 1'b0;  wr_cycle[ 2823] = 1'b1;  addr_rom[ 2823]='h00002c1c;  wr_data_rom[ 2823]='h000024f4;
    rd_cycle[ 2824] = 1'b0;  wr_cycle[ 2824] = 1'b1;  addr_rom[ 2824]='h00002c20;  wr_data_rom[ 2824]='h00003db4;
    rd_cycle[ 2825] = 1'b0;  wr_cycle[ 2825] = 1'b1;  addr_rom[ 2825]='h00002c24;  wr_data_rom[ 2825]='h00003365;
    rd_cycle[ 2826] = 1'b0;  wr_cycle[ 2826] = 1'b1;  addr_rom[ 2826]='h00002c28;  wr_data_rom[ 2826]='h00003c9f;
    rd_cycle[ 2827] = 1'b0;  wr_cycle[ 2827] = 1'b1;  addr_rom[ 2827]='h00002c2c;  wr_data_rom[ 2827]='h0000262f;
    rd_cycle[ 2828] = 1'b0;  wr_cycle[ 2828] = 1'b1;  addr_rom[ 2828]='h00002c30;  wr_data_rom[ 2828]='h00003530;
    rd_cycle[ 2829] = 1'b0;  wr_cycle[ 2829] = 1'b1;  addr_rom[ 2829]='h00002c34;  wr_data_rom[ 2829]='h00002334;
    rd_cycle[ 2830] = 1'b0;  wr_cycle[ 2830] = 1'b1;  addr_rom[ 2830]='h00002c38;  wr_data_rom[ 2830]='h0000091c;
    rd_cycle[ 2831] = 1'b0;  wr_cycle[ 2831] = 1'b1;  addr_rom[ 2831]='h00002c3c;  wr_data_rom[ 2831]='h00000dd9;
    rd_cycle[ 2832] = 1'b0;  wr_cycle[ 2832] = 1'b1;  addr_rom[ 2832]='h00002c40;  wr_data_rom[ 2832]='h00002df3;
    rd_cycle[ 2833] = 1'b0;  wr_cycle[ 2833] = 1'b1;  addr_rom[ 2833]='h00002c44;  wr_data_rom[ 2833]='h0000315d;
    rd_cycle[ 2834] = 1'b0;  wr_cycle[ 2834] = 1'b1;  addr_rom[ 2834]='h00002c48;  wr_data_rom[ 2834]='h0000078b;
    rd_cycle[ 2835] = 1'b0;  wr_cycle[ 2835] = 1'b1;  addr_rom[ 2835]='h00002c4c;  wr_data_rom[ 2835]='h00000b00;
    rd_cycle[ 2836] = 1'b0;  wr_cycle[ 2836] = 1'b1;  addr_rom[ 2836]='h00002c50;  wr_data_rom[ 2836]='h00000bba;
    rd_cycle[ 2837] = 1'b0;  wr_cycle[ 2837] = 1'b1;  addr_rom[ 2837]='h00002c54;  wr_data_rom[ 2837]='h00002e46;
    rd_cycle[ 2838] = 1'b0;  wr_cycle[ 2838] = 1'b1;  addr_rom[ 2838]='h00002c58;  wr_data_rom[ 2838]='h00001fa2;
    rd_cycle[ 2839] = 1'b0;  wr_cycle[ 2839] = 1'b1;  addr_rom[ 2839]='h00002c5c;  wr_data_rom[ 2839]='h00003ac4;
    rd_cycle[ 2840] = 1'b0;  wr_cycle[ 2840] = 1'b1;  addr_rom[ 2840]='h00002c60;  wr_data_rom[ 2840]='h000016e2;
    rd_cycle[ 2841] = 1'b0;  wr_cycle[ 2841] = 1'b1;  addr_rom[ 2841]='h00002c64;  wr_data_rom[ 2841]='h00001869;
    rd_cycle[ 2842] = 1'b0;  wr_cycle[ 2842] = 1'b1;  addr_rom[ 2842]='h00002c68;  wr_data_rom[ 2842]='h0000299a;
    rd_cycle[ 2843] = 1'b0;  wr_cycle[ 2843] = 1'b1;  addr_rom[ 2843]='h00002c6c;  wr_data_rom[ 2843]='h00000136;
    rd_cycle[ 2844] = 1'b0;  wr_cycle[ 2844] = 1'b1;  addr_rom[ 2844]='h00002c70;  wr_data_rom[ 2844]='h000016c0;
    rd_cycle[ 2845] = 1'b0;  wr_cycle[ 2845] = 1'b1;  addr_rom[ 2845]='h00002c74;  wr_data_rom[ 2845]='h000020f2;
    rd_cycle[ 2846] = 1'b0;  wr_cycle[ 2846] = 1'b1;  addr_rom[ 2846]='h00002c78;  wr_data_rom[ 2846]='h00000c5f;
    rd_cycle[ 2847] = 1'b0;  wr_cycle[ 2847] = 1'b1;  addr_rom[ 2847]='h00002c7c;  wr_data_rom[ 2847]='h000023c7;
    rd_cycle[ 2848] = 1'b0;  wr_cycle[ 2848] = 1'b1;  addr_rom[ 2848]='h00002c80;  wr_data_rom[ 2848]='h00001229;
    rd_cycle[ 2849] = 1'b0;  wr_cycle[ 2849] = 1'b1;  addr_rom[ 2849]='h00002c84;  wr_data_rom[ 2849]='h00003acf;
    rd_cycle[ 2850] = 1'b0;  wr_cycle[ 2850] = 1'b1;  addr_rom[ 2850]='h00002c88;  wr_data_rom[ 2850]='h00001f43;
    rd_cycle[ 2851] = 1'b0;  wr_cycle[ 2851] = 1'b1;  addr_rom[ 2851]='h00002c8c;  wr_data_rom[ 2851]='h0000234b;
    rd_cycle[ 2852] = 1'b0;  wr_cycle[ 2852] = 1'b1;  addr_rom[ 2852]='h00002c90;  wr_data_rom[ 2852]='h0000002e;
    rd_cycle[ 2853] = 1'b0;  wr_cycle[ 2853] = 1'b1;  addr_rom[ 2853]='h00002c94;  wr_data_rom[ 2853]='h000019ba;
    rd_cycle[ 2854] = 1'b0;  wr_cycle[ 2854] = 1'b1;  addr_rom[ 2854]='h00002c98;  wr_data_rom[ 2854]='h00000ae0;
    rd_cycle[ 2855] = 1'b0;  wr_cycle[ 2855] = 1'b1;  addr_rom[ 2855]='h00002c9c;  wr_data_rom[ 2855]='h00003d9c;
    rd_cycle[ 2856] = 1'b0;  wr_cycle[ 2856] = 1'b1;  addr_rom[ 2856]='h00002ca0;  wr_data_rom[ 2856]='h00003d2b;
    rd_cycle[ 2857] = 1'b0;  wr_cycle[ 2857] = 1'b1;  addr_rom[ 2857]='h00002ca4;  wr_data_rom[ 2857]='h000025f2;
    rd_cycle[ 2858] = 1'b0;  wr_cycle[ 2858] = 1'b1;  addr_rom[ 2858]='h00002ca8;  wr_data_rom[ 2858]='h000017de;
    rd_cycle[ 2859] = 1'b0;  wr_cycle[ 2859] = 1'b1;  addr_rom[ 2859]='h00002cac;  wr_data_rom[ 2859]='h00000fe4;
    rd_cycle[ 2860] = 1'b0;  wr_cycle[ 2860] = 1'b1;  addr_rom[ 2860]='h00002cb0;  wr_data_rom[ 2860]='h00001d32;
    rd_cycle[ 2861] = 1'b0;  wr_cycle[ 2861] = 1'b1;  addr_rom[ 2861]='h00002cb4;  wr_data_rom[ 2861]='h00003996;
    rd_cycle[ 2862] = 1'b0;  wr_cycle[ 2862] = 1'b1;  addr_rom[ 2862]='h00002cb8;  wr_data_rom[ 2862]='h00003967;
    rd_cycle[ 2863] = 1'b0;  wr_cycle[ 2863] = 1'b1;  addr_rom[ 2863]='h00002cbc;  wr_data_rom[ 2863]='h00002abd;
    rd_cycle[ 2864] = 1'b0;  wr_cycle[ 2864] = 1'b1;  addr_rom[ 2864]='h00002cc0;  wr_data_rom[ 2864]='h00000380;
    rd_cycle[ 2865] = 1'b0;  wr_cycle[ 2865] = 1'b1;  addr_rom[ 2865]='h00002cc4;  wr_data_rom[ 2865]='h0000219c;
    rd_cycle[ 2866] = 1'b0;  wr_cycle[ 2866] = 1'b1;  addr_rom[ 2866]='h00002cc8;  wr_data_rom[ 2866]='h000011cd;
    rd_cycle[ 2867] = 1'b0;  wr_cycle[ 2867] = 1'b1;  addr_rom[ 2867]='h00002ccc;  wr_data_rom[ 2867]='h0000143c;
    rd_cycle[ 2868] = 1'b0;  wr_cycle[ 2868] = 1'b1;  addr_rom[ 2868]='h00002cd0;  wr_data_rom[ 2868]='h0000111e;
    rd_cycle[ 2869] = 1'b0;  wr_cycle[ 2869] = 1'b1;  addr_rom[ 2869]='h00002cd4;  wr_data_rom[ 2869]='h00003648;
    rd_cycle[ 2870] = 1'b0;  wr_cycle[ 2870] = 1'b1;  addr_rom[ 2870]='h00002cd8;  wr_data_rom[ 2870]='h00000e49;
    rd_cycle[ 2871] = 1'b0;  wr_cycle[ 2871] = 1'b1;  addr_rom[ 2871]='h00002cdc;  wr_data_rom[ 2871]='h00001d67;
    rd_cycle[ 2872] = 1'b0;  wr_cycle[ 2872] = 1'b1;  addr_rom[ 2872]='h00002ce0;  wr_data_rom[ 2872]='h00000bf4;
    rd_cycle[ 2873] = 1'b0;  wr_cycle[ 2873] = 1'b1;  addr_rom[ 2873]='h00002ce4;  wr_data_rom[ 2873]='h000018b0;
    rd_cycle[ 2874] = 1'b0;  wr_cycle[ 2874] = 1'b1;  addr_rom[ 2874]='h00002ce8;  wr_data_rom[ 2874]='h0000122b;
    rd_cycle[ 2875] = 1'b0;  wr_cycle[ 2875] = 1'b1;  addr_rom[ 2875]='h00002cec;  wr_data_rom[ 2875]='h000024c8;
    rd_cycle[ 2876] = 1'b0;  wr_cycle[ 2876] = 1'b1;  addr_rom[ 2876]='h00002cf0;  wr_data_rom[ 2876]='h000011a5;
    rd_cycle[ 2877] = 1'b0;  wr_cycle[ 2877] = 1'b1;  addr_rom[ 2877]='h00002cf4;  wr_data_rom[ 2877]='h0000120b;
    rd_cycle[ 2878] = 1'b0;  wr_cycle[ 2878] = 1'b1;  addr_rom[ 2878]='h00002cf8;  wr_data_rom[ 2878]='h00003c89;
    rd_cycle[ 2879] = 1'b0;  wr_cycle[ 2879] = 1'b1;  addr_rom[ 2879]='h00002cfc;  wr_data_rom[ 2879]='h00000ab9;
    rd_cycle[ 2880] = 1'b0;  wr_cycle[ 2880] = 1'b1;  addr_rom[ 2880]='h00002d00;  wr_data_rom[ 2880]='h0000383f;
    rd_cycle[ 2881] = 1'b0;  wr_cycle[ 2881] = 1'b1;  addr_rom[ 2881]='h00002d04;  wr_data_rom[ 2881]='h00001a55;
    rd_cycle[ 2882] = 1'b0;  wr_cycle[ 2882] = 1'b1;  addr_rom[ 2882]='h00002d08;  wr_data_rom[ 2882]='h00000c8b;
    rd_cycle[ 2883] = 1'b0;  wr_cycle[ 2883] = 1'b1;  addr_rom[ 2883]='h00002d0c;  wr_data_rom[ 2883]='h00003f0f;
    rd_cycle[ 2884] = 1'b0;  wr_cycle[ 2884] = 1'b1;  addr_rom[ 2884]='h00002d10;  wr_data_rom[ 2884]='h00001ba2;
    rd_cycle[ 2885] = 1'b0;  wr_cycle[ 2885] = 1'b1;  addr_rom[ 2885]='h00002d14;  wr_data_rom[ 2885]='h00001f10;
    rd_cycle[ 2886] = 1'b0;  wr_cycle[ 2886] = 1'b1;  addr_rom[ 2886]='h00002d18;  wr_data_rom[ 2886]='h00000a9d;
    rd_cycle[ 2887] = 1'b0;  wr_cycle[ 2887] = 1'b1;  addr_rom[ 2887]='h00002d1c;  wr_data_rom[ 2887]='h000022da;
    rd_cycle[ 2888] = 1'b0;  wr_cycle[ 2888] = 1'b1;  addr_rom[ 2888]='h00002d20;  wr_data_rom[ 2888]='h00001c0e;
    rd_cycle[ 2889] = 1'b0;  wr_cycle[ 2889] = 1'b1;  addr_rom[ 2889]='h00002d24;  wr_data_rom[ 2889]='h00000215;
    rd_cycle[ 2890] = 1'b0;  wr_cycle[ 2890] = 1'b1;  addr_rom[ 2890]='h00002d28;  wr_data_rom[ 2890]='h00003c9d;
    rd_cycle[ 2891] = 1'b0;  wr_cycle[ 2891] = 1'b1;  addr_rom[ 2891]='h00002d2c;  wr_data_rom[ 2891]='h00000c7f;
    rd_cycle[ 2892] = 1'b0;  wr_cycle[ 2892] = 1'b1;  addr_rom[ 2892]='h00002d30;  wr_data_rom[ 2892]='h000008c8;
    rd_cycle[ 2893] = 1'b0;  wr_cycle[ 2893] = 1'b1;  addr_rom[ 2893]='h00002d34;  wr_data_rom[ 2893]='h00002593;
    rd_cycle[ 2894] = 1'b0;  wr_cycle[ 2894] = 1'b1;  addr_rom[ 2894]='h00002d38;  wr_data_rom[ 2894]='h00003d92;
    rd_cycle[ 2895] = 1'b0;  wr_cycle[ 2895] = 1'b1;  addr_rom[ 2895]='h00002d3c;  wr_data_rom[ 2895]='h00000758;
    rd_cycle[ 2896] = 1'b0;  wr_cycle[ 2896] = 1'b1;  addr_rom[ 2896]='h00002d40;  wr_data_rom[ 2896]='h0000158b;
    rd_cycle[ 2897] = 1'b0;  wr_cycle[ 2897] = 1'b1;  addr_rom[ 2897]='h00002d44;  wr_data_rom[ 2897]='h000033ba;
    rd_cycle[ 2898] = 1'b0;  wr_cycle[ 2898] = 1'b1;  addr_rom[ 2898]='h00002d48;  wr_data_rom[ 2898]='h000005b5;
    rd_cycle[ 2899] = 1'b0;  wr_cycle[ 2899] = 1'b1;  addr_rom[ 2899]='h00002d4c;  wr_data_rom[ 2899]='h000020de;
    rd_cycle[ 2900] = 1'b0;  wr_cycle[ 2900] = 1'b1;  addr_rom[ 2900]='h00002d50;  wr_data_rom[ 2900]='h0000071c;
    rd_cycle[ 2901] = 1'b0;  wr_cycle[ 2901] = 1'b1;  addr_rom[ 2901]='h00002d54;  wr_data_rom[ 2901]='h000029e3;
    rd_cycle[ 2902] = 1'b0;  wr_cycle[ 2902] = 1'b1;  addr_rom[ 2902]='h00002d58;  wr_data_rom[ 2902]='h00000c0c;
    rd_cycle[ 2903] = 1'b0;  wr_cycle[ 2903] = 1'b1;  addr_rom[ 2903]='h00002d5c;  wr_data_rom[ 2903]='h00000e2f;
    rd_cycle[ 2904] = 1'b0;  wr_cycle[ 2904] = 1'b1;  addr_rom[ 2904]='h00002d60;  wr_data_rom[ 2904]='h00000502;
    rd_cycle[ 2905] = 1'b0;  wr_cycle[ 2905] = 1'b1;  addr_rom[ 2905]='h00002d64;  wr_data_rom[ 2905]='h00001488;
    rd_cycle[ 2906] = 1'b0;  wr_cycle[ 2906] = 1'b1;  addr_rom[ 2906]='h00002d68;  wr_data_rom[ 2906]='h00000d16;
    rd_cycle[ 2907] = 1'b0;  wr_cycle[ 2907] = 1'b1;  addr_rom[ 2907]='h00002d6c;  wr_data_rom[ 2907]='h00001527;
    rd_cycle[ 2908] = 1'b0;  wr_cycle[ 2908] = 1'b1;  addr_rom[ 2908]='h00002d70;  wr_data_rom[ 2908]='h0000170d;
    rd_cycle[ 2909] = 1'b0;  wr_cycle[ 2909] = 1'b1;  addr_rom[ 2909]='h00002d74;  wr_data_rom[ 2909]='h00002d68;
    rd_cycle[ 2910] = 1'b0;  wr_cycle[ 2910] = 1'b1;  addr_rom[ 2910]='h00002d78;  wr_data_rom[ 2910]='h000024ee;
    rd_cycle[ 2911] = 1'b0;  wr_cycle[ 2911] = 1'b1;  addr_rom[ 2911]='h00002d7c;  wr_data_rom[ 2911]='h00003389;
    rd_cycle[ 2912] = 1'b0;  wr_cycle[ 2912] = 1'b1;  addr_rom[ 2912]='h00002d80;  wr_data_rom[ 2912]='h000028db;
    rd_cycle[ 2913] = 1'b0;  wr_cycle[ 2913] = 1'b1;  addr_rom[ 2913]='h00002d84;  wr_data_rom[ 2913]='h000023ff;
    rd_cycle[ 2914] = 1'b0;  wr_cycle[ 2914] = 1'b1;  addr_rom[ 2914]='h00002d88;  wr_data_rom[ 2914]='h00003379;
    rd_cycle[ 2915] = 1'b0;  wr_cycle[ 2915] = 1'b1;  addr_rom[ 2915]='h00002d8c;  wr_data_rom[ 2915]='h0000375f;
    rd_cycle[ 2916] = 1'b0;  wr_cycle[ 2916] = 1'b1;  addr_rom[ 2916]='h00002d90;  wr_data_rom[ 2916]='h000011e9;
    rd_cycle[ 2917] = 1'b0;  wr_cycle[ 2917] = 1'b1;  addr_rom[ 2917]='h00002d94;  wr_data_rom[ 2917]='h00000059;
    rd_cycle[ 2918] = 1'b0;  wr_cycle[ 2918] = 1'b1;  addr_rom[ 2918]='h00002d98;  wr_data_rom[ 2918]='h0000346d;
    rd_cycle[ 2919] = 1'b0;  wr_cycle[ 2919] = 1'b1;  addr_rom[ 2919]='h00002d9c;  wr_data_rom[ 2919]='h000039b1;
    rd_cycle[ 2920] = 1'b0;  wr_cycle[ 2920] = 1'b1;  addr_rom[ 2920]='h00002da0;  wr_data_rom[ 2920]='h00001f57;
    rd_cycle[ 2921] = 1'b0;  wr_cycle[ 2921] = 1'b1;  addr_rom[ 2921]='h00002da4;  wr_data_rom[ 2921]='h000024c4;
    rd_cycle[ 2922] = 1'b0;  wr_cycle[ 2922] = 1'b1;  addr_rom[ 2922]='h00002da8;  wr_data_rom[ 2922]='h0000265c;
    rd_cycle[ 2923] = 1'b0;  wr_cycle[ 2923] = 1'b1;  addr_rom[ 2923]='h00002dac;  wr_data_rom[ 2923]='h0000374a;
    rd_cycle[ 2924] = 1'b0;  wr_cycle[ 2924] = 1'b1;  addr_rom[ 2924]='h00002db0;  wr_data_rom[ 2924]='h00002182;
    rd_cycle[ 2925] = 1'b0;  wr_cycle[ 2925] = 1'b1;  addr_rom[ 2925]='h00002db4;  wr_data_rom[ 2925]='h0000079c;
    rd_cycle[ 2926] = 1'b0;  wr_cycle[ 2926] = 1'b1;  addr_rom[ 2926]='h00002db8;  wr_data_rom[ 2926]='h0000204b;
    rd_cycle[ 2927] = 1'b0;  wr_cycle[ 2927] = 1'b1;  addr_rom[ 2927]='h00002dbc;  wr_data_rom[ 2927]='h00003115;
    rd_cycle[ 2928] = 1'b0;  wr_cycle[ 2928] = 1'b1;  addr_rom[ 2928]='h00002dc0;  wr_data_rom[ 2928]='h00001587;
    rd_cycle[ 2929] = 1'b0;  wr_cycle[ 2929] = 1'b1;  addr_rom[ 2929]='h00002dc4;  wr_data_rom[ 2929]='h000025d5;
    rd_cycle[ 2930] = 1'b0;  wr_cycle[ 2930] = 1'b1;  addr_rom[ 2930]='h00002dc8;  wr_data_rom[ 2930]='h000005ce;
    rd_cycle[ 2931] = 1'b0;  wr_cycle[ 2931] = 1'b1;  addr_rom[ 2931]='h00002dcc;  wr_data_rom[ 2931]='h00000a5e;
    rd_cycle[ 2932] = 1'b0;  wr_cycle[ 2932] = 1'b1;  addr_rom[ 2932]='h00002dd0;  wr_data_rom[ 2932]='h0000014a;
    rd_cycle[ 2933] = 1'b0;  wr_cycle[ 2933] = 1'b1;  addr_rom[ 2933]='h00002dd4;  wr_data_rom[ 2933]='h000017e9;
    rd_cycle[ 2934] = 1'b0;  wr_cycle[ 2934] = 1'b1;  addr_rom[ 2934]='h00002dd8;  wr_data_rom[ 2934]='h00000012;
    rd_cycle[ 2935] = 1'b0;  wr_cycle[ 2935] = 1'b1;  addr_rom[ 2935]='h00002ddc;  wr_data_rom[ 2935]='h000023d2;
    rd_cycle[ 2936] = 1'b0;  wr_cycle[ 2936] = 1'b1;  addr_rom[ 2936]='h00002de0;  wr_data_rom[ 2936]='h000027ef;
    rd_cycle[ 2937] = 1'b0;  wr_cycle[ 2937] = 1'b1;  addr_rom[ 2937]='h00002de4;  wr_data_rom[ 2937]='h000032f8;
    rd_cycle[ 2938] = 1'b0;  wr_cycle[ 2938] = 1'b1;  addr_rom[ 2938]='h00002de8;  wr_data_rom[ 2938]='h00001842;
    rd_cycle[ 2939] = 1'b0;  wr_cycle[ 2939] = 1'b1;  addr_rom[ 2939]='h00002dec;  wr_data_rom[ 2939]='h00001777;
    rd_cycle[ 2940] = 1'b0;  wr_cycle[ 2940] = 1'b1;  addr_rom[ 2940]='h00002df0;  wr_data_rom[ 2940]='h00003a83;
    rd_cycle[ 2941] = 1'b0;  wr_cycle[ 2941] = 1'b1;  addr_rom[ 2941]='h00002df4;  wr_data_rom[ 2941]='h0000220c;
    rd_cycle[ 2942] = 1'b0;  wr_cycle[ 2942] = 1'b1;  addr_rom[ 2942]='h00002df8;  wr_data_rom[ 2942]='h00002b13;
    rd_cycle[ 2943] = 1'b0;  wr_cycle[ 2943] = 1'b1;  addr_rom[ 2943]='h00002dfc;  wr_data_rom[ 2943]='h000020a3;
    rd_cycle[ 2944] = 1'b0;  wr_cycle[ 2944] = 1'b1;  addr_rom[ 2944]='h00002e00;  wr_data_rom[ 2944]='h00003c73;
    rd_cycle[ 2945] = 1'b0;  wr_cycle[ 2945] = 1'b1;  addr_rom[ 2945]='h00002e04;  wr_data_rom[ 2945]='h00002b3d;
    rd_cycle[ 2946] = 1'b0;  wr_cycle[ 2946] = 1'b1;  addr_rom[ 2946]='h00002e08;  wr_data_rom[ 2946]='h000005b0;
    rd_cycle[ 2947] = 1'b0;  wr_cycle[ 2947] = 1'b1;  addr_rom[ 2947]='h00002e0c;  wr_data_rom[ 2947]='h0000189e;
    rd_cycle[ 2948] = 1'b0;  wr_cycle[ 2948] = 1'b1;  addr_rom[ 2948]='h00002e10;  wr_data_rom[ 2948]='h000012ff;
    rd_cycle[ 2949] = 1'b0;  wr_cycle[ 2949] = 1'b1;  addr_rom[ 2949]='h00002e14;  wr_data_rom[ 2949]='h0000148b;
    rd_cycle[ 2950] = 1'b0;  wr_cycle[ 2950] = 1'b1;  addr_rom[ 2950]='h00002e18;  wr_data_rom[ 2950]='h00000df7;
    rd_cycle[ 2951] = 1'b0;  wr_cycle[ 2951] = 1'b1;  addr_rom[ 2951]='h00002e1c;  wr_data_rom[ 2951]='h00003687;
    rd_cycle[ 2952] = 1'b0;  wr_cycle[ 2952] = 1'b1;  addr_rom[ 2952]='h00002e20;  wr_data_rom[ 2952]='h0000375b;
    rd_cycle[ 2953] = 1'b0;  wr_cycle[ 2953] = 1'b1;  addr_rom[ 2953]='h00002e24;  wr_data_rom[ 2953]='h000010a5;
    rd_cycle[ 2954] = 1'b0;  wr_cycle[ 2954] = 1'b1;  addr_rom[ 2954]='h00002e28;  wr_data_rom[ 2954]='h00001944;
    rd_cycle[ 2955] = 1'b0;  wr_cycle[ 2955] = 1'b1;  addr_rom[ 2955]='h00002e2c;  wr_data_rom[ 2955]='h00002f30;
    rd_cycle[ 2956] = 1'b0;  wr_cycle[ 2956] = 1'b1;  addr_rom[ 2956]='h00002e30;  wr_data_rom[ 2956]='h00002c4f;
    rd_cycle[ 2957] = 1'b0;  wr_cycle[ 2957] = 1'b1;  addr_rom[ 2957]='h00002e34;  wr_data_rom[ 2957]='h00003213;
    rd_cycle[ 2958] = 1'b0;  wr_cycle[ 2958] = 1'b1;  addr_rom[ 2958]='h00002e38;  wr_data_rom[ 2958]='h00001e27;
    rd_cycle[ 2959] = 1'b0;  wr_cycle[ 2959] = 1'b1;  addr_rom[ 2959]='h00002e3c;  wr_data_rom[ 2959]='h00002883;
    rd_cycle[ 2960] = 1'b0;  wr_cycle[ 2960] = 1'b1;  addr_rom[ 2960]='h00002e40;  wr_data_rom[ 2960]='h000035a1;
    rd_cycle[ 2961] = 1'b0;  wr_cycle[ 2961] = 1'b1;  addr_rom[ 2961]='h00002e44;  wr_data_rom[ 2961]='h000031c7;
    rd_cycle[ 2962] = 1'b0;  wr_cycle[ 2962] = 1'b1;  addr_rom[ 2962]='h00002e48;  wr_data_rom[ 2962]='h000026cb;
    rd_cycle[ 2963] = 1'b0;  wr_cycle[ 2963] = 1'b1;  addr_rom[ 2963]='h00002e4c;  wr_data_rom[ 2963]='h0000109a;
    rd_cycle[ 2964] = 1'b0;  wr_cycle[ 2964] = 1'b1;  addr_rom[ 2964]='h00002e50;  wr_data_rom[ 2964]='h000029c0;
    rd_cycle[ 2965] = 1'b0;  wr_cycle[ 2965] = 1'b1;  addr_rom[ 2965]='h00002e54;  wr_data_rom[ 2965]='h00001fd1;
    rd_cycle[ 2966] = 1'b0;  wr_cycle[ 2966] = 1'b1;  addr_rom[ 2966]='h00002e58;  wr_data_rom[ 2966]='h000015d9;
    rd_cycle[ 2967] = 1'b0;  wr_cycle[ 2967] = 1'b1;  addr_rom[ 2967]='h00002e5c;  wr_data_rom[ 2967]='h00001f20;
    rd_cycle[ 2968] = 1'b0;  wr_cycle[ 2968] = 1'b1;  addr_rom[ 2968]='h00002e60;  wr_data_rom[ 2968]='h000000f8;
    rd_cycle[ 2969] = 1'b0;  wr_cycle[ 2969] = 1'b1;  addr_rom[ 2969]='h00002e64;  wr_data_rom[ 2969]='h00003e04;
    rd_cycle[ 2970] = 1'b0;  wr_cycle[ 2970] = 1'b1;  addr_rom[ 2970]='h00002e68;  wr_data_rom[ 2970]='h000035e6;
    rd_cycle[ 2971] = 1'b0;  wr_cycle[ 2971] = 1'b1;  addr_rom[ 2971]='h00002e6c;  wr_data_rom[ 2971]='h000035c0;
    rd_cycle[ 2972] = 1'b0;  wr_cycle[ 2972] = 1'b1;  addr_rom[ 2972]='h00002e70;  wr_data_rom[ 2972]='h00000732;
    rd_cycle[ 2973] = 1'b0;  wr_cycle[ 2973] = 1'b1;  addr_rom[ 2973]='h00002e74;  wr_data_rom[ 2973]='h00003559;
    rd_cycle[ 2974] = 1'b0;  wr_cycle[ 2974] = 1'b1;  addr_rom[ 2974]='h00002e78;  wr_data_rom[ 2974]='h000006d3;
    rd_cycle[ 2975] = 1'b0;  wr_cycle[ 2975] = 1'b1;  addr_rom[ 2975]='h00002e7c;  wr_data_rom[ 2975]='h00000e09;
    rd_cycle[ 2976] = 1'b0;  wr_cycle[ 2976] = 1'b1;  addr_rom[ 2976]='h00002e80;  wr_data_rom[ 2976]='h00000c64;
    rd_cycle[ 2977] = 1'b0;  wr_cycle[ 2977] = 1'b1;  addr_rom[ 2977]='h00002e84;  wr_data_rom[ 2977]='h00002d5a;
    rd_cycle[ 2978] = 1'b0;  wr_cycle[ 2978] = 1'b1;  addr_rom[ 2978]='h00002e88;  wr_data_rom[ 2978]='h00000a3b;
    rd_cycle[ 2979] = 1'b0;  wr_cycle[ 2979] = 1'b1;  addr_rom[ 2979]='h00002e8c;  wr_data_rom[ 2979]='h00002c2d;
    rd_cycle[ 2980] = 1'b0;  wr_cycle[ 2980] = 1'b1;  addr_rom[ 2980]='h00002e90;  wr_data_rom[ 2980]='h00003f72;
    rd_cycle[ 2981] = 1'b0;  wr_cycle[ 2981] = 1'b1;  addr_rom[ 2981]='h00002e94;  wr_data_rom[ 2981]='h00002670;
    rd_cycle[ 2982] = 1'b0;  wr_cycle[ 2982] = 1'b1;  addr_rom[ 2982]='h00002e98;  wr_data_rom[ 2982]='h00000fe5;
    rd_cycle[ 2983] = 1'b0;  wr_cycle[ 2983] = 1'b1;  addr_rom[ 2983]='h00002e9c;  wr_data_rom[ 2983]='h000017d8;
    rd_cycle[ 2984] = 1'b0;  wr_cycle[ 2984] = 1'b1;  addr_rom[ 2984]='h00002ea0;  wr_data_rom[ 2984]='h000015ff;
    rd_cycle[ 2985] = 1'b0;  wr_cycle[ 2985] = 1'b1;  addr_rom[ 2985]='h00002ea4;  wr_data_rom[ 2985]='h0000049b;
    rd_cycle[ 2986] = 1'b0;  wr_cycle[ 2986] = 1'b1;  addr_rom[ 2986]='h00002ea8;  wr_data_rom[ 2986]='h0000143b;
    rd_cycle[ 2987] = 1'b0;  wr_cycle[ 2987] = 1'b1;  addr_rom[ 2987]='h00002eac;  wr_data_rom[ 2987]='h00000a0e;
    rd_cycle[ 2988] = 1'b0;  wr_cycle[ 2988] = 1'b1;  addr_rom[ 2988]='h00002eb0;  wr_data_rom[ 2988]='h00002a41;
    rd_cycle[ 2989] = 1'b0;  wr_cycle[ 2989] = 1'b1;  addr_rom[ 2989]='h00002eb4;  wr_data_rom[ 2989]='h000027e3;
    rd_cycle[ 2990] = 1'b0;  wr_cycle[ 2990] = 1'b1;  addr_rom[ 2990]='h00002eb8;  wr_data_rom[ 2990]='h00000475;
    rd_cycle[ 2991] = 1'b0;  wr_cycle[ 2991] = 1'b1;  addr_rom[ 2991]='h00002ebc;  wr_data_rom[ 2991]='h0000143d;
    rd_cycle[ 2992] = 1'b0;  wr_cycle[ 2992] = 1'b1;  addr_rom[ 2992]='h00002ec0;  wr_data_rom[ 2992]='h00001ea7;
    rd_cycle[ 2993] = 1'b0;  wr_cycle[ 2993] = 1'b1;  addr_rom[ 2993]='h00002ec4;  wr_data_rom[ 2993]='h00001d1d;
    rd_cycle[ 2994] = 1'b0;  wr_cycle[ 2994] = 1'b1;  addr_rom[ 2994]='h00002ec8;  wr_data_rom[ 2994]='h00000638;
    rd_cycle[ 2995] = 1'b0;  wr_cycle[ 2995] = 1'b1;  addr_rom[ 2995]='h00002ecc;  wr_data_rom[ 2995]='h000008d0;
    rd_cycle[ 2996] = 1'b0;  wr_cycle[ 2996] = 1'b1;  addr_rom[ 2996]='h00002ed0;  wr_data_rom[ 2996]='h00002eb9;
    rd_cycle[ 2997] = 1'b0;  wr_cycle[ 2997] = 1'b1;  addr_rom[ 2997]='h00002ed4;  wr_data_rom[ 2997]='h000006ab;
    rd_cycle[ 2998] = 1'b0;  wr_cycle[ 2998] = 1'b1;  addr_rom[ 2998]='h00002ed8;  wr_data_rom[ 2998]='h00001aef;
    rd_cycle[ 2999] = 1'b0;  wr_cycle[ 2999] = 1'b1;  addr_rom[ 2999]='h00002edc;  wr_data_rom[ 2999]='h000009ce;
    rd_cycle[ 3000] = 1'b0;  wr_cycle[ 3000] = 1'b1;  addr_rom[ 3000]='h00002ee0;  wr_data_rom[ 3000]='h00000452;
    rd_cycle[ 3001] = 1'b0;  wr_cycle[ 3001] = 1'b1;  addr_rom[ 3001]='h00002ee4;  wr_data_rom[ 3001]='h0000040b;
    rd_cycle[ 3002] = 1'b0;  wr_cycle[ 3002] = 1'b1;  addr_rom[ 3002]='h00002ee8;  wr_data_rom[ 3002]='h00000ba0;
    rd_cycle[ 3003] = 1'b0;  wr_cycle[ 3003] = 1'b1;  addr_rom[ 3003]='h00002eec;  wr_data_rom[ 3003]='h00002cbf;
    rd_cycle[ 3004] = 1'b0;  wr_cycle[ 3004] = 1'b1;  addr_rom[ 3004]='h00002ef0;  wr_data_rom[ 3004]='h000034d5;
    rd_cycle[ 3005] = 1'b0;  wr_cycle[ 3005] = 1'b1;  addr_rom[ 3005]='h00002ef4;  wr_data_rom[ 3005]='h00001a79;
    rd_cycle[ 3006] = 1'b0;  wr_cycle[ 3006] = 1'b1;  addr_rom[ 3006]='h00002ef8;  wr_data_rom[ 3006]='h00001d60;
    rd_cycle[ 3007] = 1'b0;  wr_cycle[ 3007] = 1'b1;  addr_rom[ 3007]='h00002efc;  wr_data_rom[ 3007]='h0000227a;
    rd_cycle[ 3008] = 1'b0;  wr_cycle[ 3008] = 1'b1;  addr_rom[ 3008]='h00002f00;  wr_data_rom[ 3008]='h000038df;
    rd_cycle[ 3009] = 1'b0;  wr_cycle[ 3009] = 1'b1;  addr_rom[ 3009]='h00002f04;  wr_data_rom[ 3009]='h0000369d;
    rd_cycle[ 3010] = 1'b0;  wr_cycle[ 3010] = 1'b1;  addr_rom[ 3010]='h00002f08;  wr_data_rom[ 3010]='h00003178;
    rd_cycle[ 3011] = 1'b0;  wr_cycle[ 3011] = 1'b1;  addr_rom[ 3011]='h00002f0c;  wr_data_rom[ 3011]='h0000171e;
    rd_cycle[ 3012] = 1'b0;  wr_cycle[ 3012] = 1'b1;  addr_rom[ 3012]='h00002f10;  wr_data_rom[ 3012]='h000026aa;
    rd_cycle[ 3013] = 1'b0;  wr_cycle[ 3013] = 1'b1;  addr_rom[ 3013]='h00002f14;  wr_data_rom[ 3013]='h000032da;
    rd_cycle[ 3014] = 1'b0;  wr_cycle[ 3014] = 1'b1;  addr_rom[ 3014]='h00002f18;  wr_data_rom[ 3014]='h00002a58;
    rd_cycle[ 3015] = 1'b0;  wr_cycle[ 3015] = 1'b1;  addr_rom[ 3015]='h00002f1c;  wr_data_rom[ 3015]='h000032cc;
    rd_cycle[ 3016] = 1'b0;  wr_cycle[ 3016] = 1'b1;  addr_rom[ 3016]='h00002f20;  wr_data_rom[ 3016]='h00002826;
    rd_cycle[ 3017] = 1'b0;  wr_cycle[ 3017] = 1'b1;  addr_rom[ 3017]='h00002f24;  wr_data_rom[ 3017]='h00002f95;
    rd_cycle[ 3018] = 1'b0;  wr_cycle[ 3018] = 1'b1;  addr_rom[ 3018]='h00002f28;  wr_data_rom[ 3018]='h00003727;
    rd_cycle[ 3019] = 1'b0;  wr_cycle[ 3019] = 1'b1;  addr_rom[ 3019]='h00002f2c;  wr_data_rom[ 3019]='h00000e76;
    rd_cycle[ 3020] = 1'b0;  wr_cycle[ 3020] = 1'b1;  addr_rom[ 3020]='h00002f30;  wr_data_rom[ 3020]='h000018e5;
    rd_cycle[ 3021] = 1'b0;  wr_cycle[ 3021] = 1'b1;  addr_rom[ 3021]='h00002f34;  wr_data_rom[ 3021]='h00002c73;
    rd_cycle[ 3022] = 1'b0;  wr_cycle[ 3022] = 1'b1;  addr_rom[ 3022]='h00002f38;  wr_data_rom[ 3022]='h0000225c;
    rd_cycle[ 3023] = 1'b0;  wr_cycle[ 3023] = 1'b1;  addr_rom[ 3023]='h00002f3c;  wr_data_rom[ 3023]='h00003b26;
    rd_cycle[ 3024] = 1'b0;  wr_cycle[ 3024] = 1'b1;  addr_rom[ 3024]='h00002f40;  wr_data_rom[ 3024]='h00003303;
    rd_cycle[ 3025] = 1'b0;  wr_cycle[ 3025] = 1'b1;  addr_rom[ 3025]='h00002f44;  wr_data_rom[ 3025]='h000007a0;
    rd_cycle[ 3026] = 1'b0;  wr_cycle[ 3026] = 1'b1;  addr_rom[ 3026]='h00002f48;  wr_data_rom[ 3026]='h000004e5;
    rd_cycle[ 3027] = 1'b0;  wr_cycle[ 3027] = 1'b1;  addr_rom[ 3027]='h00002f4c;  wr_data_rom[ 3027]='h00001c92;
    rd_cycle[ 3028] = 1'b0;  wr_cycle[ 3028] = 1'b1;  addr_rom[ 3028]='h00002f50;  wr_data_rom[ 3028]='h00002c38;
    rd_cycle[ 3029] = 1'b0;  wr_cycle[ 3029] = 1'b1;  addr_rom[ 3029]='h00002f54;  wr_data_rom[ 3029]='h0000380f;
    rd_cycle[ 3030] = 1'b0;  wr_cycle[ 3030] = 1'b1;  addr_rom[ 3030]='h00002f58;  wr_data_rom[ 3030]='h000025a0;
    rd_cycle[ 3031] = 1'b0;  wr_cycle[ 3031] = 1'b1;  addr_rom[ 3031]='h00002f5c;  wr_data_rom[ 3031]='h0000359e;
    rd_cycle[ 3032] = 1'b0;  wr_cycle[ 3032] = 1'b1;  addr_rom[ 3032]='h00002f60;  wr_data_rom[ 3032]='h0000308d;
    rd_cycle[ 3033] = 1'b0;  wr_cycle[ 3033] = 1'b1;  addr_rom[ 3033]='h00002f64;  wr_data_rom[ 3033]='h000022e1;
    rd_cycle[ 3034] = 1'b0;  wr_cycle[ 3034] = 1'b1;  addr_rom[ 3034]='h00002f68;  wr_data_rom[ 3034]='h000020ed;
    rd_cycle[ 3035] = 1'b0;  wr_cycle[ 3035] = 1'b1;  addr_rom[ 3035]='h00002f6c;  wr_data_rom[ 3035]='h00002e41;
    rd_cycle[ 3036] = 1'b0;  wr_cycle[ 3036] = 1'b1;  addr_rom[ 3036]='h00002f70;  wr_data_rom[ 3036]='h00003ce8;
    rd_cycle[ 3037] = 1'b0;  wr_cycle[ 3037] = 1'b1;  addr_rom[ 3037]='h00002f74;  wr_data_rom[ 3037]='h0000132b;
    rd_cycle[ 3038] = 1'b0;  wr_cycle[ 3038] = 1'b1;  addr_rom[ 3038]='h00002f78;  wr_data_rom[ 3038]='h000001ae;
    rd_cycle[ 3039] = 1'b0;  wr_cycle[ 3039] = 1'b1;  addr_rom[ 3039]='h00002f7c;  wr_data_rom[ 3039]='h0000011e;
    rd_cycle[ 3040] = 1'b0;  wr_cycle[ 3040] = 1'b1;  addr_rom[ 3040]='h00002f80;  wr_data_rom[ 3040]='h00003a4f;
    rd_cycle[ 3041] = 1'b0;  wr_cycle[ 3041] = 1'b1;  addr_rom[ 3041]='h00002f84;  wr_data_rom[ 3041]='h000033ef;
    rd_cycle[ 3042] = 1'b0;  wr_cycle[ 3042] = 1'b1;  addr_rom[ 3042]='h00002f88;  wr_data_rom[ 3042]='h00001bfc;
    rd_cycle[ 3043] = 1'b0;  wr_cycle[ 3043] = 1'b1;  addr_rom[ 3043]='h00002f8c;  wr_data_rom[ 3043]='h00000552;
    rd_cycle[ 3044] = 1'b0;  wr_cycle[ 3044] = 1'b1;  addr_rom[ 3044]='h00002f90;  wr_data_rom[ 3044]='h0000145a;
    rd_cycle[ 3045] = 1'b0;  wr_cycle[ 3045] = 1'b1;  addr_rom[ 3045]='h00002f94;  wr_data_rom[ 3045]='h00000e83;
    rd_cycle[ 3046] = 1'b0;  wr_cycle[ 3046] = 1'b1;  addr_rom[ 3046]='h00002f98;  wr_data_rom[ 3046]='h00000f23;
    rd_cycle[ 3047] = 1'b0;  wr_cycle[ 3047] = 1'b1;  addr_rom[ 3047]='h00002f9c;  wr_data_rom[ 3047]='h0000295c;
    rd_cycle[ 3048] = 1'b0;  wr_cycle[ 3048] = 1'b1;  addr_rom[ 3048]='h00002fa0;  wr_data_rom[ 3048]='h00001c0e;
    rd_cycle[ 3049] = 1'b0;  wr_cycle[ 3049] = 1'b1;  addr_rom[ 3049]='h00002fa4;  wr_data_rom[ 3049]='h00002844;
    rd_cycle[ 3050] = 1'b0;  wr_cycle[ 3050] = 1'b1;  addr_rom[ 3050]='h00002fa8;  wr_data_rom[ 3050]='h00000a11;
    rd_cycle[ 3051] = 1'b0;  wr_cycle[ 3051] = 1'b1;  addr_rom[ 3051]='h00002fac;  wr_data_rom[ 3051]='h0000325e;
    rd_cycle[ 3052] = 1'b0;  wr_cycle[ 3052] = 1'b1;  addr_rom[ 3052]='h00002fb0;  wr_data_rom[ 3052]='h000026de;
    rd_cycle[ 3053] = 1'b0;  wr_cycle[ 3053] = 1'b1;  addr_rom[ 3053]='h00002fb4;  wr_data_rom[ 3053]='h00002064;
    rd_cycle[ 3054] = 1'b0;  wr_cycle[ 3054] = 1'b1;  addr_rom[ 3054]='h00002fb8;  wr_data_rom[ 3054]='h00002265;
    rd_cycle[ 3055] = 1'b0;  wr_cycle[ 3055] = 1'b1;  addr_rom[ 3055]='h00002fbc;  wr_data_rom[ 3055]='h00003976;
    rd_cycle[ 3056] = 1'b0;  wr_cycle[ 3056] = 1'b1;  addr_rom[ 3056]='h00002fc0;  wr_data_rom[ 3056]='h00002051;
    rd_cycle[ 3057] = 1'b0;  wr_cycle[ 3057] = 1'b1;  addr_rom[ 3057]='h00002fc4;  wr_data_rom[ 3057]='h00001069;
    rd_cycle[ 3058] = 1'b0;  wr_cycle[ 3058] = 1'b1;  addr_rom[ 3058]='h00002fc8;  wr_data_rom[ 3058]='h0000267f;
    rd_cycle[ 3059] = 1'b0;  wr_cycle[ 3059] = 1'b1;  addr_rom[ 3059]='h00002fcc;  wr_data_rom[ 3059]='h00000e65;
    rd_cycle[ 3060] = 1'b0;  wr_cycle[ 3060] = 1'b1;  addr_rom[ 3060]='h00002fd0;  wr_data_rom[ 3060]='h00001103;
    rd_cycle[ 3061] = 1'b0;  wr_cycle[ 3061] = 1'b1;  addr_rom[ 3061]='h00002fd4;  wr_data_rom[ 3061]='h00001a30;
    rd_cycle[ 3062] = 1'b0;  wr_cycle[ 3062] = 1'b1;  addr_rom[ 3062]='h00002fd8;  wr_data_rom[ 3062]='h00002361;
    rd_cycle[ 3063] = 1'b0;  wr_cycle[ 3063] = 1'b1;  addr_rom[ 3063]='h00002fdc;  wr_data_rom[ 3063]='h00000513;
    rd_cycle[ 3064] = 1'b0;  wr_cycle[ 3064] = 1'b1;  addr_rom[ 3064]='h00002fe0;  wr_data_rom[ 3064]='h00000452;
    rd_cycle[ 3065] = 1'b0;  wr_cycle[ 3065] = 1'b1;  addr_rom[ 3065]='h00002fe4;  wr_data_rom[ 3065]='h00002011;
    rd_cycle[ 3066] = 1'b0;  wr_cycle[ 3066] = 1'b1;  addr_rom[ 3066]='h00002fe8;  wr_data_rom[ 3066]='h00002343;
    rd_cycle[ 3067] = 1'b0;  wr_cycle[ 3067] = 1'b1;  addr_rom[ 3067]='h00002fec;  wr_data_rom[ 3067]='h00003d48;
    rd_cycle[ 3068] = 1'b0;  wr_cycle[ 3068] = 1'b1;  addr_rom[ 3068]='h00002ff0;  wr_data_rom[ 3068]='h000034ea;
    rd_cycle[ 3069] = 1'b0;  wr_cycle[ 3069] = 1'b1;  addr_rom[ 3069]='h00002ff4;  wr_data_rom[ 3069]='h00001fd7;
    rd_cycle[ 3070] = 1'b0;  wr_cycle[ 3070] = 1'b1;  addr_rom[ 3070]='h00002ff8;  wr_data_rom[ 3070]='h00003094;
    rd_cycle[ 3071] = 1'b0;  wr_cycle[ 3071] = 1'b1;  addr_rom[ 3071]='h00002ffc;  wr_data_rom[ 3071]='h00002012;
    rd_cycle[ 3072] = 1'b0;  wr_cycle[ 3072] = 1'b1;  addr_rom[ 3072]='h00003000;  wr_data_rom[ 3072]='h000029ea;
    rd_cycle[ 3073] = 1'b0;  wr_cycle[ 3073] = 1'b1;  addr_rom[ 3073]='h00003004;  wr_data_rom[ 3073]='h00001aa9;
    rd_cycle[ 3074] = 1'b0;  wr_cycle[ 3074] = 1'b1;  addr_rom[ 3074]='h00003008;  wr_data_rom[ 3074]='h00001205;
    rd_cycle[ 3075] = 1'b0;  wr_cycle[ 3075] = 1'b1;  addr_rom[ 3075]='h0000300c;  wr_data_rom[ 3075]='h000006a6;
    rd_cycle[ 3076] = 1'b0;  wr_cycle[ 3076] = 1'b1;  addr_rom[ 3076]='h00003010;  wr_data_rom[ 3076]='h000017a9;
    rd_cycle[ 3077] = 1'b0;  wr_cycle[ 3077] = 1'b1;  addr_rom[ 3077]='h00003014;  wr_data_rom[ 3077]='h000001a0;
    rd_cycle[ 3078] = 1'b0;  wr_cycle[ 3078] = 1'b1;  addr_rom[ 3078]='h00003018;  wr_data_rom[ 3078]='h00001329;
    rd_cycle[ 3079] = 1'b0;  wr_cycle[ 3079] = 1'b1;  addr_rom[ 3079]='h0000301c;  wr_data_rom[ 3079]='h00000d01;
    rd_cycle[ 3080] = 1'b0;  wr_cycle[ 3080] = 1'b1;  addr_rom[ 3080]='h00003020;  wr_data_rom[ 3080]='h00000ead;
    rd_cycle[ 3081] = 1'b0;  wr_cycle[ 3081] = 1'b1;  addr_rom[ 3081]='h00003024;  wr_data_rom[ 3081]='h00003e88;
    rd_cycle[ 3082] = 1'b0;  wr_cycle[ 3082] = 1'b1;  addr_rom[ 3082]='h00003028;  wr_data_rom[ 3082]='h00001a38;
    rd_cycle[ 3083] = 1'b0;  wr_cycle[ 3083] = 1'b1;  addr_rom[ 3083]='h0000302c;  wr_data_rom[ 3083]='h00000792;
    rd_cycle[ 3084] = 1'b0;  wr_cycle[ 3084] = 1'b1;  addr_rom[ 3084]='h00003030;  wr_data_rom[ 3084]='h00001962;
    rd_cycle[ 3085] = 1'b0;  wr_cycle[ 3085] = 1'b1;  addr_rom[ 3085]='h00003034;  wr_data_rom[ 3085]='h00003d3c;
    rd_cycle[ 3086] = 1'b0;  wr_cycle[ 3086] = 1'b1;  addr_rom[ 3086]='h00003038;  wr_data_rom[ 3086]='h00002588;
    rd_cycle[ 3087] = 1'b0;  wr_cycle[ 3087] = 1'b1;  addr_rom[ 3087]='h0000303c;  wr_data_rom[ 3087]='h00003bab;
    rd_cycle[ 3088] = 1'b0;  wr_cycle[ 3088] = 1'b1;  addr_rom[ 3088]='h00003040;  wr_data_rom[ 3088]='h00002144;
    rd_cycle[ 3089] = 1'b0;  wr_cycle[ 3089] = 1'b1;  addr_rom[ 3089]='h00003044;  wr_data_rom[ 3089]='h00002ab8;
    rd_cycle[ 3090] = 1'b0;  wr_cycle[ 3090] = 1'b1;  addr_rom[ 3090]='h00003048;  wr_data_rom[ 3090]='h00001ba6;
    rd_cycle[ 3091] = 1'b0;  wr_cycle[ 3091] = 1'b1;  addr_rom[ 3091]='h0000304c;  wr_data_rom[ 3091]='h00000736;
    rd_cycle[ 3092] = 1'b0;  wr_cycle[ 3092] = 1'b1;  addr_rom[ 3092]='h00003050;  wr_data_rom[ 3092]='h00001255;
    rd_cycle[ 3093] = 1'b0;  wr_cycle[ 3093] = 1'b1;  addr_rom[ 3093]='h00003054;  wr_data_rom[ 3093]='h00000525;
    rd_cycle[ 3094] = 1'b0;  wr_cycle[ 3094] = 1'b1;  addr_rom[ 3094]='h00003058;  wr_data_rom[ 3094]='h00002386;
    rd_cycle[ 3095] = 1'b0;  wr_cycle[ 3095] = 1'b1;  addr_rom[ 3095]='h0000305c;  wr_data_rom[ 3095]='h00001aab;
    rd_cycle[ 3096] = 1'b0;  wr_cycle[ 3096] = 1'b1;  addr_rom[ 3096]='h00003060;  wr_data_rom[ 3096]='h00000359;
    rd_cycle[ 3097] = 1'b0;  wr_cycle[ 3097] = 1'b1;  addr_rom[ 3097]='h00003064;  wr_data_rom[ 3097]='h00003906;
    rd_cycle[ 3098] = 1'b0;  wr_cycle[ 3098] = 1'b1;  addr_rom[ 3098]='h00003068;  wr_data_rom[ 3098]='h0000275b;
    rd_cycle[ 3099] = 1'b0;  wr_cycle[ 3099] = 1'b1;  addr_rom[ 3099]='h0000306c;  wr_data_rom[ 3099]='h00002eae;
    rd_cycle[ 3100] = 1'b0;  wr_cycle[ 3100] = 1'b1;  addr_rom[ 3100]='h00003070;  wr_data_rom[ 3100]='h00000303;
    rd_cycle[ 3101] = 1'b0;  wr_cycle[ 3101] = 1'b1;  addr_rom[ 3101]='h00003074;  wr_data_rom[ 3101]='h000021dd;
    rd_cycle[ 3102] = 1'b0;  wr_cycle[ 3102] = 1'b1;  addr_rom[ 3102]='h00003078;  wr_data_rom[ 3102]='h00002fa0;
    rd_cycle[ 3103] = 1'b0;  wr_cycle[ 3103] = 1'b1;  addr_rom[ 3103]='h0000307c;  wr_data_rom[ 3103]='h00000a2e;
    rd_cycle[ 3104] = 1'b0;  wr_cycle[ 3104] = 1'b1;  addr_rom[ 3104]='h00003080;  wr_data_rom[ 3104]='h0000000f;
    rd_cycle[ 3105] = 1'b0;  wr_cycle[ 3105] = 1'b1;  addr_rom[ 3105]='h00003084;  wr_data_rom[ 3105]='h00000e52;
    rd_cycle[ 3106] = 1'b0;  wr_cycle[ 3106] = 1'b1;  addr_rom[ 3106]='h00003088;  wr_data_rom[ 3106]='h00000bd6;
    rd_cycle[ 3107] = 1'b0;  wr_cycle[ 3107] = 1'b1;  addr_rom[ 3107]='h0000308c;  wr_data_rom[ 3107]='h00001ae8;
    rd_cycle[ 3108] = 1'b0;  wr_cycle[ 3108] = 1'b1;  addr_rom[ 3108]='h00003090;  wr_data_rom[ 3108]='h00003744;
    rd_cycle[ 3109] = 1'b0;  wr_cycle[ 3109] = 1'b1;  addr_rom[ 3109]='h00003094;  wr_data_rom[ 3109]='h00002471;
    rd_cycle[ 3110] = 1'b0;  wr_cycle[ 3110] = 1'b1;  addr_rom[ 3110]='h00003098;  wr_data_rom[ 3110]='h000017c1;
    rd_cycle[ 3111] = 1'b0;  wr_cycle[ 3111] = 1'b1;  addr_rom[ 3111]='h0000309c;  wr_data_rom[ 3111]='h00002108;
    rd_cycle[ 3112] = 1'b0;  wr_cycle[ 3112] = 1'b1;  addr_rom[ 3112]='h000030a0;  wr_data_rom[ 3112]='h00002b58;
    rd_cycle[ 3113] = 1'b0;  wr_cycle[ 3113] = 1'b1;  addr_rom[ 3113]='h000030a4;  wr_data_rom[ 3113]='h0000301f;
    rd_cycle[ 3114] = 1'b0;  wr_cycle[ 3114] = 1'b1;  addr_rom[ 3114]='h000030a8;  wr_data_rom[ 3114]='h0000354e;
    rd_cycle[ 3115] = 1'b0;  wr_cycle[ 3115] = 1'b1;  addr_rom[ 3115]='h000030ac;  wr_data_rom[ 3115]='h00000e6e;
    rd_cycle[ 3116] = 1'b0;  wr_cycle[ 3116] = 1'b1;  addr_rom[ 3116]='h000030b0;  wr_data_rom[ 3116]='h000023eb;
    rd_cycle[ 3117] = 1'b0;  wr_cycle[ 3117] = 1'b1;  addr_rom[ 3117]='h000030b4;  wr_data_rom[ 3117]='h00003326;
    rd_cycle[ 3118] = 1'b0;  wr_cycle[ 3118] = 1'b1;  addr_rom[ 3118]='h000030b8;  wr_data_rom[ 3118]='h0000041a;
    rd_cycle[ 3119] = 1'b0;  wr_cycle[ 3119] = 1'b1;  addr_rom[ 3119]='h000030bc;  wr_data_rom[ 3119]='h00001702;
    rd_cycle[ 3120] = 1'b0;  wr_cycle[ 3120] = 1'b1;  addr_rom[ 3120]='h000030c0;  wr_data_rom[ 3120]='h000015fe;
    rd_cycle[ 3121] = 1'b0;  wr_cycle[ 3121] = 1'b1;  addr_rom[ 3121]='h000030c4;  wr_data_rom[ 3121]='h00001db5;
    rd_cycle[ 3122] = 1'b0;  wr_cycle[ 3122] = 1'b1;  addr_rom[ 3122]='h000030c8;  wr_data_rom[ 3122]='h000016e1;
    rd_cycle[ 3123] = 1'b0;  wr_cycle[ 3123] = 1'b1;  addr_rom[ 3123]='h000030cc;  wr_data_rom[ 3123]='h00000cc7;
    rd_cycle[ 3124] = 1'b0;  wr_cycle[ 3124] = 1'b1;  addr_rom[ 3124]='h000030d0;  wr_data_rom[ 3124]='h00003ab1;
    rd_cycle[ 3125] = 1'b0;  wr_cycle[ 3125] = 1'b1;  addr_rom[ 3125]='h000030d4;  wr_data_rom[ 3125]='h00000ae5;
    rd_cycle[ 3126] = 1'b0;  wr_cycle[ 3126] = 1'b1;  addr_rom[ 3126]='h000030d8;  wr_data_rom[ 3126]='h00003681;
    rd_cycle[ 3127] = 1'b0;  wr_cycle[ 3127] = 1'b1;  addr_rom[ 3127]='h000030dc;  wr_data_rom[ 3127]='h000007eb;
    rd_cycle[ 3128] = 1'b0;  wr_cycle[ 3128] = 1'b1;  addr_rom[ 3128]='h000030e0;  wr_data_rom[ 3128]='h000031eb;
    rd_cycle[ 3129] = 1'b0;  wr_cycle[ 3129] = 1'b1;  addr_rom[ 3129]='h000030e4;  wr_data_rom[ 3129]='h00000a3c;
    rd_cycle[ 3130] = 1'b0;  wr_cycle[ 3130] = 1'b1;  addr_rom[ 3130]='h000030e8;  wr_data_rom[ 3130]='h00000434;
    rd_cycle[ 3131] = 1'b0;  wr_cycle[ 3131] = 1'b1;  addr_rom[ 3131]='h000030ec;  wr_data_rom[ 3131]='h000015ee;
    rd_cycle[ 3132] = 1'b0;  wr_cycle[ 3132] = 1'b1;  addr_rom[ 3132]='h000030f0;  wr_data_rom[ 3132]='h000002e6;
    rd_cycle[ 3133] = 1'b0;  wr_cycle[ 3133] = 1'b1;  addr_rom[ 3133]='h000030f4;  wr_data_rom[ 3133]='h000001b4;
    rd_cycle[ 3134] = 1'b0;  wr_cycle[ 3134] = 1'b1;  addr_rom[ 3134]='h000030f8;  wr_data_rom[ 3134]='h00003edb;
    rd_cycle[ 3135] = 1'b0;  wr_cycle[ 3135] = 1'b1;  addr_rom[ 3135]='h000030fc;  wr_data_rom[ 3135]='h000013f5;
    rd_cycle[ 3136] = 1'b0;  wr_cycle[ 3136] = 1'b1;  addr_rom[ 3136]='h00003100;  wr_data_rom[ 3136]='h0000162b;
    rd_cycle[ 3137] = 1'b0;  wr_cycle[ 3137] = 1'b1;  addr_rom[ 3137]='h00003104;  wr_data_rom[ 3137]='h00003065;
    rd_cycle[ 3138] = 1'b0;  wr_cycle[ 3138] = 1'b1;  addr_rom[ 3138]='h00003108;  wr_data_rom[ 3138]='h00001589;
    rd_cycle[ 3139] = 1'b0;  wr_cycle[ 3139] = 1'b1;  addr_rom[ 3139]='h0000310c;  wr_data_rom[ 3139]='h00001fa5;
    rd_cycle[ 3140] = 1'b0;  wr_cycle[ 3140] = 1'b1;  addr_rom[ 3140]='h00003110;  wr_data_rom[ 3140]='h00003e23;
    rd_cycle[ 3141] = 1'b0;  wr_cycle[ 3141] = 1'b1;  addr_rom[ 3141]='h00003114;  wr_data_rom[ 3141]='h00000acf;
    rd_cycle[ 3142] = 1'b0;  wr_cycle[ 3142] = 1'b1;  addr_rom[ 3142]='h00003118;  wr_data_rom[ 3142]='h000025a2;
    rd_cycle[ 3143] = 1'b0;  wr_cycle[ 3143] = 1'b1;  addr_rom[ 3143]='h0000311c;  wr_data_rom[ 3143]='h00003d4c;
    rd_cycle[ 3144] = 1'b0;  wr_cycle[ 3144] = 1'b1;  addr_rom[ 3144]='h00003120;  wr_data_rom[ 3144]='h000001cc;
    rd_cycle[ 3145] = 1'b0;  wr_cycle[ 3145] = 1'b1;  addr_rom[ 3145]='h00003124;  wr_data_rom[ 3145]='h00001ad7;
    rd_cycle[ 3146] = 1'b0;  wr_cycle[ 3146] = 1'b1;  addr_rom[ 3146]='h00003128;  wr_data_rom[ 3146]='h00000c17;
    rd_cycle[ 3147] = 1'b0;  wr_cycle[ 3147] = 1'b1;  addr_rom[ 3147]='h0000312c;  wr_data_rom[ 3147]='h000037b1;
    rd_cycle[ 3148] = 1'b0;  wr_cycle[ 3148] = 1'b1;  addr_rom[ 3148]='h00003130;  wr_data_rom[ 3148]='h00000b69;
    rd_cycle[ 3149] = 1'b0;  wr_cycle[ 3149] = 1'b1;  addr_rom[ 3149]='h00003134;  wr_data_rom[ 3149]='h00002567;
    rd_cycle[ 3150] = 1'b0;  wr_cycle[ 3150] = 1'b1;  addr_rom[ 3150]='h00003138;  wr_data_rom[ 3150]='h00000fd7;
    rd_cycle[ 3151] = 1'b0;  wr_cycle[ 3151] = 1'b1;  addr_rom[ 3151]='h0000313c;  wr_data_rom[ 3151]='h00003711;
    rd_cycle[ 3152] = 1'b0;  wr_cycle[ 3152] = 1'b1;  addr_rom[ 3152]='h00003140;  wr_data_rom[ 3152]='h000025d5;
    rd_cycle[ 3153] = 1'b0;  wr_cycle[ 3153] = 1'b1;  addr_rom[ 3153]='h00003144;  wr_data_rom[ 3153]='h000024bf;
    rd_cycle[ 3154] = 1'b0;  wr_cycle[ 3154] = 1'b1;  addr_rom[ 3154]='h00003148;  wr_data_rom[ 3154]='h000038df;
    rd_cycle[ 3155] = 1'b0;  wr_cycle[ 3155] = 1'b1;  addr_rom[ 3155]='h0000314c;  wr_data_rom[ 3155]='h000017c3;
    rd_cycle[ 3156] = 1'b0;  wr_cycle[ 3156] = 1'b1;  addr_rom[ 3156]='h00003150;  wr_data_rom[ 3156]='h00003424;
    rd_cycle[ 3157] = 1'b0;  wr_cycle[ 3157] = 1'b1;  addr_rom[ 3157]='h00003154;  wr_data_rom[ 3157]='h00002306;
    rd_cycle[ 3158] = 1'b0;  wr_cycle[ 3158] = 1'b1;  addr_rom[ 3158]='h00003158;  wr_data_rom[ 3158]='h00001b14;
    rd_cycle[ 3159] = 1'b0;  wr_cycle[ 3159] = 1'b1;  addr_rom[ 3159]='h0000315c;  wr_data_rom[ 3159]='h000000fe;
    rd_cycle[ 3160] = 1'b0;  wr_cycle[ 3160] = 1'b1;  addr_rom[ 3160]='h00003160;  wr_data_rom[ 3160]='h0000344b;
    rd_cycle[ 3161] = 1'b0;  wr_cycle[ 3161] = 1'b1;  addr_rom[ 3161]='h00003164;  wr_data_rom[ 3161]='h000004bf;
    rd_cycle[ 3162] = 1'b0;  wr_cycle[ 3162] = 1'b1;  addr_rom[ 3162]='h00003168;  wr_data_rom[ 3162]='h00003fc3;
    rd_cycle[ 3163] = 1'b0;  wr_cycle[ 3163] = 1'b1;  addr_rom[ 3163]='h0000316c;  wr_data_rom[ 3163]='h00001fd6;
    rd_cycle[ 3164] = 1'b0;  wr_cycle[ 3164] = 1'b1;  addr_rom[ 3164]='h00003170;  wr_data_rom[ 3164]='h00003ee7;
    rd_cycle[ 3165] = 1'b0;  wr_cycle[ 3165] = 1'b1;  addr_rom[ 3165]='h00003174;  wr_data_rom[ 3165]='h00001a3d;
    rd_cycle[ 3166] = 1'b0;  wr_cycle[ 3166] = 1'b1;  addr_rom[ 3166]='h00003178;  wr_data_rom[ 3166]='h000002d1;
    rd_cycle[ 3167] = 1'b0;  wr_cycle[ 3167] = 1'b1;  addr_rom[ 3167]='h0000317c;  wr_data_rom[ 3167]='h00001313;
    rd_cycle[ 3168] = 1'b0;  wr_cycle[ 3168] = 1'b1;  addr_rom[ 3168]='h00003180;  wr_data_rom[ 3168]='h000016bb;
    rd_cycle[ 3169] = 1'b0;  wr_cycle[ 3169] = 1'b1;  addr_rom[ 3169]='h00003184;  wr_data_rom[ 3169]='h00001bba;
    rd_cycle[ 3170] = 1'b0;  wr_cycle[ 3170] = 1'b1;  addr_rom[ 3170]='h00003188;  wr_data_rom[ 3170]='h00003de7;
    rd_cycle[ 3171] = 1'b0;  wr_cycle[ 3171] = 1'b1;  addr_rom[ 3171]='h0000318c;  wr_data_rom[ 3171]='h00003869;
    rd_cycle[ 3172] = 1'b0;  wr_cycle[ 3172] = 1'b1;  addr_rom[ 3172]='h00003190;  wr_data_rom[ 3172]='h00002147;
    rd_cycle[ 3173] = 1'b0;  wr_cycle[ 3173] = 1'b1;  addr_rom[ 3173]='h00003194;  wr_data_rom[ 3173]='h00003973;
    rd_cycle[ 3174] = 1'b0;  wr_cycle[ 3174] = 1'b1;  addr_rom[ 3174]='h00003198;  wr_data_rom[ 3174]='h00003f64;
    rd_cycle[ 3175] = 1'b0;  wr_cycle[ 3175] = 1'b1;  addr_rom[ 3175]='h0000319c;  wr_data_rom[ 3175]='h00002550;
    rd_cycle[ 3176] = 1'b0;  wr_cycle[ 3176] = 1'b1;  addr_rom[ 3176]='h000031a0;  wr_data_rom[ 3176]='h00001634;
    rd_cycle[ 3177] = 1'b0;  wr_cycle[ 3177] = 1'b1;  addr_rom[ 3177]='h000031a4;  wr_data_rom[ 3177]='h0000035f;
    rd_cycle[ 3178] = 1'b0;  wr_cycle[ 3178] = 1'b1;  addr_rom[ 3178]='h000031a8;  wr_data_rom[ 3178]='h00003256;
    rd_cycle[ 3179] = 1'b0;  wr_cycle[ 3179] = 1'b1;  addr_rom[ 3179]='h000031ac;  wr_data_rom[ 3179]='h000013e3;
    rd_cycle[ 3180] = 1'b0;  wr_cycle[ 3180] = 1'b1;  addr_rom[ 3180]='h000031b0;  wr_data_rom[ 3180]='h00003ed4;
    rd_cycle[ 3181] = 1'b0;  wr_cycle[ 3181] = 1'b1;  addr_rom[ 3181]='h000031b4;  wr_data_rom[ 3181]='h000016b8;
    rd_cycle[ 3182] = 1'b0;  wr_cycle[ 3182] = 1'b1;  addr_rom[ 3182]='h000031b8;  wr_data_rom[ 3182]='h0000040a;
    rd_cycle[ 3183] = 1'b0;  wr_cycle[ 3183] = 1'b1;  addr_rom[ 3183]='h000031bc;  wr_data_rom[ 3183]='h000039c9;
    rd_cycle[ 3184] = 1'b0;  wr_cycle[ 3184] = 1'b1;  addr_rom[ 3184]='h000031c0;  wr_data_rom[ 3184]='h00001898;
    rd_cycle[ 3185] = 1'b0;  wr_cycle[ 3185] = 1'b1;  addr_rom[ 3185]='h000031c4;  wr_data_rom[ 3185]='h00003151;
    rd_cycle[ 3186] = 1'b0;  wr_cycle[ 3186] = 1'b1;  addr_rom[ 3186]='h000031c8;  wr_data_rom[ 3186]='h00003516;
    rd_cycle[ 3187] = 1'b0;  wr_cycle[ 3187] = 1'b1;  addr_rom[ 3187]='h000031cc;  wr_data_rom[ 3187]='h0000015d;
    rd_cycle[ 3188] = 1'b0;  wr_cycle[ 3188] = 1'b1;  addr_rom[ 3188]='h000031d0;  wr_data_rom[ 3188]='h00001aef;
    rd_cycle[ 3189] = 1'b0;  wr_cycle[ 3189] = 1'b1;  addr_rom[ 3189]='h000031d4;  wr_data_rom[ 3189]='h00003e35;
    rd_cycle[ 3190] = 1'b0;  wr_cycle[ 3190] = 1'b1;  addr_rom[ 3190]='h000031d8;  wr_data_rom[ 3190]='h000011cd;
    rd_cycle[ 3191] = 1'b0;  wr_cycle[ 3191] = 1'b1;  addr_rom[ 3191]='h000031dc;  wr_data_rom[ 3191]='h00003883;
    rd_cycle[ 3192] = 1'b0;  wr_cycle[ 3192] = 1'b1;  addr_rom[ 3192]='h000031e0;  wr_data_rom[ 3192]='h000012a7;
    rd_cycle[ 3193] = 1'b0;  wr_cycle[ 3193] = 1'b1;  addr_rom[ 3193]='h000031e4;  wr_data_rom[ 3193]='h000017e0;
    rd_cycle[ 3194] = 1'b0;  wr_cycle[ 3194] = 1'b1;  addr_rom[ 3194]='h000031e8;  wr_data_rom[ 3194]='h00002ad2;
    rd_cycle[ 3195] = 1'b0;  wr_cycle[ 3195] = 1'b1;  addr_rom[ 3195]='h000031ec;  wr_data_rom[ 3195]='h00001cd2;
    rd_cycle[ 3196] = 1'b0;  wr_cycle[ 3196] = 1'b1;  addr_rom[ 3196]='h000031f0;  wr_data_rom[ 3196]='h00003112;
    rd_cycle[ 3197] = 1'b0;  wr_cycle[ 3197] = 1'b1;  addr_rom[ 3197]='h000031f4;  wr_data_rom[ 3197]='h000002bb;
    rd_cycle[ 3198] = 1'b0;  wr_cycle[ 3198] = 1'b1;  addr_rom[ 3198]='h000031f8;  wr_data_rom[ 3198]='h00003436;
    rd_cycle[ 3199] = 1'b0;  wr_cycle[ 3199] = 1'b1;  addr_rom[ 3199]='h000031fc;  wr_data_rom[ 3199]='h0000207d;
    rd_cycle[ 3200] = 1'b0;  wr_cycle[ 3200] = 1'b1;  addr_rom[ 3200]='h00003200;  wr_data_rom[ 3200]='h000038eb;
    rd_cycle[ 3201] = 1'b0;  wr_cycle[ 3201] = 1'b1;  addr_rom[ 3201]='h00003204;  wr_data_rom[ 3201]='h00001c7f;
    rd_cycle[ 3202] = 1'b0;  wr_cycle[ 3202] = 1'b1;  addr_rom[ 3202]='h00003208;  wr_data_rom[ 3202]='h00003753;
    rd_cycle[ 3203] = 1'b0;  wr_cycle[ 3203] = 1'b1;  addr_rom[ 3203]='h0000320c;  wr_data_rom[ 3203]='h00000983;
    rd_cycle[ 3204] = 1'b0;  wr_cycle[ 3204] = 1'b1;  addr_rom[ 3204]='h00003210;  wr_data_rom[ 3204]='h00001a87;
    rd_cycle[ 3205] = 1'b0;  wr_cycle[ 3205] = 1'b1;  addr_rom[ 3205]='h00003214;  wr_data_rom[ 3205]='h0000312f;
    rd_cycle[ 3206] = 1'b0;  wr_cycle[ 3206] = 1'b1;  addr_rom[ 3206]='h00003218;  wr_data_rom[ 3206]='h000033e1;
    rd_cycle[ 3207] = 1'b0;  wr_cycle[ 3207] = 1'b1;  addr_rom[ 3207]='h0000321c;  wr_data_rom[ 3207]='h0000006f;
    rd_cycle[ 3208] = 1'b0;  wr_cycle[ 3208] = 1'b1;  addr_rom[ 3208]='h00003220;  wr_data_rom[ 3208]='h00000d6a;
    rd_cycle[ 3209] = 1'b0;  wr_cycle[ 3209] = 1'b1;  addr_rom[ 3209]='h00003224;  wr_data_rom[ 3209]='h000006a5;
    rd_cycle[ 3210] = 1'b0;  wr_cycle[ 3210] = 1'b1;  addr_rom[ 3210]='h00003228;  wr_data_rom[ 3210]='h00000483;
    rd_cycle[ 3211] = 1'b0;  wr_cycle[ 3211] = 1'b1;  addr_rom[ 3211]='h0000322c;  wr_data_rom[ 3211]='h00001b11;
    rd_cycle[ 3212] = 1'b0;  wr_cycle[ 3212] = 1'b1;  addr_rom[ 3212]='h00003230;  wr_data_rom[ 3212]='h000016e8;
    rd_cycle[ 3213] = 1'b0;  wr_cycle[ 3213] = 1'b1;  addr_rom[ 3213]='h00003234;  wr_data_rom[ 3213]='h00003c1e;
    rd_cycle[ 3214] = 1'b0;  wr_cycle[ 3214] = 1'b1;  addr_rom[ 3214]='h00003238;  wr_data_rom[ 3214]='h000019e0;
    rd_cycle[ 3215] = 1'b0;  wr_cycle[ 3215] = 1'b1;  addr_rom[ 3215]='h0000323c;  wr_data_rom[ 3215]='h00000203;
    rd_cycle[ 3216] = 1'b0;  wr_cycle[ 3216] = 1'b1;  addr_rom[ 3216]='h00003240;  wr_data_rom[ 3216]='h00003a03;
    rd_cycle[ 3217] = 1'b0;  wr_cycle[ 3217] = 1'b1;  addr_rom[ 3217]='h00003244;  wr_data_rom[ 3217]='h0000004c;
    rd_cycle[ 3218] = 1'b0;  wr_cycle[ 3218] = 1'b1;  addr_rom[ 3218]='h00003248;  wr_data_rom[ 3218]='h00000cba;
    rd_cycle[ 3219] = 1'b0;  wr_cycle[ 3219] = 1'b1;  addr_rom[ 3219]='h0000324c;  wr_data_rom[ 3219]='h00001e0c;
    rd_cycle[ 3220] = 1'b0;  wr_cycle[ 3220] = 1'b1;  addr_rom[ 3220]='h00003250;  wr_data_rom[ 3220]='h0000051b;
    rd_cycle[ 3221] = 1'b0;  wr_cycle[ 3221] = 1'b1;  addr_rom[ 3221]='h00003254;  wr_data_rom[ 3221]='h00003db8;
    rd_cycle[ 3222] = 1'b0;  wr_cycle[ 3222] = 1'b1;  addr_rom[ 3222]='h00003258;  wr_data_rom[ 3222]='h000003d6;
    rd_cycle[ 3223] = 1'b0;  wr_cycle[ 3223] = 1'b1;  addr_rom[ 3223]='h0000325c;  wr_data_rom[ 3223]='h0000068e;
    rd_cycle[ 3224] = 1'b0;  wr_cycle[ 3224] = 1'b1;  addr_rom[ 3224]='h00003260;  wr_data_rom[ 3224]='h00002818;
    rd_cycle[ 3225] = 1'b0;  wr_cycle[ 3225] = 1'b1;  addr_rom[ 3225]='h00003264;  wr_data_rom[ 3225]='h00003031;
    rd_cycle[ 3226] = 1'b0;  wr_cycle[ 3226] = 1'b1;  addr_rom[ 3226]='h00003268;  wr_data_rom[ 3226]='h000017f5;
    rd_cycle[ 3227] = 1'b0;  wr_cycle[ 3227] = 1'b1;  addr_rom[ 3227]='h0000326c;  wr_data_rom[ 3227]='h00001d15;
    rd_cycle[ 3228] = 1'b0;  wr_cycle[ 3228] = 1'b1;  addr_rom[ 3228]='h00003270;  wr_data_rom[ 3228]='h00003c8f;
    rd_cycle[ 3229] = 1'b0;  wr_cycle[ 3229] = 1'b1;  addr_rom[ 3229]='h00003274;  wr_data_rom[ 3229]='h000020b9;
    rd_cycle[ 3230] = 1'b0;  wr_cycle[ 3230] = 1'b1;  addr_rom[ 3230]='h00003278;  wr_data_rom[ 3230]='h0000103b;
    rd_cycle[ 3231] = 1'b0;  wr_cycle[ 3231] = 1'b1;  addr_rom[ 3231]='h0000327c;  wr_data_rom[ 3231]='h00003d4e;
    rd_cycle[ 3232] = 1'b0;  wr_cycle[ 3232] = 1'b1;  addr_rom[ 3232]='h00003280;  wr_data_rom[ 3232]='h00000889;
    rd_cycle[ 3233] = 1'b0;  wr_cycle[ 3233] = 1'b1;  addr_rom[ 3233]='h00003284;  wr_data_rom[ 3233]='h0000280f;
    rd_cycle[ 3234] = 1'b0;  wr_cycle[ 3234] = 1'b1;  addr_rom[ 3234]='h00003288;  wr_data_rom[ 3234]='h00000321;
    rd_cycle[ 3235] = 1'b0;  wr_cycle[ 3235] = 1'b1;  addr_rom[ 3235]='h0000328c;  wr_data_rom[ 3235]='h00002f98;
    rd_cycle[ 3236] = 1'b0;  wr_cycle[ 3236] = 1'b1;  addr_rom[ 3236]='h00003290;  wr_data_rom[ 3236]='h0000191e;
    rd_cycle[ 3237] = 1'b0;  wr_cycle[ 3237] = 1'b1;  addr_rom[ 3237]='h00003294;  wr_data_rom[ 3237]='h00003596;
    rd_cycle[ 3238] = 1'b0;  wr_cycle[ 3238] = 1'b1;  addr_rom[ 3238]='h00003298;  wr_data_rom[ 3238]='h00003579;
    rd_cycle[ 3239] = 1'b0;  wr_cycle[ 3239] = 1'b1;  addr_rom[ 3239]='h0000329c;  wr_data_rom[ 3239]='h000005e8;
    rd_cycle[ 3240] = 1'b0;  wr_cycle[ 3240] = 1'b1;  addr_rom[ 3240]='h000032a0;  wr_data_rom[ 3240]='h000012d8;
    rd_cycle[ 3241] = 1'b0;  wr_cycle[ 3241] = 1'b1;  addr_rom[ 3241]='h000032a4;  wr_data_rom[ 3241]='h000038c9;
    rd_cycle[ 3242] = 1'b0;  wr_cycle[ 3242] = 1'b1;  addr_rom[ 3242]='h000032a8;  wr_data_rom[ 3242]='h00002859;
    rd_cycle[ 3243] = 1'b0;  wr_cycle[ 3243] = 1'b1;  addr_rom[ 3243]='h000032ac;  wr_data_rom[ 3243]='h00001601;
    rd_cycle[ 3244] = 1'b0;  wr_cycle[ 3244] = 1'b1;  addr_rom[ 3244]='h000032b0;  wr_data_rom[ 3244]='h00000716;
    rd_cycle[ 3245] = 1'b0;  wr_cycle[ 3245] = 1'b1;  addr_rom[ 3245]='h000032b4;  wr_data_rom[ 3245]='h00002b92;
    rd_cycle[ 3246] = 1'b0;  wr_cycle[ 3246] = 1'b1;  addr_rom[ 3246]='h000032b8;  wr_data_rom[ 3246]='h000013d0;
    rd_cycle[ 3247] = 1'b0;  wr_cycle[ 3247] = 1'b1;  addr_rom[ 3247]='h000032bc;  wr_data_rom[ 3247]='h00000202;
    rd_cycle[ 3248] = 1'b0;  wr_cycle[ 3248] = 1'b1;  addr_rom[ 3248]='h000032c0;  wr_data_rom[ 3248]='h00002f9f;
    rd_cycle[ 3249] = 1'b0;  wr_cycle[ 3249] = 1'b1;  addr_rom[ 3249]='h000032c4;  wr_data_rom[ 3249]='h000000bb;
    rd_cycle[ 3250] = 1'b0;  wr_cycle[ 3250] = 1'b1;  addr_rom[ 3250]='h000032c8;  wr_data_rom[ 3250]='h00001ebe;
    rd_cycle[ 3251] = 1'b0;  wr_cycle[ 3251] = 1'b1;  addr_rom[ 3251]='h000032cc;  wr_data_rom[ 3251]='h00001148;
    rd_cycle[ 3252] = 1'b0;  wr_cycle[ 3252] = 1'b1;  addr_rom[ 3252]='h000032d0;  wr_data_rom[ 3252]='h000026a8;
    rd_cycle[ 3253] = 1'b0;  wr_cycle[ 3253] = 1'b1;  addr_rom[ 3253]='h000032d4;  wr_data_rom[ 3253]='h0000024b;
    rd_cycle[ 3254] = 1'b0;  wr_cycle[ 3254] = 1'b1;  addr_rom[ 3254]='h000032d8;  wr_data_rom[ 3254]='h00001509;
    rd_cycle[ 3255] = 1'b0;  wr_cycle[ 3255] = 1'b1;  addr_rom[ 3255]='h000032dc;  wr_data_rom[ 3255]='h000019a3;
    rd_cycle[ 3256] = 1'b0;  wr_cycle[ 3256] = 1'b1;  addr_rom[ 3256]='h000032e0;  wr_data_rom[ 3256]='h0000063b;
    rd_cycle[ 3257] = 1'b0;  wr_cycle[ 3257] = 1'b1;  addr_rom[ 3257]='h000032e4;  wr_data_rom[ 3257]='h00000ed2;
    rd_cycle[ 3258] = 1'b0;  wr_cycle[ 3258] = 1'b1;  addr_rom[ 3258]='h000032e8;  wr_data_rom[ 3258]='h000026e4;
    rd_cycle[ 3259] = 1'b0;  wr_cycle[ 3259] = 1'b1;  addr_rom[ 3259]='h000032ec;  wr_data_rom[ 3259]='h0000328c;
    rd_cycle[ 3260] = 1'b0;  wr_cycle[ 3260] = 1'b1;  addr_rom[ 3260]='h000032f0;  wr_data_rom[ 3260]='h00001f25;
    rd_cycle[ 3261] = 1'b0;  wr_cycle[ 3261] = 1'b1;  addr_rom[ 3261]='h000032f4;  wr_data_rom[ 3261]='h0000288d;
    rd_cycle[ 3262] = 1'b0;  wr_cycle[ 3262] = 1'b1;  addr_rom[ 3262]='h000032f8;  wr_data_rom[ 3262]='h000035f5;
    rd_cycle[ 3263] = 1'b0;  wr_cycle[ 3263] = 1'b1;  addr_rom[ 3263]='h000032fc;  wr_data_rom[ 3263]='h000001e3;
    rd_cycle[ 3264] = 1'b0;  wr_cycle[ 3264] = 1'b1;  addr_rom[ 3264]='h00003300;  wr_data_rom[ 3264]='h000014c2;
    rd_cycle[ 3265] = 1'b0;  wr_cycle[ 3265] = 1'b1;  addr_rom[ 3265]='h00003304;  wr_data_rom[ 3265]='h000020d4;
    rd_cycle[ 3266] = 1'b0;  wr_cycle[ 3266] = 1'b1;  addr_rom[ 3266]='h00003308;  wr_data_rom[ 3266]='h00000c63;
    rd_cycle[ 3267] = 1'b0;  wr_cycle[ 3267] = 1'b1;  addr_rom[ 3267]='h0000330c;  wr_data_rom[ 3267]='h000019d0;
    rd_cycle[ 3268] = 1'b0;  wr_cycle[ 3268] = 1'b1;  addr_rom[ 3268]='h00003310;  wr_data_rom[ 3268]='h00000413;
    rd_cycle[ 3269] = 1'b0;  wr_cycle[ 3269] = 1'b1;  addr_rom[ 3269]='h00003314;  wr_data_rom[ 3269]='h0000352e;
    rd_cycle[ 3270] = 1'b0;  wr_cycle[ 3270] = 1'b1;  addr_rom[ 3270]='h00003318;  wr_data_rom[ 3270]='h000003c4;
    rd_cycle[ 3271] = 1'b0;  wr_cycle[ 3271] = 1'b1;  addr_rom[ 3271]='h0000331c;  wr_data_rom[ 3271]='h00000cf9;
    rd_cycle[ 3272] = 1'b0;  wr_cycle[ 3272] = 1'b1;  addr_rom[ 3272]='h00003320;  wr_data_rom[ 3272]='h000001b1;
    rd_cycle[ 3273] = 1'b0;  wr_cycle[ 3273] = 1'b1;  addr_rom[ 3273]='h00003324;  wr_data_rom[ 3273]='h00003725;
    rd_cycle[ 3274] = 1'b0;  wr_cycle[ 3274] = 1'b1;  addr_rom[ 3274]='h00003328;  wr_data_rom[ 3274]='h00001fa9;
    rd_cycle[ 3275] = 1'b0;  wr_cycle[ 3275] = 1'b1;  addr_rom[ 3275]='h0000332c;  wr_data_rom[ 3275]='h00001e43;
    rd_cycle[ 3276] = 1'b0;  wr_cycle[ 3276] = 1'b1;  addr_rom[ 3276]='h00003330;  wr_data_rom[ 3276]='h00002715;
    rd_cycle[ 3277] = 1'b0;  wr_cycle[ 3277] = 1'b1;  addr_rom[ 3277]='h00003334;  wr_data_rom[ 3277]='h000020a8;
    rd_cycle[ 3278] = 1'b0;  wr_cycle[ 3278] = 1'b1;  addr_rom[ 3278]='h00003338;  wr_data_rom[ 3278]='h0000000e;
    rd_cycle[ 3279] = 1'b0;  wr_cycle[ 3279] = 1'b1;  addr_rom[ 3279]='h0000333c;  wr_data_rom[ 3279]='h00003c01;
    rd_cycle[ 3280] = 1'b0;  wr_cycle[ 3280] = 1'b1;  addr_rom[ 3280]='h00003340;  wr_data_rom[ 3280]='h0000269f;
    rd_cycle[ 3281] = 1'b0;  wr_cycle[ 3281] = 1'b1;  addr_rom[ 3281]='h00003344;  wr_data_rom[ 3281]='h000013ee;
    rd_cycle[ 3282] = 1'b0;  wr_cycle[ 3282] = 1'b1;  addr_rom[ 3282]='h00003348;  wr_data_rom[ 3282]='h00001108;
    rd_cycle[ 3283] = 1'b0;  wr_cycle[ 3283] = 1'b1;  addr_rom[ 3283]='h0000334c;  wr_data_rom[ 3283]='h000033f7;
    rd_cycle[ 3284] = 1'b0;  wr_cycle[ 3284] = 1'b1;  addr_rom[ 3284]='h00003350;  wr_data_rom[ 3284]='h00003ae6;
    rd_cycle[ 3285] = 1'b0;  wr_cycle[ 3285] = 1'b1;  addr_rom[ 3285]='h00003354;  wr_data_rom[ 3285]='h0000040f;
    rd_cycle[ 3286] = 1'b0;  wr_cycle[ 3286] = 1'b1;  addr_rom[ 3286]='h00003358;  wr_data_rom[ 3286]='h00001ed9;
    rd_cycle[ 3287] = 1'b0;  wr_cycle[ 3287] = 1'b1;  addr_rom[ 3287]='h0000335c;  wr_data_rom[ 3287]='h00003346;
    rd_cycle[ 3288] = 1'b0;  wr_cycle[ 3288] = 1'b1;  addr_rom[ 3288]='h00003360;  wr_data_rom[ 3288]='h000005e3;
    rd_cycle[ 3289] = 1'b0;  wr_cycle[ 3289] = 1'b1;  addr_rom[ 3289]='h00003364;  wr_data_rom[ 3289]='h0000389a;
    rd_cycle[ 3290] = 1'b0;  wr_cycle[ 3290] = 1'b1;  addr_rom[ 3290]='h00003368;  wr_data_rom[ 3290]='h00002817;
    rd_cycle[ 3291] = 1'b0;  wr_cycle[ 3291] = 1'b1;  addr_rom[ 3291]='h0000336c;  wr_data_rom[ 3291]='h000004ce;
    rd_cycle[ 3292] = 1'b0;  wr_cycle[ 3292] = 1'b1;  addr_rom[ 3292]='h00003370;  wr_data_rom[ 3292]='h0000106f;
    rd_cycle[ 3293] = 1'b0;  wr_cycle[ 3293] = 1'b1;  addr_rom[ 3293]='h00003374;  wr_data_rom[ 3293]='h00001aad;
    rd_cycle[ 3294] = 1'b0;  wr_cycle[ 3294] = 1'b1;  addr_rom[ 3294]='h00003378;  wr_data_rom[ 3294]='h00000273;
    rd_cycle[ 3295] = 1'b0;  wr_cycle[ 3295] = 1'b1;  addr_rom[ 3295]='h0000337c;  wr_data_rom[ 3295]='h00000a9c;
    rd_cycle[ 3296] = 1'b0;  wr_cycle[ 3296] = 1'b1;  addr_rom[ 3296]='h00003380;  wr_data_rom[ 3296]='h00003b85;
    rd_cycle[ 3297] = 1'b0;  wr_cycle[ 3297] = 1'b1;  addr_rom[ 3297]='h00003384;  wr_data_rom[ 3297]='h000032a0;
    rd_cycle[ 3298] = 1'b0;  wr_cycle[ 3298] = 1'b1;  addr_rom[ 3298]='h00003388;  wr_data_rom[ 3298]='h00000788;
    rd_cycle[ 3299] = 1'b0;  wr_cycle[ 3299] = 1'b1;  addr_rom[ 3299]='h0000338c;  wr_data_rom[ 3299]='h00003972;
    rd_cycle[ 3300] = 1'b0;  wr_cycle[ 3300] = 1'b1;  addr_rom[ 3300]='h00003390;  wr_data_rom[ 3300]='h000001f8;
    rd_cycle[ 3301] = 1'b0;  wr_cycle[ 3301] = 1'b1;  addr_rom[ 3301]='h00003394;  wr_data_rom[ 3301]='h0000148c;
    rd_cycle[ 3302] = 1'b0;  wr_cycle[ 3302] = 1'b1;  addr_rom[ 3302]='h00003398;  wr_data_rom[ 3302]='h0000336d;
    rd_cycle[ 3303] = 1'b0;  wr_cycle[ 3303] = 1'b1;  addr_rom[ 3303]='h0000339c;  wr_data_rom[ 3303]='h0000227c;
    rd_cycle[ 3304] = 1'b0;  wr_cycle[ 3304] = 1'b1;  addr_rom[ 3304]='h000033a0;  wr_data_rom[ 3304]='h00001d32;
    rd_cycle[ 3305] = 1'b0;  wr_cycle[ 3305] = 1'b1;  addr_rom[ 3305]='h000033a4;  wr_data_rom[ 3305]='h0000210b;
    rd_cycle[ 3306] = 1'b0;  wr_cycle[ 3306] = 1'b1;  addr_rom[ 3306]='h000033a8;  wr_data_rom[ 3306]='h000023c2;
    rd_cycle[ 3307] = 1'b0;  wr_cycle[ 3307] = 1'b1;  addr_rom[ 3307]='h000033ac;  wr_data_rom[ 3307]='h00002029;
    rd_cycle[ 3308] = 1'b0;  wr_cycle[ 3308] = 1'b1;  addr_rom[ 3308]='h000033b0;  wr_data_rom[ 3308]='h000035b9;
    rd_cycle[ 3309] = 1'b0;  wr_cycle[ 3309] = 1'b1;  addr_rom[ 3309]='h000033b4;  wr_data_rom[ 3309]='h00002bee;
    rd_cycle[ 3310] = 1'b0;  wr_cycle[ 3310] = 1'b1;  addr_rom[ 3310]='h000033b8;  wr_data_rom[ 3310]='h00000ea4;
    rd_cycle[ 3311] = 1'b0;  wr_cycle[ 3311] = 1'b1;  addr_rom[ 3311]='h000033bc;  wr_data_rom[ 3311]='h0000272d;
    rd_cycle[ 3312] = 1'b0;  wr_cycle[ 3312] = 1'b1;  addr_rom[ 3312]='h000033c0;  wr_data_rom[ 3312]='h00001823;
    rd_cycle[ 3313] = 1'b0;  wr_cycle[ 3313] = 1'b1;  addr_rom[ 3313]='h000033c4;  wr_data_rom[ 3313]='h000000ec;
    rd_cycle[ 3314] = 1'b0;  wr_cycle[ 3314] = 1'b1;  addr_rom[ 3314]='h000033c8;  wr_data_rom[ 3314]='h0000048c;
    rd_cycle[ 3315] = 1'b0;  wr_cycle[ 3315] = 1'b1;  addr_rom[ 3315]='h000033cc;  wr_data_rom[ 3315]='h0000267c;
    rd_cycle[ 3316] = 1'b0;  wr_cycle[ 3316] = 1'b1;  addr_rom[ 3316]='h000033d0;  wr_data_rom[ 3316]='h00001c86;
    rd_cycle[ 3317] = 1'b0;  wr_cycle[ 3317] = 1'b1;  addr_rom[ 3317]='h000033d4;  wr_data_rom[ 3317]='h00001438;
    rd_cycle[ 3318] = 1'b0;  wr_cycle[ 3318] = 1'b1;  addr_rom[ 3318]='h000033d8;  wr_data_rom[ 3318]='h00000fb7;
    rd_cycle[ 3319] = 1'b0;  wr_cycle[ 3319] = 1'b1;  addr_rom[ 3319]='h000033dc;  wr_data_rom[ 3319]='h00003fd1;
    rd_cycle[ 3320] = 1'b0;  wr_cycle[ 3320] = 1'b1;  addr_rom[ 3320]='h000033e0;  wr_data_rom[ 3320]='h00000f6e;
    rd_cycle[ 3321] = 1'b0;  wr_cycle[ 3321] = 1'b1;  addr_rom[ 3321]='h000033e4;  wr_data_rom[ 3321]='h0000348f;
    rd_cycle[ 3322] = 1'b0;  wr_cycle[ 3322] = 1'b1;  addr_rom[ 3322]='h000033e8;  wr_data_rom[ 3322]='h00003ea5;
    rd_cycle[ 3323] = 1'b0;  wr_cycle[ 3323] = 1'b1;  addr_rom[ 3323]='h000033ec;  wr_data_rom[ 3323]='h00002834;
    rd_cycle[ 3324] = 1'b0;  wr_cycle[ 3324] = 1'b1;  addr_rom[ 3324]='h000033f0;  wr_data_rom[ 3324]='h00001836;
    rd_cycle[ 3325] = 1'b0;  wr_cycle[ 3325] = 1'b1;  addr_rom[ 3325]='h000033f4;  wr_data_rom[ 3325]='h00000620;
    rd_cycle[ 3326] = 1'b0;  wr_cycle[ 3326] = 1'b1;  addr_rom[ 3326]='h000033f8;  wr_data_rom[ 3326]='h0000024e;
    rd_cycle[ 3327] = 1'b0;  wr_cycle[ 3327] = 1'b1;  addr_rom[ 3327]='h000033fc;  wr_data_rom[ 3327]='h00001ddb;
    rd_cycle[ 3328] = 1'b0;  wr_cycle[ 3328] = 1'b1;  addr_rom[ 3328]='h00003400;  wr_data_rom[ 3328]='h00003924;
    rd_cycle[ 3329] = 1'b0;  wr_cycle[ 3329] = 1'b1;  addr_rom[ 3329]='h00003404;  wr_data_rom[ 3329]='h0000359c;
    rd_cycle[ 3330] = 1'b0;  wr_cycle[ 3330] = 1'b1;  addr_rom[ 3330]='h00003408;  wr_data_rom[ 3330]='h0000249e;
    rd_cycle[ 3331] = 1'b0;  wr_cycle[ 3331] = 1'b1;  addr_rom[ 3331]='h0000340c;  wr_data_rom[ 3331]='h00002318;
    rd_cycle[ 3332] = 1'b0;  wr_cycle[ 3332] = 1'b1;  addr_rom[ 3332]='h00003410;  wr_data_rom[ 3332]='h00002cba;
    rd_cycle[ 3333] = 1'b0;  wr_cycle[ 3333] = 1'b1;  addr_rom[ 3333]='h00003414;  wr_data_rom[ 3333]='h0000048c;
    rd_cycle[ 3334] = 1'b0;  wr_cycle[ 3334] = 1'b1;  addr_rom[ 3334]='h00003418;  wr_data_rom[ 3334]='h00002bbc;
    rd_cycle[ 3335] = 1'b0;  wr_cycle[ 3335] = 1'b1;  addr_rom[ 3335]='h0000341c;  wr_data_rom[ 3335]='h0000347e;
    rd_cycle[ 3336] = 1'b0;  wr_cycle[ 3336] = 1'b1;  addr_rom[ 3336]='h00003420;  wr_data_rom[ 3336]='h0000366d;
    rd_cycle[ 3337] = 1'b0;  wr_cycle[ 3337] = 1'b1;  addr_rom[ 3337]='h00003424;  wr_data_rom[ 3337]='h0000076d;
    rd_cycle[ 3338] = 1'b0;  wr_cycle[ 3338] = 1'b1;  addr_rom[ 3338]='h00003428;  wr_data_rom[ 3338]='h00003e9a;
    rd_cycle[ 3339] = 1'b0;  wr_cycle[ 3339] = 1'b1;  addr_rom[ 3339]='h0000342c;  wr_data_rom[ 3339]='h000009a8;
    rd_cycle[ 3340] = 1'b0;  wr_cycle[ 3340] = 1'b1;  addr_rom[ 3340]='h00003430;  wr_data_rom[ 3340]='h00001322;
    rd_cycle[ 3341] = 1'b0;  wr_cycle[ 3341] = 1'b1;  addr_rom[ 3341]='h00003434;  wr_data_rom[ 3341]='h00003421;
    rd_cycle[ 3342] = 1'b0;  wr_cycle[ 3342] = 1'b1;  addr_rom[ 3342]='h00003438;  wr_data_rom[ 3342]='h0000044c;
    rd_cycle[ 3343] = 1'b0;  wr_cycle[ 3343] = 1'b1;  addr_rom[ 3343]='h0000343c;  wr_data_rom[ 3343]='h00001e6a;
    rd_cycle[ 3344] = 1'b0;  wr_cycle[ 3344] = 1'b1;  addr_rom[ 3344]='h00003440;  wr_data_rom[ 3344]='h00000dca;
    rd_cycle[ 3345] = 1'b0;  wr_cycle[ 3345] = 1'b1;  addr_rom[ 3345]='h00003444;  wr_data_rom[ 3345]='h000027c2;
    rd_cycle[ 3346] = 1'b0;  wr_cycle[ 3346] = 1'b1;  addr_rom[ 3346]='h00003448;  wr_data_rom[ 3346]='h00002512;
    rd_cycle[ 3347] = 1'b0;  wr_cycle[ 3347] = 1'b1;  addr_rom[ 3347]='h0000344c;  wr_data_rom[ 3347]='h00002576;
    rd_cycle[ 3348] = 1'b0;  wr_cycle[ 3348] = 1'b1;  addr_rom[ 3348]='h00003450;  wr_data_rom[ 3348]='h000033d2;
    rd_cycle[ 3349] = 1'b0;  wr_cycle[ 3349] = 1'b1;  addr_rom[ 3349]='h00003454;  wr_data_rom[ 3349]='h000030b6;
    rd_cycle[ 3350] = 1'b0;  wr_cycle[ 3350] = 1'b1;  addr_rom[ 3350]='h00003458;  wr_data_rom[ 3350]='h00001b7c;
    rd_cycle[ 3351] = 1'b0;  wr_cycle[ 3351] = 1'b1;  addr_rom[ 3351]='h0000345c;  wr_data_rom[ 3351]='h000002f6;
    rd_cycle[ 3352] = 1'b0;  wr_cycle[ 3352] = 1'b1;  addr_rom[ 3352]='h00003460;  wr_data_rom[ 3352]='h00003dd5;
    rd_cycle[ 3353] = 1'b0;  wr_cycle[ 3353] = 1'b1;  addr_rom[ 3353]='h00003464;  wr_data_rom[ 3353]='h00002f33;
    rd_cycle[ 3354] = 1'b0;  wr_cycle[ 3354] = 1'b1;  addr_rom[ 3354]='h00003468;  wr_data_rom[ 3354]='h00003fb0;
    rd_cycle[ 3355] = 1'b0;  wr_cycle[ 3355] = 1'b1;  addr_rom[ 3355]='h0000346c;  wr_data_rom[ 3355]='h0000259e;
    rd_cycle[ 3356] = 1'b0;  wr_cycle[ 3356] = 1'b1;  addr_rom[ 3356]='h00003470;  wr_data_rom[ 3356]='h00000688;
    rd_cycle[ 3357] = 1'b0;  wr_cycle[ 3357] = 1'b1;  addr_rom[ 3357]='h00003474;  wr_data_rom[ 3357]='h00003285;
    rd_cycle[ 3358] = 1'b0;  wr_cycle[ 3358] = 1'b1;  addr_rom[ 3358]='h00003478;  wr_data_rom[ 3358]='h00001f15;
    rd_cycle[ 3359] = 1'b0;  wr_cycle[ 3359] = 1'b1;  addr_rom[ 3359]='h0000347c;  wr_data_rom[ 3359]='h000009c8;
    rd_cycle[ 3360] = 1'b0;  wr_cycle[ 3360] = 1'b1;  addr_rom[ 3360]='h00003480;  wr_data_rom[ 3360]='h000014eb;
    rd_cycle[ 3361] = 1'b0;  wr_cycle[ 3361] = 1'b1;  addr_rom[ 3361]='h00003484;  wr_data_rom[ 3361]='h00000aa7;
    rd_cycle[ 3362] = 1'b0;  wr_cycle[ 3362] = 1'b1;  addr_rom[ 3362]='h00003488;  wr_data_rom[ 3362]='h0000202b;
    rd_cycle[ 3363] = 1'b0;  wr_cycle[ 3363] = 1'b1;  addr_rom[ 3363]='h0000348c;  wr_data_rom[ 3363]='h00001cdb;
    rd_cycle[ 3364] = 1'b0;  wr_cycle[ 3364] = 1'b1;  addr_rom[ 3364]='h00003490;  wr_data_rom[ 3364]='h000035d4;
    rd_cycle[ 3365] = 1'b0;  wr_cycle[ 3365] = 1'b1;  addr_rom[ 3365]='h00003494;  wr_data_rom[ 3365]='h00000a60;
    rd_cycle[ 3366] = 1'b0;  wr_cycle[ 3366] = 1'b1;  addr_rom[ 3366]='h00003498;  wr_data_rom[ 3366]='h00002590;
    rd_cycle[ 3367] = 1'b0;  wr_cycle[ 3367] = 1'b1;  addr_rom[ 3367]='h0000349c;  wr_data_rom[ 3367]='h0000195b;
    rd_cycle[ 3368] = 1'b0;  wr_cycle[ 3368] = 1'b1;  addr_rom[ 3368]='h000034a0;  wr_data_rom[ 3368]='h0000021e;
    rd_cycle[ 3369] = 1'b0;  wr_cycle[ 3369] = 1'b1;  addr_rom[ 3369]='h000034a4;  wr_data_rom[ 3369]='h00002ca8;
    rd_cycle[ 3370] = 1'b0;  wr_cycle[ 3370] = 1'b1;  addr_rom[ 3370]='h000034a8;  wr_data_rom[ 3370]='h0000151d;
    rd_cycle[ 3371] = 1'b0;  wr_cycle[ 3371] = 1'b1;  addr_rom[ 3371]='h000034ac;  wr_data_rom[ 3371]='h00003c5b;
    rd_cycle[ 3372] = 1'b0;  wr_cycle[ 3372] = 1'b1;  addr_rom[ 3372]='h000034b0;  wr_data_rom[ 3372]='h00001db8;
    rd_cycle[ 3373] = 1'b0;  wr_cycle[ 3373] = 1'b1;  addr_rom[ 3373]='h000034b4;  wr_data_rom[ 3373]='h000035dd;
    rd_cycle[ 3374] = 1'b0;  wr_cycle[ 3374] = 1'b1;  addr_rom[ 3374]='h000034b8;  wr_data_rom[ 3374]='h00003d69;
    rd_cycle[ 3375] = 1'b0;  wr_cycle[ 3375] = 1'b1;  addr_rom[ 3375]='h000034bc;  wr_data_rom[ 3375]='h000035f5;
    rd_cycle[ 3376] = 1'b0;  wr_cycle[ 3376] = 1'b1;  addr_rom[ 3376]='h000034c0;  wr_data_rom[ 3376]='h00000f8a;
    rd_cycle[ 3377] = 1'b0;  wr_cycle[ 3377] = 1'b1;  addr_rom[ 3377]='h000034c4;  wr_data_rom[ 3377]='h000021e0;
    rd_cycle[ 3378] = 1'b0;  wr_cycle[ 3378] = 1'b1;  addr_rom[ 3378]='h000034c8;  wr_data_rom[ 3378]='h00001182;
    rd_cycle[ 3379] = 1'b0;  wr_cycle[ 3379] = 1'b1;  addr_rom[ 3379]='h000034cc;  wr_data_rom[ 3379]='h000018d9;
    rd_cycle[ 3380] = 1'b0;  wr_cycle[ 3380] = 1'b1;  addr_rom[ 3380]='h000034d0;  wr_data_rom[ 3380]='h000032f1;
    rd_cycle[ 3381] = 1'b0;  wr_cycle[ 3381] = 1'b1;  addr_rom[ 3381]='h000034d4;  wr_data_rom[ 3381]='h00002147;
    rd_cycle[ 3382] = 1'b0;  wr_cycle[ 3382] = 1'b1;  addr_rom[ 3382]='h000034d8;  wr_data_rom[ 3382]='h0000034c;
    rd_cycle[ 3383] = 1'b0;  wr_cycle[ 3383] = 1'b1;  addr_rom[ 3383]='h000034dc;  wr_data_rom[ 3383]='h000006e7;
    rd_cycle[ 3384] = 1'b0;  wr_cycle[ 3384] = 1'b1;  addr_rom[ 3384]='h000034e0;  wr_data_rom[ 3384]='h00002a10;
    rd_cycle[ 3385] = 1'b0;  wr_cycle[ 3385] = 1'b1;  addr_rom[ 3385]='h000034e4;  wr_data_rom[ 3385]='h00003ebf;
    rd_cycle[ 3386] = 1'b0;  wr_cycle[ 3386] = 1'b1;  addr_rom[ 3386]='h000034e8;  wr_data_rom[ 3386]='h00002d51;
    rd_cycle[ 3387] = 1'b0;  wr_cycle[ 3387] = 1'b1;  addr_rom[ 3387]='h000034ec;  wr_data_rom[ 3387]='h000010ef;
    rd_cycle[ 3388] = 1'b0;  wr_cycle[ 3388] = 1'b1;  addr_rom[ 3388]='h000034f0;  wr_data_rom[ 3388]='h0000390c;
    rd_cycle[ 3389] = 1'b0;  wr_cycle[ 3389] = 1'b1;  addr_rom[ 3389]='h000034f4;  wr_data_rom[ 3389]='h00001a88;
    rd_cycle[ 3390] = 1'b0;  wr_cycle[ 3390] = 1'b1;  addr_rom[ 3390]='h000034f8;  wr_data_rom[ 3390]='h00002a4c;
    rd_cycle[ 3391] = 1'b0;  wr_cycle[ 3391] = 1'b1;  addr_rom[ 3391]='h000034fc;  wr_data_rom[ 3391]='h00000bcb;
    rd_cycle[ 3392] = 1'b0;  wr_cycle[ 3392] = 1'b1;  addr_rom[ 3392]='h00003500;  wr_data_rom[ 3392]='h0000231b;
    rd_cycle[ 3393] = 1'b0;  wr_cycle[ 3393] = 1'b1;  addr_rom[ 3393]='h00003504;  wr_data_rom[ 3393]='h0000158d;
    rd_cycle[ 3394] = 1'b0;  wr_cycle[ 3394] = 1'b1;  addr_rom[ 3394]='h00003508;  wr_data_rom[ 3394]='h00003025;
    rd_cycle[ 3395] = 1'b0;  wr_cycle[ 3395] = 1'b1;  addr_rom[ 3395]='h0000350c;  wr_data_rom[ 3395]='h00002204;
    rd_cycle[ 3396] = 1'b0;  wr_cycle[ 3396] = 1'b1;  addr_rom[ 3396]='h00003510;  wr_data_rom[ 3396]='h0000212b;
    rd_cycle[ 3397] = 1'b0;  wr_cycle[ 3397] = 1'b1;  addr_rom[ 3397]='h00003514;  wr_data_rom[ 3397]='h00002bc6;
    rd_cycle[ 3398] = 1'b0;  wr_cycle[ 3398] = 1'b1;  addr_rom[ 3398]='h00003518;  wr_data_rom[ 3398]='h000028c8;
    rd_cycle[ 3399] = 1'b0;  wr_cycle[ 3399] = 1'b1;  addr_rom[ 3399]='h0000351c;  wr_data_rom[ 3399]='h000004c6;
    rd_cycle[ 3400] = 1'b0;  wr_cycle[ 3400] = 1'b1;  addr_rom[ 3400]='h00003520;  wr_data_rom[ 3400]='h00002c11;
    rd_cycle[ 3401] = 1'b0;  wr_cycle[ 3401] = 1'b1;  addr_rom[ 3401]='h00003524;  wr_data_rom[ 3401]='h000022d7;
    rd_cycle[ 3402] = 1'b0;  wr_cycle[ 3402] = 1'b1;  addr_rom[ 3402]='h00003528;  wr_data_rom[ 3402]='h00001fc5;
    rd_cycle[ 3403] = 1'b0;  wr_cycle[ 3403] = 1'b1;  addr_rom[ 3403]='h0000352c;  wr_data_rom[ 3403]='h00001c2f;
    rd_cycle[ 3404] = 1'b0;  wr_cycle[ 3404] = 1'b1;  addr_rom[ 3404]='h00003530;  wr_data_rom[ 3404]='h000031f8;
    rd_cycle[ 3405] = 1'b0;  wr_cycle[ 3405] = 1'b1;  addr_rom[ 3405]='h00003534;  wr_data_rom[ 3405]='h00002f57;
    rd_cycle[ 3406] = 1'b0;  wr_cycle[ 3406] = 1'b1;  addr_rom[ 3406]='h00003538;  wr_data_rom[ 3406]='h0000048c;
    rd_cycle[ 3407] = 1'b0;  wr_cycle[ 3407] = 1'b1;  addr_rom[ 3407]='h0000353c;  wr_data_rom[ 3407]='h00003547;
    rd_cycle[ 3408] = 1'b0;  wr_cycle[ 3408] = 1'b1;  addr_rom[ 3408]='h00003540;  wr_data_rom[ 3408]='h00003bc2;
    rd_cycle[ 3409] = 1'b0;  wr_cycle[ 3409] = 1'b1;  addr_rom[ 3409]='h00003544;  wr_data_rom[ 3409]='h00002ae6;
    rd_cycle[ 3410] = 1'b0;  wr_cycle[ 3410] = 1'b1;  addr_rom[ 3410]='h00003548;  wr_data_rom[ 3410]='h00000cb7;
    rd_cycle[ 3411] = 1'b0;  wr_cycle[ 3411] = 1'b1;  addr_rom[ 3411]='h0000354c;  wr_data_rom[ 3411]='h00003447;
    rd_cycle[ 3412] = 1'b0;  wr_cycle[ 3412] = 1'b1;  addr_rom[ 3412]='h00003550;  wr_data_rom[ 3412]='h000025fd;
    rd_cycle[ 3413] = 1'b0;  wr_cycle[ 3413] = 1'b1;  addr_rom[ 3413]='h00003554;  wr_data_rom[ 3413]='h00003133;
    rd_cycle[ 3414] = 1'b0;  wr_cycle[ 3414] = 1'b1;  addr_rom[ 3414]='h00003558;  wr_data_rom[ 3414]='h00002882;
    rd_cycle[ 3415] = 1'b0;  wr_cycle[ 3415] = 1'b1;  addr_rom[ 3415]='h0000355c;  wr_data_rom[ 3415]='h00000e89;
    rd_cycle[ 3416] = 1'b0;  wr_cycle[ 3416] = 1'b1;  addr_rom[ 3416]='h00003560;  wr_data_rom[ 3416]='h0000278d;
    rd_cycle[ 3417] = 1'b0;  wr_cycle[ 3417] = 1'b1;  addr_rom[ 3417]='h00003564;  wr_data_rom[ 3417]='h00000339;
    rd_cycle[ 3418] = 1'b0;  wr_cycle[ 3418] = 1'b1;  addr_rom[ 3418]='h00003568;  wr_data_rom[ 3418]='h000032d4;
    rd_cycle[ 3419] = 1'b0;  wr_cycle[ 3419] = 1'b1;  addr_rom[ 3419]='h0000356c;  wr_data_rom[ 3419]='h0000239c;
    rd_cycle[ 3420] = 1'b0;  wr_cycle[ 3420] = 1'b1;  addr_rom[ 3420]='h00003570;  wr_data_rom[ 3420]='h000012d0;
    rd_cycle[ 3421] = 1'b0;  wr_cycle[ 3421] = 1'b1;  addr_rom[ 3421]='h00003574;  wr_data_rom[ 3421]='h0000216e;
    rd_cycle[ 3422] = 1'b0;  wr_cycle[ 3422] = 1'b1;  addr_rom[ 3422]='h00003578;  wr_data_rom[ 3422]='h00003bba;
    rd_cycle[ 3423] = 1'b0;  wr_cycle[ 3423] = 1'b1;  addr_rom[ 3423]='h0000357c;  wr_data_rom[ 3423]='h000021dd;
    rd_cycle[ 3424] = 1'b0;  wr_cycle[ 3424] = 1'b1;  addr_rom[ 3424]='h00003580;  wr_data_rom[ 3424]='h00002fb7;
    rd_cycle[ 3425] = 1'b0;  wr_cycle[ 3425] = 1'b1;  addr_rom[ 3425]='h00003584;  wr_data_rom[ 3425]='h0000183c;
    rd_cycle[ 3426] = 1'b0;  wr_cycle[ 3426] = 1'b1;  addr_rom[ 3426]='h00003588;  wr_data_rom[ 3426]='h00001380;
    rd_cycle[ 3427] = 1'b0;  wr_cycle[ 3427] = 1'b1;  addr_rom[ 3427]='h0000358c;  wr_data_rom[ 3427]='h00000f3a;
    rd_cycle[ 3428] = 1'b0;  wr_cycle[ 3428] = 1'b1;  addr_rom[ 3428]='h00003590;  wr_data_rom[ 3428]='h000025e6;
    rd_cycle[ 3429] = 1'b0;  wr_cycle[ 3429] = 1'b1;  addr_rom[ 3429]='h00003594;  wr_data_rom[ 3429]='h0000185c;
    rd_cycle[ 3430] = 1'b0;  wr_cycle[ 3430] = 1'b1;  addr_rom[ 3430]='h00003598;  wr_data_rom[ 3430]='h000020de;
    rd_cycle[ 3431] = 1'b0;  wr_cycle[ 3431] = 1'b1;  addr_rom[ 3431]='h0000359c;  wr_data_rom[ 3431]='h00000696;
    rd_cycle[ 3432] = 1'b0;  wr_cycle[ 3432] = 1'b1;  addr_rom[ 3432]='h000035a0;  wr_data_rom[ 3432]='h00000196;
    rd_cycle[ 3433] = 1'b0;  wr_cycle[ 3433] = 1'b1;  addr_rom[ 3433]='h000035a4;  wr_data_rom[ 3433]='h00003694;
    rd_cycle[ 3434] = 1'b0;  wr_cycle[ 3434] = 1'b1;  addr_rom[ 3434]='h000035a8;  wr_data_rom[ 3434]='h000023d9;
    rd_cycle[ 3435] = 1'b0;  wr_cycle[ 3435] = 1'b1;  addr_rom[ 3435]='h000035ac;  wr_data_rom[ 3435]='h000013a3;
    rd_cycle[ 3436] = 1'b0;  wr_cycle[ 3436] = 1'b1;  addr_rom[ 3436]='h000035b0;  wr_data_rom[ 3436]='h00002181;
    rd_cycle[ 3437] = 1'b0;  wr_cycle[ 3437] = 1'b1;  addr_rom[ 3437]='h000035b4;  wr_data_rom[ 3437]='h00001a98;
    rd_cycle[ 3438] = 1'b0;  wr_cycle[ 3438] = 1'b1;  addr_rom[ 3438]='h000035b8;  wr_data_rom[ 3438]='h0000193b;
    rd_cycle[ 3439] = 1'b0;  wr_cycle[ 3439] = 1'b1;  addr_rom[ 3439]='h000035bc;  wr_data_rom[ 3439]='h00000850;
    rd_cycle[ 3440] = 1'b0;  wr_cycle[ 3440] = 1'b1;  addr_rom[ 3440]='h000035c0;  wr_data_rom[ 3440]='h00000226;
    rd_cycle[ 3441] = 1'b0;  wr_cycle[ 3441] = 1'b1;  addr_rom[ 3441]='h000035c4;  wr_data_rom[ 3441]='h00001bb0;
    rd_cycle[ 3442] = 1'b0;  wr_cycle[ 3442] = 1'b1;  addr_rom[ 3442]='h000035c8;  wr_data_rom[ 3442]='h000012c0;
    rd_cycle[ 3443] = 1'b0;  wr_cycle[ 3443] = 1'b1;  addr_rom[ 3443]='h000035cc;  wr_data_rom[ 3443]='h00000aa5;
    rd_cycle[ 3444] = 1'b0;  wr_cycle[ 3444] = 1'b1;  addr_rom[ 3444]='h000035d0;  wr_data_rom[ 3444]='h00000788;
    rd_cycle[ 3445] = 1'b0;  wr_cycle[ 3445] = 1'b1;  addr_rom[ 3445]='h000035d4;  wr_data_rom[ 3445]='h00002f94;
    rd_cycle[ 3446] = 1'b0;  wr_cycle[ 3446] = 1'b1;  addr_rom[ 3446]='h000035d8;  wr_data_rom[ 3446]='h000020b1;
    rd_cycle[ 3447] = 1'b0;  wr_cycle[ 3447] = 1'b1;  addr_rom[ 3447]='h000035dc;  wr_data_rom[ 3447]='h0000053a;
    rd_cycle[ 3448] = 1'b0;  wr_cycle[ 3448] = 1'b1;  addr_rom[ 3448]='h000035e0;  wr_data_rom[ 3448]='h000026e6;
    rd_cycle[ 3449] = 1'b0;  wr_cycle[ 3449] = 1'b1;  addr_rom[ 3449]='h000035e4;  wr_data_rom[ 3449]='h00000b83;
    rd_cycle[ 3450] = 1'b0;  wr_cycle[ 3450] = 1'b1;  addr_rom[ 3450]='h000035e8;  wr_data_rom[ 3450]='h00002051;
    rd_cycle[ 3451] = 1'b0;  wr_cycle[ 3451] = 1'b1;  addr_rom[ 3451]='h000035ec;  wr_data_rom[ 3451]='h000017d4;
    rd_cycle[ 3452] = 1'b0;  wr_cycle[ 3452] = 1'b1;  addr_rom[ 3452]='h000035f0;  wr_data_rom[ 3452]='h0000052b;
    rd_cycle[ 3453] = 1'b0;  wr_cycle[ 3453] = 1'b1;  addr_rom[ 3453]='h000035f4;  wr_data_rom[ 3453]='h00001994;
    rd_cycle[ 3454] = 1'b0;  wr_cycle[ 3454] = 1'b1;  addr_rom[ 3454]='h000035f8;  wr_data_rom[ 3454]='h0000306e;
    rd_cycle[ 3455] = 1'b0;  wr_cycle[ 3455] = 1'b1;  addr_rom[ 3455]='h000035fc;  wr_data_rom[ 3455]='h00003743;
    rd_cycle[ 3456] = 1'b0;  wr_cycle[ 3456] = 1'b1;  addr_rom[ 3456]='h00003600;  wr_data_rom[ 3456]='h00001b4f;
    rd_cycle[ 3457] = 1'b0;  wr_cycle[ 3457] = 1'b1;  addr_rom[ 3457]='h00003604;  wr_data_rom[ 3457]='h00003bca;
    rd_cycle[ 3458] = 1'b0;  wr_cycle[ 3458] = 1'b1;  addr_rom[ 3458]='h00003608;  wr_data_rom[ 3458]='h00000023;
    rd_cycle[ 3459] = 1'b0;  wr_cycle[ 3459] = 1'b1;  addr_rom[ 3459]='h0000360c;  wr_data_rom[ 3459]='h00001c7c;
    rd_cycle[ 3460] = 1'b0;  wr_cycle[ 3460] = 1'b1;  addr_rom[ 3460]='h00003610;  wr_data_rom[ 3460]='h00002e80;
    rd_cycle[ 3461] = 1'b0;  wr_cycle[ 3461] = 1'b1;  addr_rom[ 3461]='h00003614;  wr_data_rom[ 3461]='h00002b1b;
    rd_cycle[ 3462] = 1'b0;  wr_cycle[ 3462] = 1'b1;  addr_rom[ 3462]='h00003618;  wr_data_rom[ 3462]='h00001682;
    rd_cycle[ 3463] = 1'b0;  wr_cycle[ 3463] = 1'b1;  addr_rom[ 3463]='h0000361c;  wr_data_rom[ 3463]='h000015cd;
    rd_cycle[ 3464] = 1'b0;  wr_cycle[ 3464] = 1'b1;  addr_rom[ 3464]='h00003620;  wr_data_rom[ 3464]='h00001266;
    rd_cycle[ 3465] = 1'b0;  wr_cycle[ 3465] = 1'b1;  addr_rom[ 3465]='h00003624;  wr_data_rom[ 3465]='h00000fdb;
    rd_cycle[ 3466] = 1'b0;  wr_cycle[ 3466] = 1'b1;  addr_rom[ 3466]='h00003628;  wr_data_rom[ 3466]='h00001857;
    rd_cycle[ 3467] = 1'b0;  wr_cycle[ 3467] = 1'b1;  addr_rom[ 3467]='h0000362c;  wr_data_rom[ 3467]='h00002f1c;
    rd_cycle[ 3468] = 1'b0;  wr_cycle[ 3468] = 1'b1;  addr_rom[ 3468]='h00003630;  wr_data_rom[ 3468]='h00002e16;
    rd_cycle[ 3469] = 1'b0;  wr_cycle[ 3469] = 1'b1;  addr_rom[ 3469]='h00003634;  wr_data_rom[ 3469]='h00001860;
    rd_cycle[ 3470] = 1'b0;  wr_cycle[ 3470] = 1'b1;  addr_rom[ 3470]='h00003638;  wr_data_rom[ 3470]='h00002b95;
    rd_cycle[ 3471] = 1'b0;  wr_cycle[ 3471] = 1'b1;  addr_rom[ 3471]='h0000363c;  wr_data_rom[ 3471]='h00003581;
    rd_cycle[ 3472] = 1'b0;  wr_cycle[ 3472] = 1'b1;  addr_rom[ 3472]='h00003640;  wr_data_rom[ 3472]='h000016c5;
    rd_cycle[ 3473] = 1'b0;  wr_cycle[ 3473] = 1'b1;  addr_rom[ 3473]='h00003644;  wr_data_rom[ 3473]='h00003677;
    rd_cycle[ 3474] = 1'b0;  wr_cycle[ 3474] = 1'b1;  addr_rom[ 3474]='h00003648;  wr_data_rom[ 3474]='h00001aa6;
    rd_cycle[ 3475] = 1'b0;  wr_cycle[ 3475] = 1'b1;  addr_rom[ 3475]='h0000364c;  wr_data_rom[ 3475]='h00000952;
    rd_cycle[ 3476] = 1'b0;  wr_cycle[ 3476] = 1'b1;  addr_rom[ 3476]='h00003650;  wr_data_rom[ 3476]='h000014e6;
    rd_cycle[ 3477] = 1'b0;  wr_cycle[ 3477] = 1'b1;  addr_rom[ 3477]='h00003654;  wr_data_rom[ 3477]='h00001289;
    rd_cycle[ 3478] = 1'b0;  wr_cycle[ 3478] = 1'b1;  addr_rom[ 3478]='h00003658;  wr_data_rom[ 3478]='h000017de;
    rd_cycle[ 3479] = 1'b0;  wr_cycle[ 3479] = 1'b1;  addr_rom[ 3479]='h0000365c;  wr_data_rom[ 3479]='h00002eec;
    rd_cycle[ 3480] = 1'b0;  wr_cycle[ 3480] = 1'b1;  addr_rom[ 3480]='h00003660;  wr_data_rom[ 3480]='h0000033f;
    rd_cycle[ 3481] = 1'b0;  wr_cycle[ 3481] = 1'b1;  addr_rom[ 3481]='h00003664;  wr_data_rom[ 3481]='h0000391a;
    rd_cycle[ 3482] = 1'b0;  wr_cycle[ 3482] = 1'b1;  addr_rom[ 3482]='h00003668;  wr_data_rom[ 3482]='h0000308b;
    rd_cycle[ 3483] = 1'b0;  wr_cycle[ 3483] = 1'b1;  addr_rom[ 3483]='h0000366c;  wr_data_rom[ 3483]='h00003019;
    rd_cycle[ 3484] = 1'b0;  wr_cycle[ 3484] = 1'b1;  addr_rom[ 3484]='h00003670;  wr_data_rom[ 3484]='h00001be8;
    rd_cycle[ 3485] = 1'b0;  wr_cycle[ 3485] = 1'b1;  addr_rom[ 3485]='h00003674;  wr_data_rom[ 3485]='h00001d03;
    rd_cycle[ 3486] = 1'b0;  wr_cycle[ 3486] = 1'b1;  addr_rom[ 3486]='h00003678;  wr_data_rom[ 3486]='h00003569;
    rd_cycle[ 3487] = 1'b0;  wr_cycle[ 3487] = 1'b1;  addr_rom[ 3487]='h0000367c;  wr_data_rom[ 3487]='h00003e73;
    rd_cycle[ 3488] = 1'b0;  wr_cycle[ 3488] = 1'b1;  addr_rom[ 3488]='h00003680;  wr_data_rom[ 3488]='h0000031c;
    rd_cycle[ 3489] = 1'b0;  wr_cycle[ 3489] = 1'b1;  addr_rom[ 3489]='h00003684;  wr_data_rom[ 3489]='h0000185b;
    rd_cycle[ 3490] = 1'b0;  wr_cycle[ 3490] = 1'b1;  addr_rom[ 3490]='h00003688;  wr_data_rom[ 3490]='h00003f9d;
    rd_cycle[ 3491] = 1'b0;  wr_cycle[ 3491] = 1'b1;  addr_rom[ 3491]='h0000368c;  wr_data_rom[ 3491]='h0000182a;
    rd_cycle[ 3492] = 1'b0;  wr_cycle[ 3492] = 1'b1;  addr_rom[ 3492]='h00003690;  wr_data_rom[ 3492]='h000029a3;
    rd_cycle[ 3493] = 1'b0;  wr_cycle[ 3493] = 1'b1;  addr_rom[ 3493]='h00003694;  wr_data_rom[ 3493]='h00002651;
    rd_cycle[ 3494] = 1'b0;  wr_cycle[ 3494] = 1'b1;  addr_rom[ 3494]='h00003698;  wr_data_rom[ 3494]='h000008c3;
    rd_cycle[ 3495] = 1'b0;  wr_cycle[ 3495] = 1'b1;  addr_rom[ 3495]='h0000369c;  wr_data_rom[ 3495]='h00000ad6;
    rd_cycle[ 3496] = 1'b0;  wr_cycle[ 3496] = 1'b1;  addr_rom[ 3496]='h000036a0;  wr_data_rom[ 3496]='h00000515;
    rd_cycle[ 3497] = 1'b0;  wr_cycle[ 3497] = 1'b1;  addr_rom[ 3497]='h000036a4;  wr_data_rom[ 3497]='h00003448;
    rd_cycle[ 3498] = 1'b0;  wr_cycle[ 3498] = 1'b1;  addr_rom[ 3498]='h000036a8;  wr_data_rom[ 3498]='h000007a8;
    rd_cycle[ 3499] = 1'b0;  wr_cycle[ 3499] = 1'b1;  addr_rom[ 3499]='h000036ac;  wr_data_rom[ 3499]='h000023aa;
    rd_cycle[ 3500] = 1'b0;  wr_cycle[ 3500] = 1'b1;  addr_rom[ 3500]='h000036b0;  wr_data_rom[ 3500]='h00001699;
    rd_cycle[ 3501] = 1'b0;  wr_cycle[ 3501] = 1'b1;  addr_rom[ 3501]='h000036b4;  wr_data_rom[ 3501]='h00002346;
    rd_cycle[ 3502] = 1'b0;  wr_cycle[ 3502] = 1'b1;  addr_rom[ 3502]='h000036b8;  wr_data_rom[ 3502]='h00002382;
    rd_cycle[ 3503] = 1'b0;  wr_cycle[ 3503] = 1'b1;  addr_rom[ 3503]='h000036bc;  wr_data_rom[ 3503]='h0000337d;
    rd_cycle[ 3504] = 1'b0;  wr_cycle[ 3504] = 1'b1;  addr_rom[ 3504]='h000036c0;  wr_data_rom[ 3504]='h000005a2;
    rd_cycle[ 3505] = 1'b0;  wr_cycle[ 3505] = 1'b1;  addr_rom[ 3505]='h000036c4;  wr_data_rom[ 3505]='h00002985;
    rd_cycle[ 3506] = 1'b0;  wr_cycle[ 3506] = 1'b1;  addr_rom[ 3506]='h000036c8;  wr_data_rom[ 3506]='h00002916;
    rd_cycle[ 3507] = 1'b0;  wr_cycle[ 3507] = 1'b1;  addr_rom[ 3507]='h000036cc;  wr_data_rom[ 3507]='h000032a3;
    rd_cycle[ 3508] = 1'b0;  wr_cycle[ 3508] = 1'b1;  addr_rom[ 3508]='h000036d0;  wr_data_rom[ 3508]='h0000194b;
    rd_cycle[ 3509] = 1'b0;  wr_cycle[ 3509] = 1'b1;  addr_rom[ 3509]='h000036d4;  wr_data_rom[ 3509]='h000008ef;
    rd_cycle[ 3510] = 1'b0;  wr_cycle[ 3510] = 1'b1;  addr_rom[ 3510]='h000036d8;  wr_data_rom[ 3510]='h000005bd;
    rd_cycle[ 3511] = 1'b0;  wr_cycle[ 3511] = 1'b1;  addr_rom[ 3511]='h000036dc;  wr_data_rom[ 3511]='h00001fb3;
    rd_cycle[ 3512] = 1'b0;  wr_cycle[ 3512] = 1'b1;  addr_rom[ 3512]='h000036e0;  wr_data_rom[ 3512]='h00003912;
    rd_cycle[ 3513] = 1'b0;  wr_cycle[ 3513] = 1'b1;  addr_rom[ 3513]='h000036e4;  wr_data_rom[ 3513]='h00001984;
    rd_cycle[ 3514] = 1'b0;  wr_cycle[ 3514] = 1'b1;  addr_rom[ 3514]='h000036e8;  wr_data_rom[ 3514]='h00002548;
    rd_cycle[ 3515] = 1'b0;  wr_cycle[ 3515] = 1'b1;  addr_rom[ 3515]='h000036ec;  wr_data_rom[ 3515]='h00002f19;
    rd_cycle[ 3516] = 1'b0;  wr_cycle[ 3516] = 1'b1;  addr_rom[ 3516]='h000036f0;  wr_data_rom[ 3516]='h00000b55;
    rd_cycle[ 3517] = 1'b0;  wr_cycle[ 3517] = 1'b1;  addr_rom[ 3517]='h000036f4;  wr_data_rom[ 3517]='h000035ac;
    rd_cycle[ 3518] = 1'b0;  wr_cycle[ 3518] = 1'b1;  addr_rom[ 3518]='h000036f8;  wr_data_rom[ 3518]='h00001f95;
    rd_cycle[ 3519] = 1'b0;  wr_cycle[ 3519] = 1'b1;  addr_rom[ 3519]='h000036fc;  wr_data_rom[ 3519]='h00000cad;
    rd_cycle[ 3520] = 1'b0;  wr_cycle[ 3520] = 1'b1;  addr_rom[ 3520]='h00003700;  wr_data_rom[ 3520]='h0000187d;
    rd_cycle[ 3521] = 1'b0;  wr_cycle[ 3521] = 1'b1;  addr_rom[ 3521]='h00003704;  wr_data_rom[ 3521]='h000012e1;
    rd_cycle[ 3522] = 1'b0;  wr_cycle[ 3522] = 1'b1;  addr_rom[ 3522]='h00003708;  wr_data_rom[ 3522]='h000004d0;
    rd_cycle[ 3523] = 1'b0;  wr_cycle[ 3523] = 1'b1;  addr_rom[ 3523]='h0000370c;  wr_data_rom[ 3523]='h00000830;
    rd_cycle[ 3524] = 1'b0;  wr_cycle[ 3524] = 1'b1;  addr_rom[ 3524]='h00003710;  wr_data_rom[ 3524]='h00000381;
    rd_cycle[ 3525] = 1'b0;  wr_cycle[ 3525] = 1'b1;  addr_rom[ 3525]='h00003714;  wr_data_rom[ 3525]='h00000561;
    rd_cycle[ 3526] = 1'b0;  wr_cycle[ 3526] = 1'b1;  addr_rom[ 3526]='h00003718;  wr_data_rom[ 3526]='h000025f9;
    rd_cycle[ 3527] = 1'b0;  wr_cycle[ 3527] = 1'b1;  addr_rom[ 3527]='h0000371c;  wr_data_rom[ 3527]='h000037cd;
    rd_cycle[ 3528] = 1'b0;  wr_cycle[ 3528] = 1'b1;  addr_rom[ 3528]='h00003720;  wr_data_rom[ 3528]='h00001f8d;
    rd_cycle[ 3529] = 1'b0;  wr_cycle[ 3529] = 1'b1;  addr_rom[ 3529]='h00003724;  wr_data_rom[ 3529]='h00003e16;
    rd_cycle[ 3530] = 1'b0;  wr_cycle[ 3530] = 1'b1;  addr_rom[ 3530]='h00003728;  wr_data_rom[ 3530]='h0000293e;
    rd_cycle[ 3531] = 1'b0;  wr_cycle[ 3531] = 1'b1;  addr_rom[ 3531]='h0000372c;  wr_data_rom[ 3531]='h000024da;
    rd_cycle[ 3532] = 1'b0;  wr_cycle[ 3532] = 1'b1;  addr_rom[ 3532]='h00003730;  wr_data_rom[ 3532]='h00000a71;
    rd_cycle[ 3533] = 1'b0;  wr_cycle[ 3533] = 1'b1;  addr_rom[ 3533]='h00003734;  wr_data_rom[ 3533]='h0000354f;
    rd_cycle[ 3534] = 1'b0;  wr_cycle[ 3534] = 1'b1;  addr_rom[ 3534]='h00003738;  wr_data_rom[ 3534]='h0000095b;
    rd_cycle[ 3535] = 1'b0;  wr_cycle[ 3535] = 1'b1;  addr_rom[ 3535]='h0000373c;  wr_data_rom[ 3535]='h000033cd;
    rd_cycle[ 3536] = 1'b0;  wr_cycle[ 3536] = 1'b1;  addr_rom[ 3536]='h00003740;  wr_data_rom[ 3536]='h00000a36;
    rd_cycle[ 3537] = 1'b0;  wr_cycle[ 3537] = 1'b1;  addr_rom[ 3537]='h00003744;  wr_data_rom[ 3537]='h000027ff;
    rd_cycle[ 3538] = 1'b0;  wr_cycle[ 3538] = 1'b1;  addr_rom[ 3538]='h00003748;  wr_data_rom[ 3538]='h00000aad;
    rd_cycle[ 3539] = 1'b0;  wr_cycle[ 3539] = 1'b1;  addr_rom[ 3539]='h0000374c;  wr_data_rom[ 3539]='h0000305c;
    rd_cycle[ 3540] = 1'b0;  wr_cycle[ 3540] = 1'b1;  addr_rom[ 3540]='h00003750;  wr_data_rom[ 3540]='h0000196d;
    rd_cycle[ 3541] = 1'b0;  wr_cycle[ 3541] = 1'b1;  addr_rom[ 3541]='h00003754;  wr_data_rom[ 3541]='h00001932;
    rd_cycle[ 3542] = 1'b0;  wr_cycle[ 3542] = 1'b1;  addr_rom[ 3542]='h00003758;  wr_data_rom[ 3542]='h00002a7b;
    rd_cycle[ 3543] = 1'b0;  wr_cycle[ 3543] = 1'b1;  addr_rom[ 3543]='h0000375c;  wr_data_rom[ 3543]='h00003e6e;
    rd_cycle[ 3544] = 1'b0;  wr_cycle[ 3544] = 1'b1;  addr_rom[ 3544]='h00003760;  wr_data_rom[ 3544]='h000035ce;
    rd_cycle[ 3545] = 1'b0;  wr_cycle[ 3545] = 1'b1;  addr_rom[ 3545]='h00003764;  wr_data_rom[ 3545]='h00001506;
    rd_cycle[ 3546] = 1'b0;  wr_cycle[ 3546] = 1'b1;  addr_rom[ 3546]='h00003768;  wr_data_rom[ 3546]='h00000b06;
    rd_cycle[ 3547] = 1'b0;  wr_cycle[ 3547] = 1'b1;  addr_rom[ 3547]='h0000376c;  wr_data_rom[ 3547]='h000005ca;
    rd_cycle[ 3548] = 1'b0;  wr_cycle[ 3548] = 1'b1;  addr_rom[ 3548]='h00003770;  wr_data_rom[ 3548]='h000025c0;
    rd_cycle[ 3549] = 1'b0;  wr_cycle[ 3549] = 1'b1;  addr_rom[ 3549]='h00003774;  wr_data_rom[ 3549]='h00001111;
    rd_cycle[ 3550] = 1'b0;  wr_cycle[ 3550] = 1'b1;  addr_rom[ 3550]='h00003778;  wr_data_rom[ 3550]='h000024c9;
    rd_cycle[ 3551] = 1'b0;  wr_cycle[ 3551] = 1'b1;  addr_rom[ 3551]='h0000377c;  wr_data_rom[ 3551]='h00003bab;
    rd_cycle[ 3552] = 1'b0;  wr_cycle[ 3552] = 1'b1;  addr_rom[ 3552]='h00003780;  wr_data_rom[ 3552]='h00002a03;
    rd_cycle[ 3553] = 1'b0;  wr_cycle[ 3553] = 1'b1;  addr_rom[ 3553]='h00003784;  wr_data_rom[ 3553]='h0000050a;
    rd_cycle[ 3554] = 1'b0;  wr_cycle[ 3554] = 1'b1;  addr_rom[ 3554]='h00003788;  wr_data_rom[ 3554]='h000019e0;
    rd_cycle[ 3555] = 1'b0;  wr_cycle[ 3555] = 1'b1;  addr_rom[ 3555]='h0000378c;  wr_data_rom[ 3555]='h000015c7;
    rd_cycle[ 3556] = 1'b0;  wr_cycle[ 3556] = 1'b1;  addr_rom[ 3556]='h00003790;  wr_data_rom[ 3556]='h00002871;
    rd_cycle[ 3557] = 1'b0;  wr_cycle[ 3557] = 1'b1;  addr_rom[ 3557]='h00003794;  wr_data_rom[ 3557]='h00000393;
    rd_cycle[ 3558] = 1'b0;  wr_cycle[ 3558] = 1'b1;  addr_rom[ 3558]='h00003798;  wr_data_rom[ 3558]='h0000095d;
    rd_cycle[ 3559] = 1'b0;  wr_cycle[ 3559] = 1'b1;  addr_rom[ 3559]='h0000379c;  wr_data_rom[ 3559]='h000021ba;
    rd_cycle[ 3560] = 1'b0;  wr_cycle[ 3560] = 1'b1;  addr_rom[ 3560]='h000037a0;  wr_data_rom[ 3560]='h00001276;
    rd_cycle[ 3561] = 1'b0;  wr_cycle[ 3561] = 1'b1;  addr_rom[ 3561]='h000037a4;  wr_data_rom[ 3561]='h000029b5;
    rd_cycle[ 3562] = 1'b0;  wr_cycle[ 3562] = 1'b1;  addr_rom[ 3562]='h000037a8;  wr_data_rom[ 3562]='h00000c7e;
    rd_cycle[ 3563] = 1'b0;  wr_cycle[ 3563] = 1'b1;  addr_rom[ 3563]='h000037ac;  wr_data_rom[ 3563]='h00000cf9;
    rd_cycle[ 3564] = 1'b0;  wr_cycle[ 3564] = 1'b1;  addr_rom[ 3564]='h000037b0;  wr_data_rom[ 3564]='h000021b8;
    rd_cycle[ 3565] = 1'b0;  wr_cycle[ 3565] = 1'b1;  addr_rom[ 3565]='h000037b4;  wr_data_rom[ 3565]='h00003a2a;
    rd_cycle[ 3566] = 1'b0;  wr_cycle[ 3566] = 1'b1;  addr_rom[ 3566]='h000037b8;  wr_data_rom[ 3566]='h000026a0;
    rd_cycle[ 3567] = 1'b0;  wr_cycle[ 3567] = 1'b1;  addr_rom[ 3567]='h000037bc;  wr_data_rom[ 3567]='h00000f4c;
    rd_cycle[ 3568] = 1'b0;  wr_cycle[ 3568] = 1'b1;  addr_rom[ 3568]='h000037c0;  wr_data_rom[ 3568]='h00002832;
    rd_cycle[ 3569] = 1'b0;  wr_cycle[ 3569] = 1'b1;  addr_rom[ 3569]='h000037c4;  wr_data_rom[ 3569]='h00003b5c;
    rd_cycle[ 3570] = 1'b0;  wr_cycle[ 3570] = 1'b1;  addr_rom[ 3570]='h000037c8;  wr_data_rom[ 3570]='h000031a4;
    rd_cycle[ 3571] = 1'b0;  wr_cycle[ 3571] = 1'b1;  addr_rom[ 3571]='h000037cc;  wr_data_rom[ 3571]='h00001a16;
    rd_cycle[ 3572] = 1'b0;  wr_cycle[ 3572] = 1'b1;  addr_rom[ 3572]='h000037d0;  wr_data_rom[ 3572]='h00000c3b;
    rd_cycle[ 3573] = 1'b0;  wr_cycle[ 3573] = 1'b1;  addr_rom[ 3573]='h000037d4;  wr_data_rom[ 3573]='h00001663;
    rd_cycle[ 3574] = 1'b0;  wr_cycle[ 3574] = 1'b1;  addr_rom[ 3574]='h000037d8;  wr_data_rom[ 3574]='h00002f47;
    rd_cycle[ 3575] = 1'b0;  wr_cycle[ 3575] = 1'b1;  addr_rom[ 3575]='h000037dc;  wr_data_rom[ 3575]='h00002be4;
    rd_cycle[ 3576] = 1'b0;  wr_cycle[ 3576] = 1'b1;  addr_rom[ 3576]='h000037e0;  wr_data_rom[ 3576]='h000010b2;
    rd_cycle[ 3577] = 1'b0;  wr_cycle[ 3577] = 1'b1;  addr_rom[ 3577]='h000037e4;  wr_data_rom[ 3577]='h00001cd4;
    rd_cycle[ 3578] = 1'b0;  wr_cycle[ 3578] = 1'b1;  addr_rom[ 3578]='h000037e8;  wr_data_rom[ 3578]='h00001a13;
    rd_cycle[ 3579] = 1'b0;  wr_cycle[ 3579] = 1'b1;  addr_rom[ 3579]='h000037ec;  wr_data_rom[ 3579]='h0000064d;
    rd_cycle[ 3580] = 1'b0;  wr_cycle[ 3580] = 1'b1;  addr_rom[ 3580]='h000037f0;  wr_data_rom[ 3580]='h000004e3;
    rd_cycle[ 3581] = 1'b0;  wr_cycle[ 3581] = 1'b1;  addr_rom[ 3581]='h000037f4;  wr_data_rom[ 3581]='h000039db;
    rd_cycle[ 3582] = 1'b0;  wr_cycle[ 3582] = 1'b1;  addr_rom[ 3582]='h000037f8;  wr_data_rom[ 3582]='h00002f77;
    rd_cycle[ 3583] = 1'b0;  wr_cycle[ 3583] = 1'b1;  addr_rom[ 3583]='h000037fc;  wr_data_rom[ 3583]='h00000b84;
    rd_cycle[ 3584] = 1'b0;  wr_cycle[ 3584] = 1'b1;  addr_rom[ 3584]='h00003800;  wr_data_rom[ 3584]='h0000334f;
    rd_cycle[ 3585] = 1'b0;  wr_cycle[ 3585] = 1'b1;  addr_rom[ 3585]='h00003804;  wr_data_rom[ 3585]='h00002cb6;
    rd_cycle[ 3586] = 1'b0;  wr_cycle[ 3586] = 1'b1;  addr_rom[ 3586]='h00003808;  wr_data_rom[ 3586]='h00002a17;
    rd_cycle[ 3587] = 1'b0;  wr_cycle[ 3587] = 1'b1;  addr_rom[ 3587]='h0000380c;  wr_data_rom[ 3587]='h00002da2;
    rd_cycle[ 3588] = 1'b0;  wr_cycle[ 3588] = 1'b1;  addr_rom[ 3588]='h00003810;  wr_data_rom[ 3588]='h00000a97;
    rd_cycle[ 3589] = 1'b0;  wr_cycle[ 3589] = 1'b1;  addr_rom[ 3589]='h00003814;  wr_data_rom[ 3589]='h000023c3;
    rd_cycle[ 3590] = 1'b0;  wr_cycle[ 3590] = 1'b1;  addr_rom[ 3590]='h00003818;  wr_data_rom[ 3590]='h000021ba;
    rd_cycle[ 3591] = 1'b0;  wr_cycle[ 3591] = 1'b1;  addr_rom[ 3591]='h0000381c;  wr_data_rom[ 3591]='h00003eee;
    rd_cycle[ 3592] = 1'b0;  wr_cycle[ 3592] = 1'b1;  addr_rom[ 3592]='h00003820;  wr_data_rom[ 3592]='h000015b3;
    rd_cycle[ 3593] = 1'b0;  wr_cycle[ 3593] = 1'b1;  addr_rom[ 3593]='h00003824;  wr_data_rom[ 3593]='h00002b4b;
    rd_cycle[ 3594] = 1'b0;  wr_cycle[ 3594] = 1'b1;  addr_rom[ 3594]='h00003828;  wr_data_rom[ 3594]='h000008c2;
    rd_cycle[ 3595] = 1'b0;  wr_cycle[ 3595] = 1'b1;  addr_rom[ 3595]='h0000382c;  wr_data_rom[ 3595]='h000019ca;
    rd_cycle[ 3596] = 1'b0;  wr_cycle[ 3596] = 1'b1;  addr_rom[ 3596]='h00003830;  wr_data_rom[ 3596]='h0000154b;
    rd_cycle[ 3597] = 1'b0;  wr_cycle[ 3597] = 1'b1;  addr_rom[ 3597]='h00003834;  wr_data_rom[ 3597]='h00001e4a;
    rd_cycle[ 3598] = 1'b0;  wr_cycle[ 3598] = 1'b1;  addr_rom[ 3598]='h00003838;  wr_data_rom[ 3598]='h000018ad;
    rd_cycle[ 3599] = 1'b0;  wr_cycle[ 3599] = 1'b1;  addr_rom[ 3599]='h0000383c;  wr_data_rom[ 3599]='h00001e32;
    rd_cycle[ 3600] = 1'b0;  wr_cycle[ 3600] = 1'b1;  addr_rom[ 3600]='h00003840;  wr_data_rom[ 3600]='h000007e0;
    rd_cycle[ 3601] = 1'b0;  wr_cycle[ 3601] = 1'b1;  addr_rom[ 3601]='h00003844;  wr_data_rom[ 3601]='h000002c4;
    rd_cycle[ 3602] = 1'b0;  wr_cycle[ 3602] = 1'b1;  addr_rom[ 3602]='h00003848;  wr_data_rom[ 3602]='h0000319c;
    rd_cycle[ 3603] = 1'b0;  wr_cycle[ 3603] = 1'b1;  addr_rom[ 3603]='h0000384c;  wr_data_rom[ 3603]='h00001eb2;
    rd_cycle[ 3604] = 1'b0;  wr_cycle[ 3604] = 1'b1;  addr_rom[ 3604]='h00003850;  wr_data_rom[ 3604]='h00000fd1;
    rd_cycle[ 3605] = 1'b0;  wr_cycle[ 3605] = 1'b1;  addr_rom[ 3605]='h00003854;  wr_data_rom[ 3605]='h00003d1b;
    rd_cycle[ 3606] = 1'b0;  wr_cycle[ 3606] = 1'b1;  addr_rom[ 3606]='h00003858;  wr_data_rom[ 3606]='h00001247;
    rd_cycle[ 3607] = 1'b0;  wr_cycle[ 3607] = 1'b1;  addr_rom[ 3607]='h0000385c;  wr_data_rom[ 3607]='h00002617;
    rd_cycle[ 3608] = 1'b0;  wr_cycle[ 3608] = 1'b1;  addr_rom[ 3608]='h00003860;  wr_data_rom[ 3608]='h00002c8f;
    rd_cycle[ 3609] = 1'b0;  wr_cycle[ 3609] = 1'b1;  addr_rom[ 3609]='h00003864;  wr_data_rom[ 3609]='h00000feb;
    rd_cycle[ 3610] = 1'b0;  wr_cycle[ 3610] = 1'b1;  addr_rom[ 3610]='h00003868;  wr_data_rom[ 3610]='h00002f82;
    rd_cycle[ 3611] = 1'b0;  wr_cycle[ 3611] = 1'b1;  addr_rom[ 3611]='h0000386c;  wr_data_rom[ 3611]='h00002a57;
    rd_cycle[ 3612] = 1'b0;  wr_cycle[ 3612] = 1'b1;  addr_rom[ 3612]='h00003870;  wr_data_rom[ 3612]='h000006e2;
    rd_cycle[ 3613] = 1'b0;  wr_cycle[ 3613] = 1'b1;  addr_rom[ 3613]='h00003874;  wr_data_rom[ 3613]='h00000c0e;
    rd_cycle[ 3614] = 1'b0;  wr_cycle[ 3614] = 1'b1;  addr_rom[ 3614]='h00003878;  wr_data_rom[ 3614]='h00002ebe;
    rd_cycle[ 3615] = 1'b0;  wr_cycle[ 3615] = 1'b1;  addr_rom[ 3615]='h0000387c;  wr_data_rom[ 3615]='h000017cb;
    rd_cycle[ 3616] = 1'b0;  wr_cycle[ 3616] = 1'b1;  addr_rom[ 3616]='h00003880;  wr_data_rom[ 3616]='h0000041c;
    rd_cycle[ 3617] = 1'b0;  wr_cycle[ 3617] = 1'b1;  addr_rom[ 3617]='h00003884;  wr_data_rom[ 3617]='h0000045a;
    rd_cycle[ 3618] = 1'b0;  wr_cycle[ 3618] = 1'b1;  addr_rom[ 3618]='h00003888;  wr_data_rom[ 3618]='h00001fef;
    rd_cycle[ 3619] = 1'b0;  wr_cycle[ 3619] = 1'b1;  addr_rom[ 3619]='h0000388c;  wr_data_rom[ 3619]='h00001966;
    rd_cycle[ 3620] = 1'b0;  wr_cycle[ 3620] = 1'b1;  addr_rom[ 3620]='h00003890;  wr_data_rom[ 3620]='h000032b6;
    rd_cycle[ 3621] = 1'b0;  wr_cycle[ 3621] = 1'b1;  addr_rom[ 3621]='h00003894;  wr_data_rom[ 3621]='h00000fea;
    rd_cycle[ 3622] = 1'b0;  wr_cycle[ 3622] = 1'b1;  addr_rom[ 3622]='h00003898;  wr_data_rom[ 3622]='h00003cc9;
    rd_cycle[ 3623] = 1'b0;  wr_cycle[ 3623] = 1'b1;  addr_rom[ 3623]='h0000389c;  wr_data_rom[ 3623]='h00001290;
    rd_cycle[ 3624] = 1'b0;  wr_cycle[ 3624] = 1'b1;  addr_rom[ 3624]='h000038a0;  wr_data_rom[ 3624]='h000028e7;
    rd_cycle[ 3625] = 1'b0;  wr_cycle[ 3625] = 1'b1;  addr_rom[ 3625]='h000038a4;  wr_data_rom[ 3625]='h00001610;
    rd_cycle[ 3626] = 1'b0;  wr_cycle[ 3626] = 1'b1;  addr_rom[ 3626]='h000038a8;  wr_data_rom[ 3626]='h00001365;
    rd_cycle[ 3627] = 1'b0;  wr_cycle[ 3627] = 1'b1;  addr_rom[ 3627]='h000038ac;  wr_data_rom[ 3627]='h00001b26;
    rd_cycle[ 3628] = 1'b0;  wr_cycle[ 3628] = 1'b1;  addr_rom[ 3628]='h000038b0;  wr_data_rom[ 3628]='h000030fa;
    rd_cycle[ 3629] = 1'b0;  wr_cycle[ 3629] = 1'b1;  addr_rom[ 3629]='h000038b4;  wr_data_rom[ 3629]='h00000f2a;
    rd_cycle[ 3630] = 1'b0;  wr_cycle[ 3630] = 1'b1;  addr_rom[ 3630]='h000038b8;  wr_data_rom[ 3630]='h00000fe5;
    rd_cycle[ 3631] = 1'b0;  wr_cycle[ 3631] = 1'b1;  addr_rom[ 3631]='h000038bc;  wr_data_rom[ 3631]='h000021d7;
    rd_cycle[ 3632] = 1'b0;  wr_cycle[ 3632] = 1'b1;  addr_rom[ 3632]='h000038c0;  wr_data_rom[ 3632]='h00002862;
    rd_cycle[ 3633] = 1'b0;  wr_cycle[ 3633] = 1'b1;  addr_rom[ 3633]='h000038c4;  wr_data_rom[ 3633]='h00002167;
    rd_cycle[ 3634] = 1'b0;  wr_cycle[ 3634] = 1'b1;  addr_rom[ 3634]='h000038c8;  wr_data_rom[ 3634]='h00001e29;
    rd_cycle[ 3635] = 1'b0;  wr_cycle[ 3635] = 1'b1;  addr_rom[ 3635]='h000038cc;  wr_data_rom[ 3635]='h000009dd;
    rd_cycle[ 3636] = 1'b0;  wr_cycle[ 3636] = 1'b1;  addr_rom[ 3636]='h000038d0;  wr_data_rom[ 3636]='h00002b85;
    rd_cycle[ 3637] = 1'b0;  wr_cycle[ 3637] = 1'b1;  addr_rom[ 3637]='h000038d4;  wr_data_rom[ 3637]='h00002c65;
    rd_cycle[ 3638] = 1'b0;  wr_cycle[ 3638] = 1'b1;  addr_rom[ 3638]='h000038d8;  wr_data_rom[ 3638]='h0000346e;
    rd_cycle[ 3639] = 1'b0;  wr_cycle[ 3639] = 1'b1;  addr_rom[ 3639]='h000038dc;  wr_data_rom[ 3639]='h00002f28;
    rd_cycle[ 3640] = 1'b0;  wr_cycle[ 3640] = 1'b1;  addr_rom[ 3640]='h000038e0;  wr_data_rom[ 3640]='h000006a1;
    rd_cycle[ 3641] = 1'b0;  wr_cycle[ 3641] = 1'b1;  addr_rom[ 3641]='h000038e4;  wr_data_rom[ 3641]='h0000392f;
    rd_cycle[ 3642] = 1'b0;  wr_cycle[ 3642] = 1'b1;  addr_rom[ 3642]='h000038e8;  wr_data_rom[ 3642]='h00003258;
    rd_cycle[ 3643] = 1'b0;  wr_cycle[ 3643] = 1'b1;  addr_rom[ 3643]='h000038ec;  wr_data_rom[ 3643]='h000028f2;
    rd_cycle[ 3644] = 1'b0;  wr_cycle[ 3644] = 1'b1;  addr_rom[ 3644]='h000038f0;  wr_data_rom[ 3644]='h00001ac4;
    rd_cycle[ 3645] = 1'b0;  wr_cycle[ 3645] = 1'b1;  addr_rom[ 3645]='h000038f4;  wr_data_rom[ 3645]='h000030b6;
    rd_cycle[ 3646] = 1'b0;  wr_cycle[ 3646] = 1'b1;  addr_rom[ 3646]='h000038f8;  wr_data_rom[ 3646]='h00000b7b;
    rd_cycle[ 3647] = 1'b0;  wr_cycle[ 3647] = 1'b1;  addr_rom[ 3647]='h000038fc;  wr_data_rom[ 3647]='h0000360d;
    rd_cycle[ 3648] = 1'b0;  wr_cycle[ 3648] = 1'b1;  addr_rom[ 3648]='h00003900;  wr_data_rom[ 3648]='h00000df7;
    rd_cycle[ 3649] = 1'b0;  wr_cycle[ 3649] = 1'b1;  addr_rom[ 3649]='h00003904;  wr_data_rom[ 3649]='h0000021f;
    rd_cycle[ 3650] = 1'b0;  wr_cycle[ 3650] = 1'b1;  addr_rom[ 3650]='h00003908;  wr_data_rom[ 3650]='h000012c7;
    rd_cycle[ 3651] = 1'b0;  wr_cycle[ 3651] = 1'b1;  addr_rom[ 3651]='h0000390c;  wr_data_rom[ 3651]='h000023ca;
    rd_cycle[ 3652] = 1'b0;  wr_cycle[ 3652] = 1'b1;  addr_rom[ 3652]='h00003910;  wr_data_rom[ 3652]='h000005e2;
    rd_cycle[ 3653] = 1'b0;  wr_cycle[ 3653] = 1'b1;  addr_rom[ 3653]='h00003914;  wr_data_rom[ 3653]='h000027bc;
    rd_cycle[ 3654] = 1'b0;  wr_cycle[ 3654] = 1'b1;  addr_rom[ 3654]='h00003918;  wr_data_rom[ 3654]='h00000477;
    rd_cycle[ 3655] = 1'b0;  wr_cycle[ 3655] = 1'b1;  addr_rom[ 3655]='h0000391c;  wr_data_rom[ 3655]='h00003748;
    rd_cycle[ 3656] = 1'b0;  wr_cycle[ 3656] = 1'b1;  addr_rom[ 3656]='h00003920;  wr_data_rom[ 3656]='h00001183;
    rd_cycle[ 3657] = 1'b0;  wr_cycle[ 3657] = 1'b1;  addr_rom[ 3657]='h00003924;  wr_data_rom[ 3657]='h00003ed2;
    rd_cycle[ 3658] = 1'b0;  wr_cycle[ 3658] = 1'b1;  addr_rom[ 3658]='h00003928;  wr_data_rom[ 3658]='h00002c19;
    rd_cycle[ 3659] = 1'b0;  wr_cycle[ 3659] = 1'b1;  addr_rom[ 3659]='h0000392c;  wr_data_rom[ 3659]='h00000790;
    rd_cycle[ 3660] = 1'b0;  wr_cycle[ 3660] = 1'b1;  addr_rom[ 3660]='h00003930;  wr_data_rom[ 3660]='h0000176a;
    rd_cycle[ 3661] = 1'b0;  wr_cycle[ 3661] = 1'b1;  addr_rom[ 3661]='h00003934;  wr_data_rom[ 3661]='h00000138;
    rd_cycle[ 3662] = 1'b0;  wr_cycle[ 3662] = 1'b1;  addr_rom[ 3662]='h00003938;  wr_data_rom[ 3662]='h000034f6;
    rd_cycle[ 3663] = 1'b0;  wr_cycle[ 3663] = 1'b1;  addr_rom[ 3663]='h0000393c;  wr_data_rom[ 3663]='h000034a9;
    rd_cycle[ 3664] = 1'b0;  wr_cycle[ 3664] = 1'b1;  addr_rom[ 3664]='h00003940;  wr_data_rom[ 3664]='h000014ac;
    rd_cycle[ 3665] = 1'b0;  wr_cycle[ 3665] = 1'b1;  addr_rom[ 3665]='h00003944;  wr_data_rom[ 3665]='h00001f60;
    rd_cycle[ 3666] = 1'b0;  wr_cycle[ 3666] = 1'b1;  addr_rom[ 3666]='h00003948;  wr_data_rom[ 3666]='h00002aa5;
    rd_cycle[ 3667] = 1'b0;  wr_cycle[ 3667] = 1'b1;  addr_rom[ 3667]='h0000394c;  wr_data_rom[ 3667]='h000017ed;
    rd_cycle[ 3668] = 1'b0;  wr_cycle[ 3668] = 1'b1;  addr_rom[ 3668]='h00003950;  wr_data_rom[ 3668]='h0000199f;
    rd_cycle[ 3669] = 1'b0;  wr_cycle[ 3669] = 1'b1;  addr_rom[ 3669]='h00003954;  wr_data_rom[ 3669]='h00003c74;
    rd_cycle[ 3670] = 1'b0;  wr_cycle[ 3670] = 1'b1;  addr_rom[ 3670]='h00003958;  wr_data_rom[ 3670]='h0000103b;
    rd_cycle[ 3671] = 1'b0;  wr_cycle[ 3671] = 1'b1;  addr_rom[ 3671]='h0000395c;  wr_data_rom[ 3671]='h00002139;
    rd_cycle[ 3672] = 1'b0;  wr_cycle[ 3672] = 1'b1;  addr_rom[ 3672]='h00003960;  wr_data_rom[ 3672]='h00000d97;
    rd_cycle[ 3673] = 1'b0;  wr_cycle[ 3673] = 1'b1;  addr_rom[ 3673]='h00003964;  wr_data_rom[ 3673]='h00000159;
    rd_cycle[ 3674] = 1'b0;  wr_cycle[ 3674] = 1'b1;  addr_rom[ 3674]='h00003968;  wr_data_rom[ 3674]='h00002887;
    rd_cycle[ 3675] = 1'b0;  wr_cycle[ 3675] = 1'b1;  addr_rom[ 3675]='h0000396c;  wr_data_rom[ 3675]='h000003c6;
    rd_cycle[ 3676] = 1'b0;  wr_cycle[ 3676] = 1'b1;  addr_rom[ 3676]='h00003970;  wr_data_rom[ 3676]='h00003b2d;
    rd_cycle[ 3677] = 1'b0;  wr_cycle[ 3677] = 1'b1;  addr_rom[ 3677]='h00003974;  wr_data_rom[ 3677]='h00002736;
    rd_cycle[ 3678] = 1'b0;  wr_cycle[ 3678] = 1'b1;  addr_rom[ 3678]='h00003978;  wr_data_rom[ 3678]='h00000f09;
    rd_cycle[ 3679] = 1'b0;  wr_cycle[ 3679] = 1'b1;  addr_rom[ 3679]='h0000397c;  wr_data_rom[ 3679]='h00003220;
    rd_cycle[ 3680] = 1'b0;  wr_cycle[ 3680] = 1'b1;  addr_rom[ 3680]='h00003980;  wr_data_rom[ 3680]='h00000a67;
    rd_cycle[ 3681] = 1'b0;  wr_cycle[ 3681] = 1'b1;  addr_rom[ 3681]='h00003984;  wr_data_rom[ 3681]='h0000000c;
    rd_cycle[ 3682] = 1'b0;  wr_cycle[ 3682] = 1'b1;  addr_rom[ 3682]='h00003988;  wr_data_rom[ 3682]='h0000061c;
    rd_cycle[ 3683] = 1'b0;  wr_cycle[ 3683] = 1'b1;  addr_rom[ 3683]='h0000398c;  wr_data_rom[ 3683]='h00003f17;
    rd_cycle[ 3684] = 1'b0;  wr_cycle[ 3684] = 1'b1;  addr_rom[ 3684]='h00003990;  wr_data_rom[ 3684]='h00003c35;
    rd_cycle[ 3685] = 1'b0;  wr_cycle[ 3685] = 1'b1;  addr_rom[ 3685]='h00003994;  wr_data_rom[ 3685]='h00002126;
    rd_cycle[ 3686] = 1'b0;  wr_cycle[ 3686] = 1'b1;  addr_rom[ 3686]='h00003998;  wr_data_rom[ 3686]='h0000393c;
    rd_cycle[ 3687] = 1'b0;  wr_cycle[ 3687] = 1'b1;  addr_rom[ 3687]='h0000399c;  wr_data_rom[ 3687]='h00001a23;
    rd_cycle[ 3688] = 1'b0;  wr_cycle[ 3688] = 1'b1;  addr_rom[ 3688]='h000039a0;  wr_data_rom[ 3688]='h00000ebe;
    rd_cycle[ 3689] = 1'b0;  wr_cycle[ 3689] = 1'b1;  addr_rom[ 3689]='h000039a4;  wr_data_rom[ 3689]='h00001e4c;
    rd_cycle[ 3690] = 1'b0;  wr_cycle[ 3690] = 1'b1;  addr_rom[ 3690]='h000039a8;  wr_data_rom[ 3690]='h0000154f;
    rd_cycle[ 3691] = 1'b0;  wr_cycle[ 3691] = 1'b1;  addr_rom[ 3691]='h000039ac;  wr_data_rom[ 3691]='h00003ba1;
    rd_cycle[ 3692] = 1'b0;  wr_cycle[ 3692] = 1'b1;  addr_rom[ 3692]='h000039b0;  wr_data_rom[ 3692]='h00001e05;
    rd_cycle[ 3693] = 1'b0;  wr_cycle[ 3693] = 1'b1;  addr_rom[ 3693]='h000039b4;  wr_data_rom[ 3693]='h0000161a;
    rd_cycle[ 3694] = 1'b0;  wr_cycle[ 3694] = 1'b1;  addr_rom[ 3694]='h000039b8;  wr_data_rom[ 3694]='h00000c64;
    rd_cycle[ 3695] = 1'b0;  wr_cycle[ 3695] = 1'b1;  addr_rom[ 3695]='h000039bc;  wr_data_rom[ 3695]='h00002f3b;
    rd_cycle[ 3696] = 1'b0;  wr_cycle[ 3696] = 1'b1;  addr_rom[ 3696]='h000039c0;  wr_data_rom[ 3696]='h00002452;
    rd_cycle[ 3697] = 1'b0;  wr_cycle[ 3697] = 1'b1;  addr_rom[ 3697]='h000039c4;  wr_data_rom[ 3697]='h00000dbd;
    rd_cycle[ 3698] = 1'b0;  wr_cycle[ 3698] = 1'b1;  addr_rom[ 3698]='h000039c8;  wr_data_rom[ 3698]='h00000d73;
    rd_cycle[ 3699] = 1'b0;  wr_cycle[ 3699] = 1'b1;  addr_rom[ 3699]='h000039cc;  wr_data_rom[ 3699]='h000026e6;
    rd_cycle[ 3700] = 1'b0;  wr_cycle[ 3700] = 1'b1;  addr_rom[ 3700]='h000039d0;  wr_data_rom[ 3700]='h0000078b;
    rd_cycle[ 3701] = 1'b0;  wr_cycle[ 3701] = 1'b1;  addr_rom[ 3701]='h000039d4;  wr_data_rom[ 3701]='h00003e9c;
    rd_cycle[ 3702] = 1'b0;  wr_cycle[ 3702] = 1'b1;  addr_rom[ 3702]='h000039d8;  wr_data_rom[ 3702]='h000003ce;
    rd_cycle[ 3703] = 1'b0;  wr_cycle[ 3703] = 1'b1;  addr_rom[ 3703]='h000039dc;  wr_data_rom[ 3703]='h00002d97;
    rd_cycle[ 3704] = 1'b0;  wr_cycle[ 3704] = 1'b1;  addr_rom[ 3704]='h000039e0;  wr_data_rom[ 3704]='h000025ae;
    rd_cycle[ 3705] = 1'b0;  wr_cycle[ 3705] = 1'b1;  addr_rom[ 3705]='h000039e4;  wr_data_rom[ 3705]='h00001c25;
    rd_cycle[ 3706] = 1'b0;  wr_cycle[ 3706] = 1'b1;  addr_rom[ 3706]='h000039e8;  wr_data_rom[ 3706]='h00000ab7;
    rd_cycle[ 3707] = 1'b0;  wr_cycle[ 3707] = 1'b1;  addr_rom[ 3707]='h000039ec;  wr_data_rom[ 3707]='h0000003f;
    rd_cycle[ 3708] = 1'b0;  wr_cycle[ 3708] = 1'b1;  addr_rom[ 3708]='h000039f0;  wr_data_rom[ 3708]='h00001c9b;
    rd_cycle[ 3709] = 1'b0;  wr_cycle[ 3709] = 1'b1;  addr_rom[ 3709]='h000039f4;  wr_data_rom[ 3709]='h000024ee;
    rd_cycle[ 3710] = 1'b0;  wr_cycle[ 3710] = 1'b1;  addr_rom[ 3710]='h000039f8;  wr_data_rom[ 3710]='h0000293a;
    rd_cycle[ 3711] = 1'b0;  wr_cycle[ 3711] = 1'b1;  addr_rom[ 3711]='h000039fc;  wr_data_rom[ 3711]='h000002f3;
    rd_cycle[ 3712] = 1'b0;  wr_cycle[ 3712] = 1'b1;  addr_rom[ 3712]='h00003a00;  wr_data_rom[ 3712]='h00001ed5;
    rd_cycle[ 3713] = 1'b0;  wr_cycle[ 3713] = 1'b1;  addr_rom[ 3713]='h00003a04;  wr_data_rom[ 3713]='h000007f7;
    rd_cycle[ 3714] = 1'b0;  wr_cycle[ 3714] = 1'b1;  addr_rom[ 3714]='h00003a08;  wr_data_rom[ 3714]='h00000d3f;
    rd_cycle[ 3715] = 1'b0;  wr_cycle[ 3715] = 1'b1;  addr_rom[ 3715]='h00003a0c;  wr_data_rom[ 3715]='h00000fff;
    rd_cycle[ 3716] = 1'b0;  wr_cycle[ 3716] = 1'b1;  addr_rom[ 3716]='h00003a10;  wr_data_rom[ 3716]='h00002a69;
    rd_cycle[ 3717] = 1'b0;  wr_cycle[ 3717] = 1'b1;  addr_rom[ 3717]='h00003a14;  wr_data_rom[ 3717]='h00003394;
    rd_cycle[ 3718] = 1'b0;  wr_cycle[ 3718] = 1'b1;  addr_rom[ 3718]='h00003a18;  wr_data_rom[ 3718]='h00002c1c;
    rd_cycle[ 3719] = 1'b0;  wr_cycle[ 3719] = 1'b1;  addr_rom[ 3719]='h00003a1c;  wr_data_rom[ 3719]='h000032c1;
    rd_cycle[ 3720] = 1'b0;  wr_cycle[ 3720] = 1'b1;  addr_rom[ 3720]='h00003a20;  wr_data_rom[ 3720]='h00001596;
    rd_cycle[ 3721] = 1'b0;  wr_cycle[ 3721] = 1'b1;  addr_rom[ 3721]='h00003a24;  wr_data_rom[ 3721]='h000034d6;
    rd_cycle[ 3722] = 1'b0;  wr_cycle[ 3722] = 1'b1;  addr_rom[ 3722]='h00003a28;  wr_data_rom[ 3722]='h00002ed9;
    rd_cycle[ 3723] = 1'b0;  wr_cycle[ 3723] = 1'b1;  addr_rom[ 3723]='h00003a2c;  wr_data_rom[ 3723]='h00002b1f;
    rd_cycle[ 3724] = 1'b0;  wr_cycle[ 3724] = 1'b1;  addr_rom[ 3724]='h00003a30;  wr_data_rom[ 3724]='h00002f54;
    rd_cycle[ 3725] = 1'b0;  wr_cycle[ 3725] = 1'b1;  addr_rom[ 3725]='h00003a34;  wr_data_rom[ 3725]='h00002eb7;
    rd_cycle[ 3726] = 1'b0;  wr_cycle[ 3726] = 1'b1;  addr_rom[ 3726]='h00003a38;  wr_data_rom[ 3726]='h00003b9b;
    rd_cycle[ 3727] = 1'b0;  wr_cycle[ 3727] = 1'b1;  addr_rom[ 3727]='h00003a3c;  wr_data_rom[ 3727]='h000007f2;
    rd_cycle[ 3728] = 1'b0;  wr_cycle[ 3728] = 1'b1;  addr_rom[ 3728]='h00003a40;  wr_data_rom[ 3728]='h00001d0c;
    rd_cycle[ 3729] = 1'b0;  wr_cycle[ 3729] = 1'b1;  addr_rom[ 3729]='h00003a44;  wr_data_rom[ 3729]='h00002913;
    rd_cycle[ 3730] = 1'b0;  wr_cycle[ 3730] = 1'b1;  addr_rom[ 3730]='h00003a48;  wr_data_rom[ 3730]='h00003bb9;
    rd_cycle[ 3731] = 1'b0;  wr_cycle[ 3731] = 1'b1;  addr_rom[ 3731]='h00003a4c;  wr_data_rom[ 3731]='h00000c25;
    rd_cycle[ 3732] = 1'b0;  wr_cycle[ 3732] = 1'b1;  addr_rom[ 3732]='h00003a50;  wr_data_rom[ 3732]='h00001552;
    rd_cycle[ 3733] = 1'b0;  wr_cycle[ 3733] = 1'b1;  addr_rom[ 3733]='h00003a54;  wr_data_rom[ 3733]='h00002f9a;
    rd_cycle[ 3734] = 1'b0;  wr_cycle[ 3734] = 1'b1;  addr_rom[ 3734]='h00003a58;  wr_data_rom[ 3734]='h00000aec;
    rd_cycle[ 3735] = 1'b0;  wr_cycle[ 3735] = 1'b1;  addr_rom[ 3735]='h00003a5c;  wr_data_rom[ 3735]='h00003474;
    rd_cycle[ 3736] = 1'b0;  wr_cycle[ 3736] = 1'b1;  addr_rom[ 3736]='h00003a60;  wr_data_rom[ 3736]='h0000345a;
    rd_cycle[ 3737] = 1'b0;  wr_cycle[ 3737] = 1'b1;  addr_rom[ 3737]='h00003a64;  wr_data_rom[ 3737]='h00003b4b;
    rd_cycle[ 3738] = 1'b0;  wr_cycle[ 3738] = 1'b1;  addr_rom[ 3738]='h00003a68;  wr_data_rom[ 3738]='h00003294;
    rd_cycle[ 3739] = 1'b0;  wr_cycle[ 3739] = 1'b1;  addr_rom[ 3739]='h00003a6c;  wr_data_rom[ 3739]='h000032e7;
    rd_cycle[ 3740] = 1'b0;  wr_cycle[ 3740] = 1'b1;  addr_rom[ 3740]='h00003a70;  wr_data_rom[ 3740]='h00002a15;
    rd_cycle[ 3741] = 1'b0;  wr_cycle[ 3741] = 1'b1;  addr_rom[ 3741]='h00003a74;  wr_data_rom[ 3741]='h000037f5;
    rd_cycle[ 3742] = 1'b0;  wr_cycle[ 3742] = 1'b1;  addr_rom[ 3742]='h00003a78;  wr_data_rom[ 3742]='h00002a67;
    rd_cycle[ 3743] = 1'b0;  wr_cycle[ 3743] = 1'b1;  addr_rom[ 3743]='h00003a7c;  wr_data_rom[ 3743]='h00002847;
    rd_cycle[ 3744] = 1'b0;  wr_cycle[ 3744] = 1'b1;  addr_rom[ 3744]='h00003a80;  wr_data_rom[ 3744]='h0000300a;
    rd_cycle[ 3745] = 1'b0;  wr_cycle[ 3745] = 1'b1;  addr_rom[ 3745]='h00003a84;  wr_data_rom[ 3745]='h00000d62;
    rd_cycle[ 3746] = 1'b0;  wr_cycle[ 3746] = 1'b1;  addr_rom[ 3746]='h00003a88;  wr_data_rom[ 3746]='h00002115;
    rd_cycle[ 3747] = 1'b0;  wr_cycle[ 3747] = 1'b1;  addr_rom[ 3747]='h00003a8c;  wr_data_rom[ 3747]='h00002f11;
    rd_cycle[ 3748] = 1'b0;  wr_cycle[ 3748] = 1'b1;  addr_rom[ 3748]='h00003a90;  wr_data_rom[ 3748]='h00000845;
    rd_cycle[ 3749] = 1'b0;  wr_cycle[ 3749] = 1'b1;  addr_rom[ 3749]='h00003a94;  wr_data_rom[ 3749]='h00000dae;
    rd_cycle[ 3750] = 1'b0;  wr_cycle[ 3750] = 1'b1;  addr_rom[ 3750]='h00003a98;  wr_data_rom[ 3750]='h00003846;
    rd_cycle[ 3751] = 1'b0;  wr_cycle[ 3751] = 1'b1;  addr_rom[ 3751]='h00003a9c;  wr_data_rom[ 3751]='h000027a2;
    rd_cycle[ 3752] = 1'b0;  wr_cycle[ 3752] = 1'b1;  addr_rom[ 3752]='h00003aa0;  wr_data_rom[ 3752]='h00000d91;
    rd_cycle[ 3753] = 1'b0;  wr_cycle[ 3753] = 1'b1;  addr_rom[ 3753]='h00003aa4;  wr_data_rom[ 3753]='h000019ff;
    rd_cycle[ 3754] = 1'b0;  wr_cycle[ 3754] = 1'b1;  addr_rom[ 3754]='h00003aa8;  wr_data_rom[ 3754]='h00001ebb;
    rd_cycle[ 3755] = 1'b0;  wr_cycle[ 3755] = 1'b1;  addr_rom[ 3755]='h00003aac;  wr_data_rom[ 3755]='h00003d5d;
    rd_cycle[ 3756] = 1'b0;  wr_cycle[ 3756] = 1'b1;  addr_rom[ 3756]='h00003ab0;  wr_data_rom[ 3756]='h00000742;
    rd_cycle[ 3757] = 1'b0;  wr_cycle[ 3757] = 1'b1;  addr_rom[ 3757]='h00003ab4;  wr_data_rom[ 3757]='h00000f63;
    rd_cycle[ 3758] = 1'b0;  wr_cycle[ 3758] = 1'b1;  addr_rom[ 3758]='h00003ab8;  wr_data_rom[ 3758]='h00002304;
    rd_cycle[ 3759] = 1'b0;  wr_cycle[ 3759] = 1'b1;  addr_rom[ 3759]='h00003abc;  wr_data_rom[ 3759]='h00001b85;
    rd_cycle[ 3760] = 1'b0;  wr_cycle[ 3760] = 1'b1;  addr_rom[ 3760]='h00003ac0;  wr_data_rom[ 3760]='h00001dac;
    rd_cycle[ 3761] = 1'b0;  wr_cycle[ 3761] = 1'b1;  addr_rom[ 3761]='h00003ac4;  wr_data_rom[ 3761]='h00002b10;
    rd_cycle[ 3762] = 1'b0;  wr_cycle[ 3762] = 1'b1;  addr_rom[ 3762]='h00003ac8;  wr_data_rom[ 3762]='h00001e0a;
    rd_cycle[ 3763] = 1'b0;  wr_cycle[ 3763] = 1'b1;  addr_rom[ 3763]='h00003acc;  wr_data_rom[ 3763]='h000016a5;
    rd_cycle[ 3764] = 1'b0;  wr_cycle[ 3764] = 1'b1;  addr_rom[ 3764]='h00003ad0;  wr_data_rom[ 3764]='h00002b1f;
    rd_cycle[ 3765] = 1'b0;  wr_cycle[ 3765] = 1'b1;  addr_rom[ 3765]='h00003ad4;  wr_data_rom[ 3765]='h00002769;
    rd_cycle[ 3766] = 1'b0;  wr_cycle[ 3766] = 1'b1;  addr_rom[ 3766]='h00003ad8;  wr_data_rom[ 3766]='h00001ae4;
    rd_cycle[ 3767] = 1'b0;  wr_cycle[ 3767] = 1'b1;  addr_rom[ 3767]='h00003adc;  wr_data_rom[ 3767]='h00002cce;
    rd_cycle[ 3768] = 1'b0;  wr_cycle[ 3768] = 1'b1;  addr_rom[ 3768]='h00003ae0;  wr_data_rom[ 3768]='h00002e8e;
    rd_cycle[ 3769] = 1'b0;  wr_cycle[ 3769] = 1'b1;  addr_rom[ 3769]='h00003ae4;  wr_data_rom[ 3769]='h000031fe;
    rd_cycle[ 3770] = 1'b0;  wr_cycle[ 3770] = 1'b1;  addr_rom[ 3770]='h00003ae8;  wr_data_rom[ 3770]='h00002b8e;
    rd_cycle[ 3771] = 1'b0;  wr_cycle[ 3771] = 1'b1;  addr_rom[ 3771]='h00003aec;  wr_data_rom[ 3771]='h00001514;
    rd_cycle[ 3772] = 1'b0;  wr_cycle[ 3772] = 1'b1;  addr_rom[ 3772]='h00003af0;  wr_data_rom[ 3772]='h00001f44;
    rd_cycle[ 3773] = 1'b0;  wr_cycle[ 3773] = 1'b1;  addr_rom[ 3773]='h00003af4;  wr_data_rom[ 3773]='h000001a3;
    rd_cycle[ 3774] = 1'b0;  wr_cycle[ 3774] = 1'b1;  addr_rom[ 3774]='h00003af8;  wr_data_rom[ 3774]='h00001dc6;
    rd_cycle[ 3775] = 1'b0;  wr_cycle[ 3775] = 1'b1;  addr_rom[ 3775]='h00003afc;  wr_data_rom[ 3775]='h00003f23;
    rd_cycle[ 3776] = 1'b0;  wr_cycle[ 3776] = 1'b1;  addr_rom[ 3776]='h00003b00;  wr_data_rom[ 3776]='h000000b3;
    rd_cycle[ 3777] = 1'b0;  wr_cycle[ 3777] = 1'b1;  addr_rom[ 3777]='h00003b04;  wr_data_rom[ 3777]='h00002890;
    rd_cycle[ 3778] = 1'b0;  wr_cycle[ 3778] = 1'b1;  addr_rom[ 3778]='h00003b08;  wr_data_rom[ 3778]='h00003b1b;
    rd_cycle[ 3779] = 1'b0;  wr_cycle[ 3779] = 1'b1;  addr_rom[ 3779]='h00003b0c;  wr_data_rom[ 3779]='h00003619;
    rd_cycle[ 3780] = 1'b0;  wr_cycle[ 3780] = 1'b1;  addr_rom[ 3780]='h00003b10;  wr_data_rom[ 3780]='h000000a5;
    rd_cycle[ 3781] = 1'b0;  wr_cycle[ 3781] = 1'b1;  addr_rom[ 3781]='h00003b14;  wr_data_rom[ 3781]='h000020c2;
    rd_cycle[ 3782] = 1'b0;  wr_cycle[ 3782] = 1'b1;  addr_rom[ 3782]='h00003b18;  wr_data_rom[ 3782]='h00001f23;
    rd_cycle[ 3783] = 1'b0;  wr_cycle[ 3783] = 1'b1;  addr_rom[ 3783]='h00003b1c;  wr_data_rom[ 3783]='h000013c8;
    rd_cycle[ 3784] = 1'b0;  wr_cycle[ 3784] = 1'b1;  addr_rom[ 3784]='h00003b20;  wr_data_rom[ 3784]='h000025dd;
    rd_cycle[ 3785] = 1'b0;  wr_cycle[ 3785] = 1'b1;  addr_rom[ 3785]='h00003b24;  wr_data_rom[ 3785]='h000032f8;
    rd_cycle[ 3786] = 1'b0;  wr_cycle[ 3786] = 1'b1;  addr_rom[ 3786]='h00003b28;  wr_data_rom[ 3786]='h0000343e;
    rd_cycle[ 3787] = 1'b0;  wr_cycle[ 3787] = 1'b1;  addr_rom[ 3787]='h00003b2c;  wr_data_rom[ 3787]='h00002c91;
    rd_cycle[ 3788] = 1'b0;  wr_cycle[ 3788] = 1'b1;  addr_rom[ 3788]='h00003b30;  wr_data_rom[ 3788]='h00002e7e;
    rd_cycle[ 3789] = 1'b0;  wr_cycle[ 3789] = 1'b1;  addr_rom[ 3789]='h00003b34;  wr_data_rom[ 3789]='h00000079;
    rd_cycle[ 3790] = 1'b0;  wr_cycle[ 3790] = 1'b1;  addr_rom[ 3790]='h00003b38;  wr_data_rom[ 3790]='h0000208f;
    rd_cycle[ 3791] = 1'b0;  wr_cycle[ 3791] = 1'b1;  addr_rom[ 3791]='h00003b3c;  wr_data_rom[ 3791]='h000038c9;
    rd_cycle[ 3792] = 1'b0;  wr_cycle[ 3792] = 1'b1;  addr_rom[ 3792]='h00003b40;  wr_data_rom[ 3792]='h00001ca5;
    rd_cycle[ 3793] = 1'b0;  wr_cycle[ 3793] = 1'b1;  addr_rom[ 3793]='h00003b44;  wr_data_rom[ 3793]='h00001875;
    rd_cycle[ 3794] = 1'b0;  wr_cycle[ 3794] = 1'b1;  addr_rom[ 3794]='h00003b48;  wr_data_rom[ 3794]='h00002bf2;
    rd_cycle[ 3795] = 1'b0;  wr_cycle[ 3795] = 1'b1;  addr_rom[ 3795]='h00003b4c;  wr_data_rom[ 3795]='h000007a6;
    rd_cycle[ 3796] = 1'b0;  wr_cycle[ 3796] = 1'b1;  addr_rom[ 3796]='h00003b50;  wr_data_rom[ 3796]='h00000fa5;
    rd_cycle[ 3797] = 1'b0;  wr_cycle[ 3797] = 1'b1;  addr_rom[ 3797]='h00003b54;  wr_data_rom[ 3797]='h00001301;
    rd_cycle[ 3798] = 1'b0;  wr_cycle[ 3798] = 1'b1;  addr_rom[ 3798]='h00003b58;  wr_data_rom[ 3798]='h00001cf5;
    rd_cycle[ 3799] = 1'b0;  wr_cycle[ 3799] = 1'b1;  addr_rom[ 3799]='h00003b5c;  wr_data_rom[ 3799]='h00000c34;
    rd_cycle[ 3800] = 1'b0;  wr_cycle[ 3800] = 1'b1;  addr_rom[ 3800]='h00003b60;  wr_data_rom[ 3800]='h000023f5;
    rd_cycle[ 3801] = 1'b0;  wr_cycle[ 3801] = 1'b1;  addr_rom[ 3801]='h00003b64;  wr_data_rom[ 3801]='h00001c6e;
    rd_cycle[ 3802] = 1'b0;  wr_cycle[ 3802] = 1'b1;  addr_rom[ 3802]='h00003b68;  wr_data_rom[ 3802]='h0000179e;
    rd_cycle[ 3803] = 1'b0;  wr_cycle[ 3803] = 1'b1;  addr_rom[ 3803]='h00003b6c;  wr_data_rom[ 3803]='h00001ac8;
    rd_cycle[ 3804] = 1'b0;  wr_cycle[ 3804] = 1'b1;  addr_rom[ 3804]='h00003b70;  wr_data_rom[ 3804]='h000010fc;
    rd_cycle[ 3805] = 1'b0;  wr_cycle[ 3805] = 1'b1;  addr_rom[ 3805]='h00003b74;  wr_data_rom[ 3805]='h00002038;
    rd_cycle[ 3806] = 1'b0;  wr_cycle[ 3806] = 1'b1;  addr_rom[ 3806]='h00003b78;  wr_data_rom[ 3806]='h0000389e;
    rd_cycle[ 3807] = 1'b0;  wr_cycle[ 3807] = 1'b1;  addr_rom[ 3807]='h00003b7c;  wr_data_rom[ 3807]='h00002ad6;
    rd_cycle[ 3808] = 1'b0;  wr_cycle[ 3808] = 1'b1;  addr_rom[ 3808]='h00003b80;  wr_data_rom[ 3808]='h000023f4;
    rd_cycle[ 3809] = 1'b0;  wr_cycle[ 3809] = 1'b1;  addr_rom[ 3809]='h00003b84;  wr_data_rom[ 3809]='h00002292;
    rd_cycle[ 3810] = 1'b0;  wr_cycle[ 3810] = 1'b1;  addr_rom[ 3810]='h00003b88;  wr_data_rom[ 3810]='h00001582;
    rd_cycle[ 3811] = 1'b0;  wr_cycle[ 3811] = 1'b1;  addr_rom[ 3811]='h00003b8c;  wr_data_rom[ 3811]='h00003eb2;
    rd_cycle[ 3812] = 1'b0;  wr_cycle[ 3812] = 1'b1;  addr_rom[ 3812]='h00003b90;  wr_data_rom[ 3812]='h000006a0;
    rd_cycle[ 3813] = 1'b0;  wr_cycle[ 3813] = 1'b1;  addr_rom[ 3813]='h00003b94;  wr_data_rom[ 3813]='h0000206d;
    rd_cycle[ 3814] = 1'b0;  wr_cycle[ 3814] = 1'b1;  addr_rom[ 3814]='h00003b98;  wr_data_rom[ 3814]='h000039a7;
    rd_cycle[ 3815] = 1'b0;  wr_cycle[ 3815] = 1'b1;  addr_rom[ 3815]='h00003b9c;  wr_data_rom[ 3815]='h00002f15;
    rd_cycle[ 3816] = 1'b0;  wr_cycle[ 3816] = 1'b1;  addr_rom[ 3816]='h00003ba0;  wr_data_rom[ 3816]='h000036e2;
    rd_cycle[ 3817] = 1'b0;  wr_cycle[ 3817] = 1'b1;  addr_rom[ 3817]='h00003ba4;  wr_data_rom[ 3817]='h00001694;
    rd_cycle[ 3818] = 1'b0;  wr_cycle[ 3818] = 1'b1;  addr_rom[ 3818]='h00003ba8;  wr_data_rom[ 3818]='h00001935;
    rd_cycle[ 3819] = 1'b0;  wr_cycle[ 3819] = 1'b1;  addr_rom[ 3819]='h00003bac;  wr_data_rom[ 3819]='h00003fc9;
    rd_cycle[ 3820] = 1'b0;  wr_cycle[ 3820] = 1'b1;  addr_rom[ 3820]='h00003bb0;  wr_data_rom[ 3820]='h00003512;
    rd_cycle[ 3821] = 1'b0;  wr_cycle[ 3821] = 1'b1;  addr_rom[ 3821]='h00003bb4;  wr_data_rom[ 3821]='h00001e5f;
    rd_cycle[ 3822] = 1'b0;  wr_cycle[ 3822] = 1'b1;  addr_rom[ 3822]='h00003bb8;  wr_data_rom[ 3822]='h00003fa0;
    rd_cycle[ 3823] = 1'b0;  wr_cycle[ 3823] = 1'b1;  addr_rom[ 3823]='h00003bbc;  wr_data_rom[ 3823]='h00001a62;
    rd_cycle[ 3824] = 1'b0;  wr_cycle[ 3824] = 1'b1;  addr_rom[ 3824]='h00003bc0;  wr_data_rom[ 3824]='h0000022a;
    rd_cycle[ 3825] = 1'b0;  wr_cycle[ 3825] = 1'b1;  addr_rom[ 3825]='h00003bc4;  wr_data_rom[ 3825]='h000030af;
    rd_cycle[ 3826] = 1'b0;  wr_cycle[ 3826] = 1'b1;  addr_rom[ 3826]='h00003bc8;  wr_data_rom[ 3826]='h00000f3b;
    rd_cycle[ 3827] = 1'b0;  wr_cycle[ 3827] = 1'b1;  addr_rom[ 3827]='h00003bcc;  wr_data_rom[ 3827]='h0000292f;
    rd_cycle[ 3828] = 1'b0;  wr_cycle[ 3828] = 1'b1;  addr_rom[ 3828]='h00003bd0;  wr_data_rom[ 3828]='h000021b4;
    rd_cycle[ 3829] = 1'b0;  wr_cycle[ 3829] = 1'b1;  addr_rom[ 3829]='h00003bd4;  wr_data_rom[ 3829]='h00002ba8;
    rd_cycle[ 3830] = 1'b0;  wr_cycle[ 3830] = 1'b1;  addr_rom[ 3830]='h00003bd8;  wr_data_rom[ 3830]='h00001479;
    rd_cycle[ 3831] = 1'b0;  wr_cycle[ 3831] = 1'b1;  addr_rom[ 3831]='h00003bdc;  wr_data_rom[ 3831]='h00001155;
    rd_cycle[ 3832] = 1'b0;  wr_cycle[ 3832] = 1'b1;  addr_rom[ 3832]='h00003be0;  wr_data_rom[ 3832]='h00001607;
    rd_cycle[ 3833] = 1'b0;  wr_cycle[ 3833] = 1'b1;  addr_rom[ 3833]='h00003be4;  wr_data_rom[ 3833]='h0000296a;
    rd_cycle[ 3834] = 1'b0;  wr_cycle[ 3834] = 1'b1;  addr_rom[ 3834]='h00003be8;  wr_data_rom[ 3834]='h00001d65;
    rd_cycle[ 3835] = 1'b0;  wr_cycle[ 3835] = 1'b1;  addr_rom[ 3835]='h00003bec;  wr_data_rom[ 3835]='h00003fd9;
    rd_cycle[ 3836] = 1'b0;  wr_cycle[ 3836] = 1'b1;  addr_rom[ 3836]='h00003bf0;  wr_data_rom[ 3836]='h00003ca1;
    rd_cycle[ 3837] = 1'b0;  wr_cycle[ 3837] = 1'b1;  addr_rom[ 3837]='h00003bf4;  wr_data_rom[ 3837]='h00002918;
    rd_cycle[ 3838] = 1'b0;  wr_cycle[ 3838] = 1'b1;  addr_rom[ 3838]='h00003bf8;  wr_data_rom[ 3838]='h00002870;
    rd_cycle[ 3839] = 1'b0;  wr_cycle[ 3839] = 1'b1;  addr_rom[ 3839]='h00003bfc;  wr_data_rom[ 3839]='h0000188b;
    rd_cycle[ 3840] = 1'b0;  wr_cycle[ 3840] = 1'b1;  addr_rom[ 3840]='h00003c00;  wr_data_rom[ 3840]='h00001b83;
    rd_cycle[ 3841] = 1'b0;  wr_cycle[ 3841] = 1'b1;  addr_rom[ 3841]='h00003c04;  wr_data_rom[ 3841]='h00002967;
    rd_cycle[ 3842] = 1'b0;  wr_cycle[ 3842] = 1'b1;  addr_rom[ 3842]='h00003c08;  wr_data_rom[ 3842]='h00003a93;
    rd_cycle[ 3843] = 1'b0;  wr_cycle[ 3843] = 1'b1;  addr_rom[ 3843]='h00003c0c;  wr_data_rom[ 3843]='h000012cc;
    rd_cycle[ 3844] = 1'b0;  wr_cycle[ 3844] = 1'b1;  addr_rom[ 3844]='h00003c10;  wr_data_rom[ 3844]='h000010ae;
    rd_cycle[ 3845] = 1'b0;  wr_cycle[ 3845] = 1'b1;  addr_rom[ 3845]='h00003c14;  wr_data_rom[ 3845]='h00000a08;
    rd_cycle[ 3846] = 1'b0;  wr_cycle[ 3846] = 1'b1;  addr_rom[ 3846]='h00003c18;  wr_data_rom[ 3846]='h00002ab8;
    rd_cycle[ 3847] = 1'b0;  wr_cycle[ 3847] = 1'b1;  addr_rom[ 3847]='h00003c1c;  wr_data_rom[ 3847]='h00003ddf;
    rd_cycle[ 3848] = 1'b0;  wr_cycle[ 3848] = 1'b1;  addr_rom[ 3848]='h00003c20;  wr_data_rom[ 3848]='h00003f9b;
    rd_cycle[ 3849] = 1'b0;  wr_cycle[ 3849] = 1'b1;  addr_rom[ 3849]='h00003c24;  wr_data_rom[ 3849]='h00001b6e;
    rd_cycle[ 3850] = 1'b0;  wr_cycle[ 3850] = 1'b1;  addr_rom[ 3850]='h00003c28;  wr_data_rom[ 3850]='h000009cf;
    rd_cycle[ 3851] = 1'b0;  wr_cycle[ 3851] = 1'b1;  addr_rom[ 3851]='h00003c2c;  wr_data_rom[ 3851]='h00003209;
    rd_cycle[ 3852] = 1'b0;  wr_cycle[ 3852] = 1'b1;  addr_rom[ 3852]='h00003c30;  wr_data_rom[ 3852]='h000011b6;
    rd_cycle[ 3853] = 1'b0;  wr_cycle[ 3853] = 1'b1;  addr_rom[ 3853]='h00003c34;  wr_data_rom[ 3853]='h00002a3e;
    rd_cycle[ 3854] = 1'b0;  wr_cycle[ 3854] = 1'b1;  addr_rom[ 3854]='h00003c38;  wr_data_rom[ 3854]='h00003c59;
    rd_cycle[ 3855] = 1'b0;  wr_cycle[ 3855] = 1'b1;  addr_rom[ 3855]='h00003c3c;  wr_data_rom[ 3855]='h000014c0;
    rd_cycle[ 3856] = 1'b0;  wr_cycle[ 3856] = 1'b1;  addr_rom[ 3856]='h00003c40;  wr_data_rom[ 3856]='h000006c7;
    rd_cycle[ 3857] = 1'b0;  wr_cycle[ 3857] = 1'b1;  addr_rom[ 3857]='h00003c44;  wr_data_rom[ 3857]='h00001551;
    rd_cycle[ 3858] = 1'b0;  wr_cycle[ 3858] = 1'b1;  addr_rom[ 3858]='h00003c48;  wr_data_rom[ 3858]='h0000077a;
    rd_cycle[ 3859] = 1'b0;  wr_cycle[ 3859] = 1'b1;  addr_rom[ 3859]='h00003c4c;  wr_data_rom[ 3859]='h00002f6c;
    rd_cycle[ 3860] = 1'b0;  wr_cycle[ 3860] = 1'b1;  addr_rom[ 3860]='h00003c50;  wr_data_rom[ 3860]='h00003f62;
    rd_cycle[ 3861] = 1'b0;  wr_cycle[ 3861] = 1'b1;  addr_rom[ 3861]='h00003c54;  wr_data_rom[ 3861]='h000028b2;
    rd_cycle[ 3862] = 1'b0;  wr_cycle[ 3862] = 1'b1;  addr_rom[ 3862]='h00003c58;  wr_data_rom[ 3862]='h0000345c;
    rd_cycle[ 3863] = 1'b0;  wr_cycle[ 3863] = 1'b1;  addr_rom[ 3863]='h00003c5c;  wr_data_rom[ 3863]='h00000312;
    rd_cycle[ 3864] = 1'b0;  wr_cycle[ 3864] = 1'b1;  addr_rom[ 3864]='h00003c60;  wr_data_rom[ 3864]='h00001404;
    rd_cycle[ 3865] = 1'b0;  wr_cycle[ 3865] = 1'b1;  addr_rom[ 3865]='h00003c64;  wr_data_rom[ 3865]='h00002ef6;
    rd_cycle[ 3866] = 1'b0;  wr_cycle[ 3866] = 1'b1;  addr_rom[ 3866]='h00003c68;  wr_data_rom[ 3866]='h0000082f;
    rd_cycle[ 3867] = 1'b0;  wr_cycle[ 3867] = 1'b1;  addr_rom[ 3867]='h00003c6c;  wr_data_rom[ 3867]='h00000a21;
    rd_cycle[ 3868] = 1'b0;  wr_cycle[ 3868] = 1'b1;  addr_rom[ 3868]='h00003c70;  wr_data_rom[ 3868]='h00000117;
    rd_cycle[ 3869] = 1'b0;  wr_cycle[ 3869] = 1'b1;  addr_rom[ 3869]='h00003c74;  wr_data_rom[ 3869]='h00003e6b;
    rd_cycle[ 3870] = 1'b0;  wr_cycle[ 3870] = 1'b1;  addr_rom[ 3870]='h00003c78;  wr_data_rom[ 3870]='h000016ba;
    rd_cycle[ 3871] = 1'b0;  wr_cycle[ 3871] = 1'b1;  addr_rom[ 3871]='h00003c7c;  wr_data_rom[ 3871]='h00001313;
    rd_cycle[ 3872] = 1'b0;  wr_cycle[ 3872] = 1'b1;  addr_rom[ 3872]='h00003c80;  wr_data_rom[ 3872]='h0000367c;
    rd_cycle[ 3873] = 1'b0;  wr_cycle[ 3873] = 1'b1;  addr_rom[ 3873]='h00003c84;  wr_data_rom[ 3873]='h00002a43;
    rd_cycle[ 3874] = 1'b0;  wr_cycle[ 3874] = 1'b1;  addr_rom[ 3874]='h00003c88;  wr_data_rom[ 3874]='h00002672;
    rd_cycle[ 3875] = 1'b0;  wr_cycle[ 3875] = 1'b1;  addr_rom[ 3875]='h00003c8c;  wr_data_rom[ 3875]='h0000061c;
    rd_cycle[ 3876] = 1'b0;  wr_cycle[ 3876] = 1'b1;  addr_rom[ 3876]='h00003c90;  wr_data_rom[ 3876]='h00003d18;
    rd_cycle[ 3877] = 1'b0;  wr_cycle[ 3877] = 1'b1;  addr_rom[ 3877]='h00003c94;  wr_data_rom[ 3877]='h000009e7;
    rd_cycle[ 3878] = 1'b0;  wr_cycle[ 3878] = 1'b1;  addr_rom[ 3878]='h00003c98;  wr_data_rom[ 3878]='h00003d72;
    rd_cycle[ 3879] = 1'b0;  wr_cycle[ 3879] = 1'b1;  addr_rom[ 3879]='h00003c9c;  wr_data_rom[ 3879]='h00000fda;
    rd_cycle[ 3880] = 1'b0;  wr_cycle[ 3880] = 1'b1;  addr_rom[ 3880]='h00003ca0;  wr_data_rom[ 3880]='h00000f2f;
    rd_cycle[ 3881] = 1'b0;  wr_cycle[ 3881] = 1'b1;  addr_rom[ 3881]='h00003ca4;  wr_data_rom[ 3881]='h000022be;
    rd_cycle[ 3882] = 1'b0;  wr_cycle[ 3882] = 1'b1;  addr_rom[ 3882]='h00003ca8;  wr_data_rom[ 3882]='h00002646;
    rd_cycle[ 3883] = 1'b0;  wr_cycle[ 3883] = 1'b1;  addr_rom[ 3883]='h00003cac;  wr_data_rom[ 3883]='h00001b1c;
    rd_cycle[ 3884] = 1'b0;  wr_cycle[ 3884] = 1'b1;  addr_rom[ 3884]='h00003cb0;  wr_data_rom[ 3884]='h00003b6d;
    rd_cycle[ 3885] = 1'b0;  wr_cycle[ 3885] = 1'b1;  addr_rom[ 3885]='h00003cb4;  wr_data_rom[ 3885]='h00003a09;
    rd_cycle[ 3886] = 1'b0;  wr_cycle[ 3886] = 1'b1;  addr_rom[ 3886]='h00003cb8;  wr_data_rom[ 3886]='h000038ec;
    rd_cycle[ 3887] = 1'b0;  wr_cycle[ 3887] = 1'b1;  addr_rom[ 3887]='h00003cbc;  wr_data_rom[ 3887]='h00003c7c;
    rd_cycle[ 3888] = 1'b0;  wr_cycle[ 3888] = 1'b1;  addr_rom[ 3888]='h00003cc0;  wr_data_rom[ 3888]='h00000a40;
    rd_cycle[ 3889] = 1'b0;  wr_cycle[ 3889] = 1'b1;  addr_rom[ 3889]='h00003cc4;  wr_data_rom[ 3889]='h00003111;
    rd_cycle[ 3890] = 1'b0;  wr_cycle[ 3890] = 1'b1;  addr_rom[ 3890]='h00003cc8;  wr_data_rom[ 3890]='h00001a2a;
    rd_cycle[ 3891] = 1'b0;  wr_cycle[ 3891] = 1'b1;  addr_rom[ 3891]='h00003ccc;  wr_data_rom[ 3891]='h00000d70;
    rd_cycle[ 3892] = 1'b0;  wr_cycle[ 3892] = 1'b1;  addr_rom[ 3892]='h00003cd0;  wr_data_rom[ 3892]='h00000661;
    rd_cycle[ 3893] = 1'b0;  wr_cycle[ 3893] = 1'b1;  addr_rom[ 3893]='h00003cd4;  wr_data_rom[ 3893]='h000027b6;
    rd_cycle[ 3894] = 1'b0;  wr_cycle[ 3894] = 1'b1;  addr_rom[ 3894]='h00003cd8;  wr_data_rom[ 3894]='h00000e9b;
    rd_cycle[ 3895] = 1'b0;  wr_cycle[ 3895] = 1'b1;  addr_rom[ 3895]='h00003cdc;  wr_data_rom[ 3895]='h000020e1;
    rd_cycle[ 3896] = 1'b0;  wr_cycle[ 3896] = 1'b1;  addr_rom[ 3896]='h00003ce0;  wr_data_rom[ 3896]='h00000694;
    rd_cycle[ 3897] = 1'b0;  wr_cycle[ 3897] = 1'b1;  addr_rom[ 3897]='h00003ce4;  wr_data_rom[ 3897]='h000028a2;
    rd_cycle[ 3898] = 1'b0;  wr_cycle[ 3898] = 1'b1;  addr_rom[ 3898]='h00003ce8;  wr_data_rom[ 3898]='h00000ed9;
    rd_cycle[ 3899] = 1'b0;  wr_cycle[ 3899] = 1'b1;  addr_rom[ 3899]='h00003cec;  wr_data_rom[ 3899]='h0000322d;
    rd_cycle[ 3900] = 1'b0;  wr_cycle[ 3900] = 1'b1;  addr_rom[ 3900]='h00003cf0;  wr_data_rom[ 3900]='h000009cc;
    rd_cycle[ 3901] = 1'b0;  wr_cycle[ 3901] = 1'b1;  addr_rom[ 3901]='h00003cf4;  wr_data_rom[ 3901]='h00000e06;
    rd_cycle[ 3902] = 1'b0;  wr_cycle[ 3902] = 1'b1;  addr_rom[ 3902]='h00003cf8;  wr_data_rom[ 3902]='h000004c1;
    rd_cycle[ 3903] = 1'b0;  wr_cycle[ 3903] = 1'b1;  addr_rom[ 3903]='h00003cfc;  wr_data_rom[ 3903]='h00003643;
    rd_cycle[ 3904] = 1'b0;  wr_cycle[ 3904] = 1'b1;  addr_rom[ 3904]='h00003d00;  wr_data_rom[ 3904]='h00002ae9;
    rd_cycle[ 3905] = 1'b0;  wr_cycle[ 3905] = 1'b1;  addr_rom[ 3905]='h00003d04;  wr_data_rom[ 3905]='h00000ac3;
    rd_cycle[ 3906] = 1'b0;  wr_cycle[ 3906] = 1'b1;  addr_rom[ 3906]='h00003d08;  wr_data_rom[ 3906]='h00000bf8;
    rd_cycle[ 3907] = 1'b0;  wr_cycle[ 3907] = 1'b1;  addr_rom[ 3907]='h00003d0c;  wr_data_rom[ 3907]='h00000ba7;
    rd_cycle[ 3908] = 1'b0;  wr_cycle[ 3908] = 1'b1;  addr_rom[ 3908]='h00003d10;  wr_data_rom[ 3908]='h00000995;
    rd_cycle[ 3909] = 1'b0;  wr_cycle[ 3909] = 1'b1;  addr_rom[ 3909]='h00003d14;  wr_data_rom[ 3909]='h000032a5;
    rd_cycle[ 3910] = 1'b0;  wr_cycle[ 3910] = 1'b1;  addr_rom[ 3910]='h00003d18;  wr_data_rom[ 3910]='h000020fd;
    rd_cycle[ 3911] = 1'b0;  wr_cycle[ 3911] = 1'b1;  addr_rom[ 3911]='h00003d1c;  wr_data_rom[ 3911]='h00000730;
    rd_cycle[ 3912] = 1'b0;  wr_cycle[ 3912] = 1'b1;  addr_rom[ 3912]='h00003d20;  wr_data_rom[ 3912]='h00003fbf;
    rd_cycle[ 3913] = 1'b0;  wr_cycle[ 3913] = 1'b1;  addr_rom[ 3913]='h00003d24;  wr_data_rom[ 3913]='h00001e98;
    rd_cycle[ 3914] = 1'b0;  wr_cycle[ 3914] = 1'b1;  addr_rom[ 3914]='h00003d28;  wr_data_rom[ 3914]='h00002f4a;
    rd_cycle[ 3915] = 1'b0;  wr_cycle[ 3915] = 1'b1;  addr_rom[ 3915]='h00003d2c;  wr_data_rom[ 3915]='h00001375;
    rd_cycle[ 3916] = 1'b0;  wr_cycle[ 3916] = 1'b1;  addr_rom[ 3916]='h00003d30;  wr_data_rom[ 3916]='h000038dd;
    rd_cycle[ 3917] = 1'b0;  wr_cycle[ 3917] = 1'b1;  addr_rom[ 3917]='h00003d34;  wr_data_rom[ 3917]='h00003b7e;
    rd_cycle[ 3918] = 1'b0;  wr_cycle[ 3918] = 1'b1;  addr_rom[ 3918]='h00003d38;  wr_data_rom[ 3918]='h000006f0;
    rd_cycle[ 3919] = 1'b0;  wr_cycle[ 3919] = 1'b1;  addr_rom[ 3919]='h00003d3c;  wr_data_rom[ 3919]='h000027b6;
    rd_cycle[ 3920] = 1'b0;  wr_cycle[ 3920] = 1'b1;  addr_rom[ 3920]='h00003d40;  wr_data_rom[ 3920]='h00001e9c;
    rd_cycle[ 3921] = 1'b0;  wr_cycle[ 3921] = 1'b1;  addr_rom[ 3921]='h00003d44;  wr_data_rom[ 3921]='h000020c0;
    rd_cycle[ 3922] = 1'b0;  wr_cycle[ 3922] = 1'b1;  addr_rom[ 3922]='h00003d48;  wr_data_rom[ 3922]='h0000183d;
    rd_cycle[ 3923] = 1'b0;  wr_cycle[ 3923] = 1'b1;  addr_rom[ 3923]='h00003d4c;  wr_data_rom[ 3923]='h00001c5e;
    rd_cycle[ 3924] = 1'b0;  wr_cycle[ 3924] = 1'b1;  addr_rom[ 3924]='h00003d50;  wr_data_rom[ 3924]='h0000162e;
    rd_cycle[ 3925] = 1'b0;  wr_cycle[ 3925] = 1'b1;  addr_rom[ 3925]='h00003d54;  wr_data_rom[ 3925]='h00000cdc;
    rd_cycle[ 3926] = 1'b0;  wr_cycle[ 3926] = 1'b1;  addr_rom[ 3926]='h00003d58;  wr_data_rom[ 3926]='h000038a8;
    rd_cycle[ 3927] = 1'b0;  wr_cycle[ 3927] = 1'b1;  addr_rom[ 3927]='h00003d5c;  wr_data_rom[ 3927]='h000038ab;
    rd_cycle[ 3928] = 1'b0;  wr_cycle[ 3928] = 1'b1;  addr_rom[ 3928]='h00003d60;  wr_data_rom[ 3928]='h00002b78;
    rd_cycle[ 3929] = 1'b0;  wr_cycle[ 3929] = 1'b1;  addr_rom[ 3929]='h00003d64;  wr_data_rom[ 3929]='h000026bc;
    rd_cycle[ 3930] = 1'b0;  wr_cycle[ 3930] = 1'b1;  addr_rom[ 3930]='h00003d68;  wr_data_rom[ 3930]='h00003550;
    rd_cycle[ 3931] = 1'b0;  wr_cycle[ 3931] = 1'b1;  addr_rom[ 3931]='h00003d6c;  wr_data_rom[ 3931]='h0000387f;
    rd_cycle[ 3932] = 1'b0;  wr_cycle[ 3932] = 1'b1;  addr_rom[ 3932]='h00003d70;  wr_data_rom[ 3932]='h00002024;
    rd_cycle[ 3933] = 1'b0;  wr_cycle[ 3933] = 1'b1;  addr_rom[ 3933]='h00003d74;  wr_data_rom[ 3933]='h00000420;
    rd_cycle[ 3934] = 1'b0;  wr_cycle[ 3934] = 1'b1;  addr_rom[ 3934]='h00003d78;  wr_data_rom[ 3934]='h00001d50;
    rd_cycle[ 3935] = 1'b0;  wr_cycle[ 3935] = 1'b1;  addr_rom[ 3935]='h00003d7c;  wr_data_rom[ 3935]='h00000539;
    rd_cycle[ 3936] = 1'b0;  wr_cycle[ 3936] = 1'b1;  addr_rom[ 3936]='h00003d80;  wr_data_rom[ 3936]='h00002dd5;
    rd_cycle[ 3937] = 1'b0;  wr_cycle[ 3937] = 1'b1;  addr_rom[ 3937]='h00003d84;  wr_data_rom[ 3937]='h00000464;
    rd_cycle[ 3938] = 1'b0;  wr_cycle[ 3938] = 1'b1;  addr_rom[ 3938]='h00003d88;  wr_data_rom[ 3938]='h0000368a;
    rd_cycle[ 3939] = 1'b0;  wr_cycle[ 3939] = 1'b1;  addr_rom[ 3939]='h00003d8c;  wr_data_rom[ 3939]='h00003797;
    rd_cycle[ 3940] = 1'b0;  wr_cycle[ 3940] = 1'b1;  addr_rom[ 3940]='h00003d90;  wr_data_rom[ 3940]='h000030c2;
    rd_cycle[ 3941] = 1'b0;  wr_cycle[ 3941] = 1'b1;  addr_rom[ 3941]='h00003d94;  wr_data_rom[ 3941]='h0000257c;
    rd_cycle[ 3942] = 1'b0;  wr_cycle[ 3942] = 1'b1;  addr_rom[ 3942]='h00003d98;  wr_data_rom[ 3942]='h0000041a;
    rd_cycle[ 3943] = 1'b0;  wr_cycle[ 3943] = 1'b1;  addr_rom[ 3943]='h00003d9c;  wr_data_rom[ 3943]='h00001171;
    rd_cycle[ 3944] = 1'b0;  wr_cycle[ 3944] = 1'b1;  addr_rom[ 3944]='h00003da0;  wr_data_rom[ 3944]='h00002983;
    rd_cycle[ 3945] = 1'b0;  wr_cycle[ 3945] = 1'b1;  addr_rom[ 3945]='h00003da4;  wr_data_rom[ 3945]='h00002416;
    rd_cycle[ 3946] = 1'b0;  wr_cycle[ 3946] = 1'b1;  addr_rom[ 3946]='h00003da8;  wr_data_rom[ 3946]='h00001219;
    rd_cycle[ 3947] = 1'b0;  wr_cycle[ 3947] = 1'b1;  addr_rom[ 3947]='h00003dac;  wr_data_rom[ 3947]='h0000228a;
    rd_cycle[ 3948] = 1'b0;  wr_cycle[ 3948] = 1'b1;  addr_rom[ 3948]='h00003db0;  wr_data_rom[ 3948]='h000008f4;
    rd_cycle[ 3949] = 1'b0;  wr_cycle[ 3949] = 1'b1;  addr_rom[ 3949]='h00003db4;  wr_data_rom[ 3949]='h0000114c;
    rd_cycle[ 3950] = 1'b0;  wr_cycle[ 3950] = 1'b1;  addr_rom[ 3950]='h00003db8;  wr_data_rom[ 3950]='h0000022f;
    rd_cycle[ 3951] = 1'b0;  wr_cycle[ 3951] = 1'b1;  addr_rom[ 3951]='h00003dbc;  wr_data_rom[ 3951]='h00001136;
    rd_cycle[ 3952] = 1'b0;  wr_cycle[ 3952] = 1'b1;  addr_rom[ 3952]='h00003dc0;  wr_data_rom[ 3952]='h0000217d;
    rd_cycle[ 3953] = 1'b0;  wr_cycle[ 3953] = 1'b1;  addr_rom[ 3953]='h00003dc4;  wr_data_rom[ 3953]='h00003abf;
    rd_cycle[ 3954] = 1'b0;  wr_cycle[ 3954] = 1'b1;  addr_rom[ 3954]='h00003dc8;  wr_data_rom[ 3954]='h0000143a;
    rd_cycle[ 3955] = 1'b0;  wr_cycle[ 3955] = 1'b1;  addr_rom[ 3955]='h00003dcc;  wr_data_rom[ 3955]='h00003905;
    rd_cycle[ 3956] = 1'b0;  wr_cycle[ 3956] = 1'b1;  addr_rom[ 3956]='h00003dd0;  wr_data_rom[ 3956]='h0000128f;
    rd_cycle[ 3957] = 1'b0;  wr_cycle[ 3957] = 1'b1;  addr_rom[ 3957]='h00003dd4;  wr_data_rom[ 3957]='h000012f0;
    rd_cycle[ 3958] = 1'b0;  wr_cycle[ 3958] = 1'b1;  addr_rom[ 3958]='h00003dd8;  wr_data_rom[ 3958]='h0000098e;
    rd_cycle[ 3959] = 1'b0;  wr_cycle[ 3959] = 1'b1;  addr_rom[ 3959]='h00003ddc;  wr_data_rom[ 3959]='h00000d1c;
    rd_cycle[ 3960] = 1'b0;  wr_cycle[ 3960] = 1'b1;  addr_rom[ 3960]='h00003de0;  wr_data_rom[ 3960]='h00001c25;
    rd_cycle[ 3961] = 1'b0;  wr_cycle[ 3961] = 1'b1;  addr_rom[ 3961]='h00003de4;  wr_data_rom[ 3961]='h00000318;
    rd_cycle[ 3962] = 1'b0;  wr_cycle[ 3962] = 1'b1;  addr_rom[ 3962]='h00003de8;  wr_data_rom[ 3962]='h000024c7;
    rd_cycle[ 3963] = 1'b0;  wr_cycle[ 3963] = 1'b1;  addr_rom[ 3963]='h00003dec;  wr_data_rom[ 3963]='h000013bd;
    rd_cycle[ 3964] = 1'b0;  wr_cycle[ 3964] = 1'b1;  addr_rom[ 3964]='h00003df0;  wr_data_rom[ 3964]='h00003a63;
    rd_cycle[ 3965] = 1'b0;  wr_cycle[ 3965] = 1'b1;  addr_rom[ 3965]='h00003df4;  wr_data_rom[ 3965]='h00000a5c;
    rd_cycle[ 3966] = 1'b0;  wr_cycle[ 3966] = 1'b1;  addr_rom[ 3966]='h00003df8;  wr_data_rom[ 3966]='h00000733;
    rd_cycle[ 3967] = 1'b0;  wr_cycle[ 3967] = 1'b1;  addr_rom[ 3967]='h00003dfc;  wr_data_rom[ 3967]='h000000e2;
    rd_cycle[ 3968] = 1'b0;  wr_cycle[ 3968] = 1'b1;  addr_rom[ 3968]='h00003e00;  wr_data_rom[ 3968]='h00000331;
    rd_cycle[ 3969] = 1'b0;  wr_cycle[ 3969] = 1'b1;  addr_rom[ 3969]='h00003e04;  wr_data_rom[ 3969]='h00002bcc;
    rd_cycle[ 3970] = 1'b0;  wr_cycle[ 3970] = 1'b1;  addr_rom[ 3970]='h00003e08;  wr_data_rom[ 3970]='h00001ae1;
    rd_cycle[ 3971] = 1'b0;  wr_cycle[ 3971] = 1'b1;  addr_rom[ 3971]='h00003e0c;  wr_data_rom[ 3971]='h000015ff;
    rd_cycle[ 3972] = 1'b0;  wr_cycle[ 3972] = 1'b1;  addr_rom[ 3972]='h00003e10;  wr_data_rom[ 3972]='h000021d2;
    rd_cycle[ 3973] = 1'b0;  wr_cycle[ 3973] = 1'b1;  addr_rom[ 3973]='h00003e14;  wr_data_rom[ 3973]='h00003a57;
    rd_cycle[ 3974] = 1'b0;  wr_cycle[ 3974] = 1'b1;  addr_rom[ 3974]='h00003e18;  wr_data_rom[ 3974]='h00003412;
    rd_cycle[ 3975] = 1'b0;  wr_cycle[ 3975] = 1'b1;  addr_rom[ 3975]='h00003e1c;  wr_data_rom[ 3975]='h00000780;
    rd_cycle[ 3976] = 1'b0;  wr_cycle[ 3976] = 1'b1;  addr_rom[ 3976]='h00003e20;  wr_data_rom[ 3976]='h00003fba;
    rd_cycle[ 3977] = 1'b0;  wr_cycle[ 3977] = 1'b1;  addr_rom[ 3977]='h00003e24;  wr_data_rom[ 3977]='h000029d8;
    rd_cycle[ 3978] = 1'b0;  wr_cycle[ 3978] = 1'b1;  addr_rom[ 3978]='h00003e28;  wr_data_rom[ 3978]='h00002cef;
    rd_cycle[ 3979] = 1'b0;  wr_cycle[ 3979] = 1'b1;  addr_rom[ 3979]='h00003e2c;  wr_data_rom[ 3979]='h000015de;
    rd_cycle[ 3980] = 1'b0;  wr_cycle[ 3980] = 1'b1;  addr_rom[ 3980]='h00003e30;  wr_data_rom[ 3980]='h00001c43;
    rd_cycle[ 3981] = 1'b0;  wr_cycle[ 3981] = 1'b1;  addr_rom[ 3981]='h00003e34;  wr_data_rom[ 3981]='h00003ace;
    rd_cycle[ 3982] = 1'b0;  wr_cycle[ 3982] = 1'b1;  addr_rom[ 3982]='h00003e38;  wr_data_rom[ 3982]='h000009a7;
    rd_cycle[ 3983] = 1'b0;  wr_cycle[ 3983] = 1'b1;  addr_rom[ 3983]='h00003e3c;  wr_data_rom[ 3983]='h00000969;
    rd_cycle[ 3984] = 1'b0;  wr_cycle[ 3984] = 1'b1;  addr_rom[ 3984]='h00003e40;  wr_data_rom[ 3984]='h000023ce;
    rd_cycle[ 3985] = 1'b0;  wr_cycle[ 3985] = 1'b1;  addr_rom[ 3985]='h00003e44;  wr_data_rom[ 3985]='h00003717;
    rd_cycle[ 3986] = 1'b0;  wr_cycle[ 3986] = 1'b1;  addr_rom[ 3986]='h00003e48;  wr_data_rom[ 3986]='h00002c05;
    rd_cycle[ 3987] = 1'b0;  wr_cycle[ 3987] = 1'b1;  addr_rom[ 3987]='h00003e4c;  wr_data_rom[ 3987]='h00002a3b;
    rd_cycle[ 3988] = 1'b0;  wr_cycle[ 3988] = 1'b1;  addr_rom[ 3988]='h00003e50;  wr_data_rom[ 3988]='h000013c8;
    rd_cycle[ 3989] = 1'b0;  wr_cycle[ 3989] = 1'b1;  addr_rom[ 3989]='h00003e54;  wr_data_rom[ 3989]='h00001170;
    rd_cycle[ 3990] = 1'b0;  wr_cycle[ 3990] = 1'b1;  addr_rom[ 3990]='h00003e58;  wr_data_rom[ 3990]='h000014d6;
    rd_cycle[ 3991] = 1'b0;  wr_cycle[ 3991] = 1'b1;  addr_rom[ 3991]='h00003e5c;  wr_data_rom[ 3991]='h0000340d;
    rd_cycle[ 3992] = 1'b0;  wr_cycle[ 3992] = 1'b1;  addr_rom[ 3992]='h00003e60;  wr_data_rom[ 3992]='h00002f27;
    rd_cycle[ 3993] = 1'b0;  wr_cycle[ 3993] = 1'b1;  addr_rom[ 3993]='h00003e64;  wr_data_rom[ 3993]='h00003ac1;
    rd_cycle[ 3994] = 1'b0;  wr_cycle[ 3994] = 1'b1;  addr_rom[ 3994]='h00003e68;  wr_data_rom[ 3994]='h00001a68;
    rd_cycle[ 3995] = 1'b0;  wr_cycle[ 3995] = 1'b1;  addr_rom[ 3995]='h00003e6c;  wr_data_rom[ 3995]='h000031c7;
    rd_cycle[ 3996] = 1'b0;  wr_cycle[ 3996] = 1'b1;  addr_rom[ 3996]='h00003e70;  wr_data_rom[ 3996]='h00001128;
    rd_cycle[ 3997] = 1'b0;  wr_cycle[ 3997] = 1'b1;  addr_rom[ 3997]='h00003e74;  wr_data_rom[ 3997]='h00002320;
    rd_cycle[ 3998] = 1'b0;  wr_cycle[ 3998] = 1'b1;  addr_rom[ 3998]='h00003e78;  wr_data_rom[ 3998]='h00001325;
    rd_cycle[ 3999] = 1'b0;  wr_cycle[ 3999] = 1'b1;  addr_rom[ 3999]='h00003e7c;  wr_data_rom[ 3999]='h000013df;
    rd_cycle[ 4000] = 1'b0;  wr_cycle[ 4000] = 1'b1;  addr_rom[ 4000]='h00003e80;  wr_data_rom[ 4000]='h00001224;
    rd_cycle[ 4001] = 1'b0;  wr_cycle[ 4001] = 1'b1;  addr_rom[ 4001]='h00003e84;  wr_data_rom[ 4001]='h00003244;
    rd_cycle[ 4002] = 1'b0;  wr_cycle[ 4002] = 1'b1;  addr_rom[ 4002]='h00003e88;  wr_data_rom[ 4002]='h00000a18;
    rd_cycle[ 4003] = 1'b0;  wr_cycle[ 4003] = 1'b1;  addr_rom[ 4003]='h00003e8c;  wr_data_rom[ 4003]='h00001613;
    rd_cycle[ 4004] = 1'b0;  wr_cycle[ 4004] = 1'b1;  addr_rom[ 4004]='h00003e90;  wr_data_rom[ 4004]='h00003d3f;
    rd_cycle[ 4005] = 1'b0;  wr_cycle[ 4005] = 1'b1;  addr_rom[ 4005]='h00003e94;  wr_data_rom[ 4005]='h00001d0f;
    rd_cycle[ 4006] = 1'b0;  wr_cycle[ 4006] = 1'b1;  addr_rom[ 4006]='h00003e98;  wr_data_rom[ 4006]='h00001854;
    rd_cycle[ 4007] = 1'b0;  wr_cycle[ 4007] = 1'b1;  addr_rom[ 4007]='h00003e9c;  wr_data_rom[ 4007]='h000011e6;
    rd_cycle[ 4008] = 1'b0;  wr_cycle[ 4008] = 1'b1;  addr_rom[ 4008]='h00003ea0;  wr_data_rom[ 4008]='h00001b27;
    rd_cycle[ 4009] = 1'b0;  wr_cycle[ 4009] = 1'b1;  addr_rom[ 4009]='h00003ea4;  wr_data_rom[ 4009]='h000012b1;
    rd_cycle[ 4010] = 1'b0;  wr_cycle[ 4010] = 1'b1;  addr_rom[ 4010]='h00003ea8;  wr_data_rom[ 4010]='h0000358b;
    rd_cycle[ 4011] = 1'b0;  wr_cycle[ 4011] = 1'b1;  addr_rom[ 4011]='h00003eac;  wr_data_rom[ 4011]='h0000140d;
    rd_cycle[ 4012] = 1'b0;  wr_cycle[ 4012] = 1'b1;  addr_rom[ 4012]='h00003eb0;  wr_data_rom[ 4012]='h000002ea;
    rd_cycle[ 4013] = 1'b0;  wr_cycle[ 4013] = 1'b1;  addr_rom[ 4013]='h00003eb4;  wr_data_rom[ 4013]='h000034d6;
    rd_cycle[ 4014] = 1'b0;  wr_cycle[ 4014] = 1'b1;  addr_rom[ 4014]='h00003eb8;  wr_data_rom[ 4014]='h0000364b;
    rd_cycle[ 4015] = 1'b0;  wr_cycle[ 4015] = 1'b1;  addr_rom[ 4015]='h00003ebc;  wr_data_rom[ 4015]='h00000596;
    rd_cycle[ 4016] = 1'b0;  wr_cycle[ 4016] = 1'b1;  addr_rom[ 4016]='h00003ec0;  wr_data_rom[ 4016]='h00003b47;
    rd_cycle[ 4017] = 1'b0;  wr_cycle[ 4017] = 1'b1;  addr_rom[ 4017]='h00003ec4;  wr_data_rom[ 4017]='h000022e0;
    rd_cycle[ 4018] = 1'b0;  wr_cycle[ 4018] = 1'b1;  addr_rom[ 4018]='h00003ec8;  wr_data_rom[ 4018]='h00002f24;
    rd_cycle[ 4019] = 1'b0;  wr_cycle[ 4019] = 1'b1;  addr_rom[ 4019]='h00003ecc;  wr_data_rom[ 4019]='h00000103;
    rd_cycle[ 4020] = 1'b0;  wr_cycle[ 4020] = 1'b1;  addr_rom[ 4020]='h00003ed0;  wr_data_rom[ 4020]='h00003ee4;
    rd_cycle[ 4021] = 1'b0;  wr_cycle[ 4021] = 1'b1;  addr_rom[ 4021]='h00003ed4;  wr_data_rom[ 4021]='h00002247;
    rd_cycle[ 4022] = 1'b0;  wr_cycle[ 4022] = 1'b1;  addr_rom[ 4022]='h00003ed8;  wr_data_rom[ 4022]='h00001366;
    rd_cycle[ 4023] = 1'b0;  wr_cycle[ 4023] = 1'b1;  addr_rom[ 4023]='h00003edc;  wr_data_rom[ 4023]='h000011d6;
    rd_cycle[ 4024] = 1'b0;  wr_cycle[ 4024] = 1'b1;  addr_rom[ 4024]='h00003ee0;  wr_data_rom[ 4024]='h00003e5f;
    rd_cycle[ 4025] = 1'b0;  wr_cycle[ 4025] = 1'b1;  addr_rom[ 4025]='h00003ee4;  wr_data_rom[ 4025]='h00003393;
    rd_cycle[ 4026] = 1'b0;  wr_cycle[ 4026] = 1'b1;  addr_rom[ 4026]='h00003ee8;  wr_data_rom[ 4026]='h00003af6;
    rd_cycle[ 4027] = 1'b0;  wr_cycle[ 4027] = 1'b1;  addr_rom[ 4027]='h00003eec;  wr_data_rom[ 4027]='h000024c9;
    rd_cycle[ 4028] = 1'b0;  wr_cycle[ 4028] = 1'b1;  addr_rom[ 4028]='h00003ef0;  wr_data_rom[ 4028]='h00001b71;
    rd_cycle[ 4029] = 1'b0;  wr_cycle[ 4029] = 1'b1;  addr_rom[ 4029]='h00003ef4;  wr_data_rom[ 4029]='h00000f6a;
    rd_cycle[ 4030] = 1'b0;  wr_cycle[ 4030] = 1'b1;  addr_rom[ 4030]='h00003ef8;  wr_data_rom[ 4030]='h00001bb6;
    rd_cycle[ 4031] = 1'b0;  wr_cycle[ 4031] = 1'b1;  addr_rom[ 4031]='h00003efc;  wr_data_rom[ 4031]='h00003204;
    rd_cycle[ 4032] = 1'b0;  wr_cycle[ 4032] = 1'b1;  addr_rom[ 4032]='h00003f00;  wr_data_rom[ 4032]='h00002e31;
    rd_cycle[ 4033] = 1'b0;  wr_cycle[ 4033] = 1'b1;  addr_rom[ 4033]='h00003f04;  wr_data_rom[ 4033]='h00002e2c;
    rd_cycle[ 4034] = 1'b0;  wr_cycle[ 4034] = 1'b1;  addr_rom[ 4034]='h00003f08;  wr_data_rom[ 4034]='h0000328b;
    rd_cycle[ 4035] = 1'b0;  wr_cycle[ 4035] = 1'b1;  addr_rom[ 4035]='h00003f0c;  wr_data_rom[ 4035]='h00001e3e;
    rd_cycle[ 4036] = 1'b0;  wr_cycle[ 4036] = 1'b1;  addr_rom[ 4036]='h00003f10;  wr_data_rom[ 4036]='h000022b3;
    rd_cycle[ 4037] = 1'b0;  wr_cycle[ 4037] = 1'b1;  addr_rom[ 4037]='h00003f14;  wr_data_rom[ 4037]='h000015b3;
    rd_cycle[ 4038] = 1'b0;  wr_cycle[ 4038] = 1'b1;  addr_rom[ 4038]='h00003f18;  wr_data_rom[ 4038]='h00001ab1;
    rd_cycle[ 4039] = 1'b0;  wr_cycle[ 4039] = 1'b1;  addr_rom[ 4039]='h00003f1c;  wr_data_rom[ 4039]='h00001177;
    rd_cycle[ 4040] = 1'b0;  wr_cycle[ 4040] = 1'b1;  addr_rom[ 4040]='h00003f20;  wr_data_rom[ 4040]='h00003f0a;
    rd_cycle[ 4041] = 1'b0;  wr_cycle[ 4041] = 1'b1;  addr_rom[ 4041]='h00003f24;  wr_data_rom[ 4041]='h00000459;
    rd_cycle[ 4042] = 1'b0;  wr_cycle[ 4042] = 1'b1;  addr_rom[ 4042]='h00003f28;  wr_data_rom[ 4042]='h0000127e;
    rd_cycle[ 4043] = 1'b0;  wr_cycle[ 4043] = 1'b1;  addr_rom[ 4043]='h00003f2c;  wr_data_rom[ 4043]='h00000f03;
    rd_cycle[ 4044] = 1'b0;  wr_cycle[ 4044] = 1'b1;  addr_rom[ 4044]='h00003f30;  wr_data_rom[ 4044]='h000030b1;
    rd_cycle[ 4045] = 1'b0;  wr_cycle[ 4045] = 1'b1;  addr_rom[ 4045]='h00003f34;  wr_data_rom[ 4045]='h00002d7d;
    rd_cycle[ 4046] = 1'b0;  wr_cycle[ 4046] = 1'b1;  addr_rom[ 4046]='h00003f38;  wr_data_rom[ 4046]='h0000323f;
    rd_cycle[ 4047] = 1'b0;  wr_cycle[ 4047] = 1'b1;  addr_rom[ 4047]='h00003f3c;  wr_data_rom[ 4047]='h0000017e;
    rd_cycle[ 4048] = 1'b0;  wr_cycle[ 4048] = 1'b1;  addr_rom[ 4048]='h00003f40;  wr_data_rom[ 4048]='h000017d3;
    rd_cycle[ 4049] = 1'b0;  wr_cycle[ 4049] = 1'b1;  addr_rom[ 4049]='h00003f44;  wr_data_rom[ 4049]='h0000323e;
    rd_cycle[ 4050] = 1'b0;  wr_cycle[ 4050] = 1'b1;  addr_rom[ 4050]='h00003f48;  wr_data_rom[ 4050]='h00002a68;
    rd_cycle[ 4051] = 1'b0;  wr_cycle[ 4051] = 1'b1;  addr_rom[ 4051]='h00003f4c;  wr_data_rom[ 4051]='h00003885;
    rd_cycle[ 4052] = 1'b0;  wr_cycle[ 4052] = 1'b1;  addr_rom[ 4052]='h00003f50;  wr_data_rom[ 4052]='h000031b4;
    rd_cycle[ 4053] = 1'b0;  wr_cycle[ 4053] = 1'b1;  addr_rom[ 4053]='h00003f54;  wr_data_rom[ 4053]='h00002c6c;
    rd_cycle[ 4054] = 1'b0;  wr_cycle[ 4054] = 1'b1;  addr_rom[ 4054]='h00003f58;  wr_data_rom[ 4054]='h00000932;
    rd_cycle[ 4055] = 1'b0;  wr_cycle[ 4055] = 1'b1;  addr_rom[ 4055]='h00003f5c;  wr_data_rom[ 4055]='h000024d6;
    rd_cycle[ 4056] = 1'b0;  wr_cycle[ 4056] = 1'b1;  addr_rom[ 4056]='h00003f60;  wr_data_rom[ 4056]='h00002a8e;
    rd_cycle[ 4057] = 1'b0;  wr_cycle[ 4057] = 1'b1;  addr_rom[ 4057]='h00003f64;  wr_data_rom[ 4057]='h00001ab8;
    rd_cycle[ 4058] = 1'b0;  wr_cycle[ 4058] = 1'b1;  addr_rom[ 4058]='h00003f68;  wr_data_rom[ 4058]='h0000185d;
    rd_cycle[ 4059] = 1'b0;  wr_cycle[ 4059] = 1'b1;  addr_rom[ 4059]='h00003f6c;  wr_data_rom[ 4059]='h00002e38;
    rd_cycle[ 4060] = 1'b0;  wr_cycle[ 4060] = 1'b1;  addr_rom[ 4060]='h00003f70;  wr_data_rom[ 4060]='h0000009a;
    rd_cycle[ 4061] = 1'b0;  wr_cycle[ 4061] = 1'b1;  addr_rom[ 4061]='h00003f74;  wr_data_rom[ 4061]='h00002ce7;
    rd_cycle[ 4062] = 1'b0;  wr_cycle[ 4062] = 1'b1;  addr_rom[ 4062]='h00003f78;  wr_data_rom[ 4062]='h00001ca5;
    rd_cycle[ 4063] = 1'b0;  wr_cycle[ 4063] = 1'b1;  addr_rom[ 4063]='h00003f7c;  wr_data_rom[ 4063]='h0000161b;
    rd_cycle[ 4064] = 1'b0;  wr_cycle[ 4064] = 1'b1;  addr_rom[ 4064]='h00003f80;  wr_data_rom[ 4064]='h000004d2;
    rd_cycle[ 4065] = 1'b0;  wr_cycle[ 4065] = 1'b1;  addr_rom[ 4065]='h00003f84;  wr_data_rom[ 4065]='h000012e3;
    rd_cycle[ 4066] = 1'b0;  wr_cycle[ 4066] = 1'b1;  addr_rom[ 4066]='h00003f88;  wr_data_rom[ 4066]='h0000162b;
    rd_cycle[ 4067] = 1'b0;  wr_cycle[ 4067] = 1'b1;  addr_rom[ 4067]='h00003f8c;  wr_data_rom[ 4067]='h00001bed;
    rd_cycle[ 4068] = 1'b0;  wr_cycle[ 4068] = 1'b1;  addr_rom[ 4068]='h00003f90;  wr_data_rom[ 4068]='h0000073f;
    rd_cycle[ 4069] = 1'b0;  wr_cycle[ 4069] = 1'b1;  addr_rom[ 4069]='h00003f94;  wr_data_rom[ 4069]='h00003b88;
    rd_cycle[ 4070] = 1'b0;  wr_cycle[ 4070] = 1'b1;  addr_rom[ 4070]='h00003f98;  wr_data_rom[ 4070]='h00000bf7;
    rd_cycle[ 4071] = 1'b0;  wr_cycle[ 4071] = 1'b1;  addr_rom[ 4071]='h00003f9c;  wr_data_rom[ 4071]='h000024cd;
    rd_cycle[ 4072] = 1'b0;  wr_cycle[ 4072] = 1'b1;  addr_rom[ 4072]='h00003fa0;  wr_data_rom[ 4072]='h00002f3f;
    rd_cycle[ 4073] = 1'b0;  wr_cycle[ 4073] = 1'b1;  addr_rom[ 4073]='h00003fa4;  wr_data_rom[ 4073]='h0000293d;
    rd_cycle[ 4074] = 1'b0;  wr_cycle[ 4074] = 1'b1;  addr_rom[ 4074]='h00003fa8;  wr_data_rom[ 4074]='h00003a8f;
    rd_cycle[ 4075] = 1'b0;  wr_cycle[ 4075] = 1'b1;  addr_rom[ 4075]='h00003fac;  wr_data_rom[ 4075]='h00001a15;
    rd_cycle[ 4076] = 1'b0;  wr_cycle[ 4076] = 1'b1;  addr_rom[ 4076]='h00003fb0;  wr_data_rom[ 4076]='h00003ddd;
    rd_cycle[ 4077] = 1'b0;  wr_cycle[ 4077] = 1'b1;  addr_rom[ 4077]='h00003fb4;  wr_data_rom[ 4077]='h00000210;
    rd_cycle[ 4078] = 1'b0;  wr_cycle[ 4078] = 1'b1;  addr_rom[ 4078]='h00003fb8;  wr_data_rom[ 4078]='h000035f0;
    rd_cycle[ 4079] = 1'b0;  wr_cycle[ 4079] = 1'b1;  addr_rom[ 4079]='h00003fbc;  wr_data_rom[ 4079]='h00001065;
    rd_cycle[ 4080] = 1'b0;  wr_cycle[ 4080] = 1'b1;  addr_rom[ 4080]='h00003fc0;  wr_data_rom[ 4080]='h00000b5a;
    rd_cycle[ 4081] = 1'b0;  wr_cycle[ 4081] = 1'b1;  addr_rom[ 4081]='h00003fc4;  wr_data_rom[ 4081]='h00001e4f;
    rd_cycle[ 4082] = 1'b0;  wr_cycle[ 4082] = 1'b1;  addr_rom[ 4082]='h00003fc8;  wr_data_rom[ 4082]='h00003d14;
    rd_cycle[ 4083] = 1'b0;  wr_cycle[ 4083] = 1'b1;  addr_rom[ 4083]='h00003fcc;  wr_data_rom[ 4083]='h0000244b;
    rd_cycle[ 4084] = 1'b0;  wr_cycle[ 4084] = 1'b1;  addr_rom[ 4084]='h00003fd0;  wr_data_rom[ 4084]='h00000268;
    rd_cycle[ 4085] = 1'b0;  wr_cycle[ 4085] = 1'b1;  addr_rom[ 4085]='h00003fd4;  wr_data_rom[ 4085]='h00002087;
    rd_cycle[ 4086] = 1'b0;  wr_cycle[ 4086] = 1'b1;  addr_rom[ 4086]='h00003fd8;  wr_data_rom[ 4086]='h00002781;
    rd_cycle[ 4087] = 1'b0;  wr_cycle[ 4087] = 1'b1;  addr_rom[ 4087]='h00003fdc;  wr_data_rom[ 4087]='h0000371c;
    rd_cycle[ 4088] = 1'b0;  wr_cycle[ 4088] = 1'b1;  addr_rom[ 4088]='h00003fe0;  wr_data_rom[ 4088]='h0000366f;
    rd_cycle[ 4089] = 1'b0;  wr_cycle[ 4089] = 1'b1;  addr_rom[ 4089]='h00003fe4;  wr_data_rom[ 4089]='h000026e3;
    rd_cycle[ 4090] = 1'b0;  wr_cycle[ 4090] = 1'b1;  addr_rom[ 4090]='h00003fe8;  wr_data_rom[ 4090]='h000009ce;
    rd_cycle[ 4091] = 1'b0;  wr_cycle[ 4091] = 1'b1;  addr_rom[ 4091]='h00003fec;  wr_data_rom[ 4091]='h00003e0e;
    rd_cycle[ 4092] = 1'b0;  wr_cycle[ 4092] = 1'b1;  addr_rom[ 4092]='h00003ff0;  wr_data_rom[ 4092]='h00000d12;
    rd_cycle[ 4093] = 1'b0;  wr_cycle[ 4093] = 1'b1;  addr_rom[ 4093]='h00003ff4;  wr_data_rom[ 4093]='h00002bf9;
    rd_cycle[ 4094] = 1'b0;  wr_cycle[ 4094] = 1'b1;  addr_rom[ 4094]='h00003ff8;  wr_data_rom[ 4094]='h00000981;
    rd_cycle[ 4095] = 1'b0;  wr_cycle[ 4095] = 1'b1;  addr_rom[ 4095]='h00003ffc;  wr_data_rom[ 4095]='h00002d42;
    // 12288 random read and write cycles
    rd_cycle[ 4096] = 1'b0;  wr_cycle[ 4096] = 1'b1;  addr_rom[ 4096]='h00000634;  wr_data_rom[ 4096]='h00001de4;
    rd_cycle[ 4097] = 1'b0;  wr_cycle[ 4097] = 1'b1;  addr_rom[ 4097]='h00003cf0;  wr_data_rom[ 4097]='h0000123c;
    rd_cycle[ 4098] = 1'b1;  wr_cycle[ 4098] = 1'b0;  addr_rom[ 4098]='h00003c2c;  wr_data_rom[ 4098]='h00000000;
    rd_cycle[ 4099] = 1'b0;  wr_cycle[ 4099] = 1'b1;  addr_rom[ 4099]='h00001460;  wr_data_rom[ 4099]='h000012a3;
    rd_cycle[ 4100] = 1'b1;  wr_cycle[ 4100] = 1'b0;  addr_rom[ 4100]='h00000fe4;  wr_data_rom[ 4100]='h00000000;
    rd_cycle[ 4101] = 1'b0;  wr_cycle[ 4101] = 1'b1;  addr_rom[ 4101]='h00002060;  wr_data_rom[ 4101]='h000026ff;
    rd_cycle[ 4102] = 1'b1;  wr_cycle[ 4102] = 1'b0;  addr_rom[ 4102]='h00003e6c;  wr_data_rom[ 4102]='h00000000;
    rd_cycle[ 4103] = 1'b0;  wr_cycle[ 4103] = 1'b1;  addr_rom[ 4103]='h00002e98;  wr_data_rom[ 4103]='h00003157;
    rd_cycle[ 4104] = 1'b1;  wr_cycle[ 4104] = 1'b0;  addr_rom[ 4104]='h00002c80;  wr_data_rom[ 4104]='h00000000;
    rd_cycle[ 4105] = 1'b1;  wr_cycle[ 4105] = 1'b0;  addr_rom[ 4105]='h000033b0;  wr_data_rom[ 4105]='h00000000;
    rd_cycle[ 4106] = 1'b0;  wr_cycle[ 4106] = 1'b1;  addr_rom[ 4106]='h000022cc;  wr_data_rom[ 4106]='h00000ec4;
    rd_cycle[ 4107] = 1'b1;  wr_cycle[ 4107] = 1'b0;  addr_rom[ 4107]='h00001314;  wr_data_rom[ 4107]='h00000000;
    rd_cycle[ 4108] = 1'b0;  wr_cycle[ 4108] = 1'b1;  addr_rom[ 4108]='h000003b4;  wr_data_rom[ 4108]='h00001057;
    rd_cycle[ 4109] = 1'b1;  wr_cycle[ 4109] = 1'b0;  addr_rom[ 4109]='h00000478;  wr_data_rom[ 4109]='h00000000;
    rd_cycle[ 4110] = 1'b1;  wr_cycle[ 4110] = 1'b0;  addr_rom[ 4110]='h000003b0;  wr_data_rom[ 4110]='h00000000;
    rd_cycle[ 4111] = 1'b0;  wr_cycle[ 4111] = 1'b1;  addr_rom[ 4111]='h00000e84;  wr_data_rom[ 4111]='h00001819;
    rd_cycle[ 4112] = 1'b0;  wr_cycle[ 4112] = 1'b1;  addr_rom[ 4112]='h00000658;  wr_data_rom[ 4112]='h00002586;
    rd_cycle[ 4113] = 1'b0;  wr_cycle[ 4113] = 1'b1;  addr_rom[ 4113]='h00003178;  wr_data_rom[ 4113]='h00000734;
    rd_cycle[ 4114] = 1'b0;  wr_cycle[ 4114] = 1'b1;  addr_rom[ 4114]='h00003f6c;  wr_data_rom[ 4114]='h00003ad1;
    rd_cycle[ 4115] = 1'b1;  wr_cycle[ 4115] = 1'b0;  addr_rom[ 4115]='h00002dc8;  wr_data_rom[ 4115]='h00000000;
    rd_cycle[ 4116] = 1'b1;  wr_cycle[ 4116] = 1'b0;  addr_rom[ 4116]='h000030fc;  wr_data_rom[ 4116]='h00000000;
    rd_cycle[ 4117] = 1'b1;  wr_cycle[ 4117] = 1'b0;  addr_rom[ 4117]='h000026a4;  wr_data_rom[ 4117]='h00000000;
    rd_cycle[ 4118] = 1'b0;  wr_cycle[ 4118] = 1'b1;  addr_rom[ 4118]='h000034e0;  wr_data_rom[ 4118]='h00001518;
    rd_cycle[ 4119] = 1'b1;  wr_cycle[ 4119] = 1'b0;  addr_rom[ 4119]='h00001b78;  wr_data_rom[ 4119]='h00000000;
    rd_cycle[ 4120] = 1'b1;  wr_cycle[ 4120] = 1'b0;  addr_rom[ 4120]='h00002968;  wr_data_rom[ 4120]='h00000000;
    rd_cycle[ 4121] = 1'b0;  wr_cycle[ 4121] = 1'b1;  addr_rom[ 4121]='h00000208;  wr_data_rom[ 4121]='h00002953;
    rd_cycle[ 4122] = 1'b1;  wr_cycle[ 4122] = 1'b0;  addr_rom[ 4122]='h0000325c;  wr_data_rom[ 4122]='h00000000;
    rd_cycle[ 4123] = 1'b0;  wr_cycle[ 4123] = 1'b1;  addr_rom[ 4123]='h00000bc8;  wr_data_rom[ 4123]='h00002897;
    rd_cycle[ 4124] = 1'b1;  wr_cycle[ 4124] = 1'b0;  addr_rom[ 4124]='h0000365c;  wr_data_rom[ 4124]='h00000000;
    rd_cycle[ 4125] = 1'b1;  wr_cycle[ 4125] = 1'b0;  addr_rom[ 4125]='h000006a4;  wr_data_rom[ 4125]='h00000000;
    rd_cycle[ 4126] = 1'b1;  wr_cycle[ 4126] = 1'b0;  addr_rom[ 4126]='h00002a64;  wr_data_rom[ 4126]='h00000000;
    rd_cycle[ 4127] = 1'b1;  wr_cycle[ 4127] = 1'b0;  addr_rom[ 4127]='h00000d20;  wr_data_rom[ 4127]='h00000000;
    rd_cycle[ 4128] = 1'b1;  wr_cycle[ 4128] = 1'b0;  addr_rom[ 4128]='h0000020c;  wr_data_rom[ 4128]='h00000000;
    rd_cycle[ 4129] = 1'b0;  wr_cycle[ 4129] = 1'b1;  addr_rom[ 4129]='h000032a4;  wr_data_rom[ 4129]='h000035f5;
    rd_cycle[ 4130] = 1'b0;  wr_cycle[ 4130] = 1'b1;  addr_rom[ 4130]='h0000212c;  wr_data_rom[ 4130]='h000027cd;
    rd_cycle[ 4131] = 1'b1;  wr_cycle[ 4131] = 1'b0;  addr_rom[ 4131]='h00000778;  wr_data_rom[ 4131]='h00000000;
    rd_cycle[ 4132] = 1'b1;  wr_cycle[ 4132] = 1'b0;  addr_rom[ 4132]='h0000256c;  wr_data_rom[ 4132]='h00000000;
    rd_cycle[ 4133] = 1'b0;  wr_cycle[ 4133] = 1'b1;  addr_rom[ 4133]='h000010cc;  wr_data_rom[ 4133]='h00001946;
    rd_cycle[ 4134] = 1'b1;  wr_cycle[ 4134] = 1'b0;  addr_rom[ 4134]='h000014b4;  wr_data_rom[ 4134]='h00000000;
    rd_cycle[ 4135] = 1'b1;  wr_cycle[ 4135] = 1'b0;  addr_rom[ 4135]='h000017bc;  wr_data_rom[ 4135]='h00000000;
    rd_cycle[ 4136] = 1'b1;  wr_cycle[ 4136] = 1'b0;  addr_rom[ 4136]='h0000164c;  wr_data_rom[ 4136]='h00000000;
    rd_cycle[ 4137] = 1'b0;  wr_cycle[ 4137] = 1'b1;  addr_rom[ 4137]='h00002684;  wr_data_rom[ 4137]='h00000f91;
    rd_cycle[ 4138] = 1'b1;  wr_cycle[ 4138] = 1'b0;  addr_rom[ 4138]='h00000530;  wr_data_rom[ 4138]='h00000000;
    rd_cycle[ 4139] = 1'b1;  wr_cycle[ 4139] = 1'b0;  addr_rom[ 4139]='h00003724;  wr_data_rom[ 4139]='h00000000;
    rd_cycle[ 4140] = 1'b0;  wr_cycle[ 4140] = 1'b1;  addr_rom[ 4140]='h000015a8;  wr_data_rom[ 4140]='h00002bc0;
    rd_cycle[ 4141] = 1'b1;  wr_cycle[ 4141] = 1'b0;  addr_rom[ 4141]='h00003140;  wr_data_rom[ 4141]='h00000000;
    rd_cycle[ 4142] = 1'b0;  wr_cycle[ 4142] = 1'b1;  addr_rom[ 4142]='h000023a0;  wr_data_rom[ 4142]='h00000a9c;
    rd_cycle[ 4143] = 1'b1;  wr_cycle[ 4143] = 1'b0;  addr_rom[ 4143]='h000012f4;  wr_data_rom[ 4143]='h00000000;
    rd_cycle[ 4144] = 1'b0;  wr_cycle[ 4144] = 1'b1;  addr_rom[ 4144]='h000024d0;  wr_data_rom[ 4144]='h00000557;
    rd_cycle[ 4145] = 1'b1;  wr_cycle[ 4145] = 1'b0;  addr_rom[ 4145]='h00003b18;  wr_data_rom[ 4145]='h00000000;
    rd_cycle[ 4146] = 1'b0;  wr_cycle[ 4146] = 1'b1;  addr_rom[ 4146]='h00001470;  wr_data_rom[ 4146]='h00000fa7;
    rd_cycle[ 4147] = 1'b0;  wr_cycle[ 4147] = 1'b1;  addr_rom[ 4147]='h000035e4;  wr_data_rom[ 4147]='h0000349a;
    rd_cycle[ 4148] = 1'b1;  wr_cycle[ 4148] = 1'b0;  addr_rom[ 4148]='h000037c8;  wr_data_rom[ 4148]='h00000000;
    rd_cycle[ 4149] = 1'b1;  wr_cycle[ 4149] = 1'b0;  addr_rom[ 4149]='h00002078;  wr_data_rom[ 4149]='h00000000;
    rd_cycle[ 4150] = 1'b0;  wr_cycle[ 4150] = 1'b1;  addr_rom[ 4150]='h00002b08;  wr_data_rom[ 4150]='h00003e8e;
    rd_cycle[ 4151] = 1'b0;  wr_cycle[ 4151] = 1'b1;  addr_rom[ 4151]='h00002f30;  wr_data_rom[ 4151]='h00000705;
    rd_cycle[ 4152] = 1'b1;  wr_cycle[ 4152] = 1'b0;  addr_rom[ 4152]='h00002230;  wr_data_rom[ 4152]='h00000000;
    rd_cycle[ 4153] = 1'b0;  wr_cycle[ 4153] = 1'b1;  addr_rom[ 4153]='h00001108;  wr_data_rom[ 4153]='h000036a3;
    rd_cycle[ 4154] = 1'b1;  wr_cycle[ 4154] = 1'b0;  addr_rom[ 4154]='h000006b0;  wr_data_rom[ 4154]='h00000000;
    rd_cycle[ 4155] = 1'b1;  wr_cycle[ 4155] = 1'b0;  addr_rom[ 4155]='h00001524;  wr_data_rom[ 4155]='h00000000;
    rd_cycle[ 4156] = 1'b0;  wr_cycle[ 4156] = 1'b1;  addr_rom[ 4156]='h000039a0;  wr_data_rom[ 4156]='h000020f7;
    rd_cycle[ 4157] = 1'b0;  wr_cycle[ 4157] = 1'b1;  addr_rom[ 4157]='h0000320c;  wr_data_rom[ 4157]='h00003b66;
    rd_cycle[ 4158] = 1'b1;  wr_cycle[ 4158] = 1'b0;  addr_rom[ 4158]='h00003bac;  wr_data_rom[ 4158]='h00000000;
    rd_cycle[ 4159] = 1'b0;  wr_cycle[ 4159] = 1'b1;  addr_rom[ 4159]='h00001c04;  wr_data_rom[ 4159]='h00000dc9;
    rd_cycle[ 4160] = 1'b1;  wr_cycle[ 4160] = 1'b0;  addr_rom[ 4160]='h00002938;  wr_data_rom[ 4160]='h00000000;
    rd_cycle[ 4161] = 1'b0;  wr_cycle[ 4161] = 1'b1;  addr_rom[ 4161]='h00003f30;  wr_data_rom[ 4161]='h00002c7b;
    rd_cycle[ 4162] = 1'b1;  wr_cycle[ 4162] = 1'b0;  addr_rom[ 4162]='h00002a28;  wr_data_rom[ 4162]='h00000000;
    rd_cycle[ 4163] = 1'b0;  wr_cycle[ 4163] = 1'b1;  addr_rom[ 4163]='h00003acc;  wr_data_rom[ 4163]='h00000986;
    rd_cycle[ 4164] = 1'b1;  wr_cycle[ 4164] = 1'b0;  addr_rom[ 4164]='h000015a0;  wr_data_rom[ 4164]='h00000000;
    rd_cycle[ 4165] = 1'b1;  wr_cycle[ 4165] = 1'b0;  addr_rom[ 4165]='h00003188;  wr_data_rom[ 4165]='h00000000;
    rd_cycle[ 4166] = 1'b1;  wr_cycle[ 4166] = 1'b0;  addr_rom[ 4166]='h00003d7c;  wr_data_rom[ 4166]='h00000000;
    rd_cycle[ 4167] = 1'b1;  wr_cycle[ 4167] = 1'b0;  addr_rom[ 4167]='h00003ff4;  wr_data_rom[ 4167]='h00000000;
    rd_cycle[ 4168] = 1'b0;  wr_cycle[ 4168] = 1'b1;  addr_rom[ 4168]='h0000060c;  wr_data_rom[ 4168]='h000025fd;
    rd_cycle[ 4169] = 1'b1;  wr_cycle[ 4169] = 1'b0;  addr_rom[ 4169]='h00000010;  wr_data_rom[ 4169]='h00000000;
    rd_cycle[ 4170] = 1'b0;  wr_cycle[ 4170] = 1'b1;  addr_rom[ 4170]='h000019ec;  wr_data_rom[ 4170]='h00002d10;
    rd_cycle[ 4171] = 1'b0;  wr_cycle[ 4171] = 1'b1;  addr_rom[ 4171]='h000020f8;  wr_data_rom[ 4171]='h000029d7;
    rd_cycle[ 4172] = 1'b0;  wr_cycle[ 4172] = 1'b1;  addr_rom[ 4172]='h00000f80;  wr_data_rom[ 4172]='h000029ac;
    rd_cycle[ 4173] = 1'b0;  wr_cycle[ 4173] = 1'b1;  addr_rom[ 4173]='h0000390c;  wr_data_rom[ 4173]='h00001cd0;
    rd_cycle[ 4174] = 1'b0;  wr_cycle[ 4174] = 1'b1;  addr_rom[ 4174]='h0000085c;  wr_data_rom[ 4174]='h000035e7;
    rd_cycle[ 4175] = 1'b0;  wr_cycle[ 4175] = 1'b1;  addr_rom[ 4175]='h000003ac;  wr_data_rom[ 4175]='h000016e5;
    rd_cycle[ 4176] = 1'b0;  wr_cycle[ 4176] = 1'b1;  addr_rom[ 4176]='h00003a60;  wr_data_rom[ 4176]='h00000a0e;
    rd_cycle[ 4177] = 1'b0;  wr_cycle[ 4177] = 1'b1;  addr_rom[ 4177]='h00001664;  wr_data_rom[ 4177]='h000028be;
    rd_cycle[ 4178] = 1'b1;  wr_cycle[ 4178] = 1'b0;  addr_rom[ 4178]='h00000a38;  wr_data_rom[ 4178]='h00000000;
    rd_cycle[ 4179] = 1'b1;  wr_cycle[ 4179] = 1'b0;  addr_rom[ 4179]='h00001cf8;  wr_data_rom[ 4179]='h00000000;
    rd_cycle[ 4180] = 1'b1;  wr_cycle[ 4180] = 1'b0;  addr_rom[ 4180]='h000007e4;  wr_data_rom[ 4180]='h00000000;
    rd_cycle[ 4181] = 1'b1;  wr_cycle[ 4181] = 1'b0;  addr_rom[ 4181]='h00000874;  wr_data_rom[ 4181]='h00000000;
    rd_cycle[ 4182] = 1'b0;  wr_cycle[ 4182] = 1'b1;  addr_rom[ 4182]='h000006f4;  wr_data_rom[ 4182]='h000021a2;
    rd_cycle[ 4183] = 1'b1;  wr_cycle[ 4183] = 1'b0;  addr_rom[ 4183]='h00001f34;  wr_data_rom[ 4183]='h00000000;
    rd_cycle[ 4184] = 1'b1;  wr_cycle[ 4184] = 1'b0;  addr_rom[ 4184]='h00002b44;  wr_data_rom[ 4184]='h00000000;
    rd_cycle[ 4185] = 1'b1;  wr_cycle[ 4185] = 1'b0;  addr_rom[ 4185]='h00001354;  wr_data_rom[ 4185]='h00000000;
    rd_cycle[ 4186] = 1'b1;  wr_cycle[ 4186] = 1'b0;  addr_rom[ 4186]='h00000768;  wr_data_rom[ 4186]='h00000000;
    rd_cycle[ 4187] = 1'b1;  wr_cycle[ 4187] = 1'b0;  addr_rom[ 4187]='h00002230;  wr_data_rom[ 4187]='h00000000;
    rd_cycle[ 4188] = 1'b1;  wr_cycle[ 4188] = 1'b0;  addr_rom[ 4188]='h00003510;  wr_data_rom[ 4188]='h00000000;
    rd_cycle[ 4189] = 1'b1;  wr_cycle[ 4189] = 1'b0;  addr_rom[ 4189]='h000028c8;  wr_data_rom[ 4189]='h00000000;
    rd_cycle[ 4190] = 1'b0;  wr_cycle[ 4190] = 1'b1;  addr_rom[ 4190]='h00000034;  wr_data_rom[ 4190]='h0000281e;
    rd_cycle[ 4191] = 1'b0;  wr_cycle[ 4191] = 1'b1;  addr_rom[ 4191]='h00002418;  wr_data_rom[ 4191]='h00000a05;
    rd_cycle[ 4192] = 1'b1;  wr_cycle[ 4192] = 1'b0;  addr_rom[ 4192]='h00000e80;  wr_data_rom[ 4192]='h00000000;
    rd_cycle[ 4193] = 1'b0;  wr_cycle[ 4193] = 1'b1;  addr_rom[ 4193]='h00000308;  wr_data_rom[ 4193]='h000023b5;
    rd_cycle[ 4194] = 1'b1;  wr_cycle[ 4194] = 1'b0;  addr_rom[ 4194]='h00001ef4;  wr_data_rom[ 4194]='h00000000;
    rd_cycle[ 4195] = 1'b1;  wr_cycle[ 4195] = 1'b0;  addr_rom[ 4195]='h00001850;  wr_data_rom[ 4195]='h00000000;
    rd_cycle[ 4196] = 1'b0;  wr_cycle[ 4196] = 1'b1;  addr_rom[ 4196]='h00002dec;  wr_data_rom[ 4196]='h00002dc7;
    rd_cycle[ 4197] = 1'b0;  wr_cycle[ 4197] = 1'b1;  addr_rom[ 4197]='h00000748;  wr_data_rom[ 4197]='h00001ea1;
    rd_cycle[ 4198] = 1'b0;  wr_cycle[ 4198] = 1'b1;  addr_rom[ 4198]='h00003cc4;  wr_data_rom[ 4198]='h00002723;
    rd_cycle[ 4199] = 1'b0;  wr_cycle[ 4199] = 1'b1;  addr_rom[ 4199]='h00002054;  wr_data_rom[ 4199]='h00003596;
    rd_cycle[ 4200] = 1'b1;  wr_cycle[ 4200] = 1'b0;  addr_rom[ 4200]='h000017c0;  wr_data_rom[ 4200]='h00000000;
    rd_cycle[ 4201] = 1'b0;  wr_cycle[ 4201] = 1'b1;  addr_rom[ 4201]='h00001c48;  wr_data_rom[ 4201]='h00000976;
    rd_cycle[ 4202] = 1'b1;  wr_cycle[ 4202] = 1'b0;  addr_rom[ 4202]='h00000f00;  wr_data_rom[ 4202]='h00000000;
    rd_cycle[ 4203] = 1'b1;  wr_cycle[ 4203] = 1'b0;  addr_rom[ 4203]='h0000277c;  wr_data_rom[ 4203]='h00000000;
    rd_cycle[ 4204] = 1'b1;  wr_cycle[ 4204] = 1'b0;  addr_rom[ 4204]='h00002db4;  wr_data_rom[ 4204]='h00000000;
    rd_cycle[ 4205] = 1'b0;  wr_cycle[ 4205] = 1'b1;  addr_rom[ 4205]='h000034e0;  wr_data_rom[ 4205]='h00000c0a;
    rd_cycle[ 4206] = 1'b1;  wr_cycle[ 4206] = 1'b0;  addr_rom[ 4206]='h00000a7c;  wr_data_rom[ 4206]='h00000000;
    rd_cycle[ 4207] = 1'b1;  wr_cycle[ 4207] = 1'b0;  addr_rom[ 4207]='h00001004;  wr_data_rom[ 4207]='h00000000;
    rd_cycle[ 4208] = 1'b0;  wr_cycle[ 4208] = 1'b1;  addr_rom[ 4208]='h000027d0;  wr_data_rom[ 4208]='h00001944;
    rd_cycle[ 4209] = 1'b1;  wr_cycle[ 4209] = 1'b0;  addr_rom[ 4209]='h000004c4;  wr_data_rom[ 4209]='h00000000;
    rd_cycle[ 4210] = 1'b1;  wr_cycle[ 4210] = 1'b0;  addr_rom[ 4210]='h00001110;  wr_data_rom[ 4210]='h00000000;
    rd_cycle[ 4211] = 1'b0;  wr_cycle[ 4211] = 1'b1;  addr_rom[ 4211]='h000022e0;  wr_data_rom[ 4211]='h00002f6d;
    rd_cycle[ 4212] = 1'b0;  wr_cycle[ 4212] = 1'b1;  addr_rom[ 4212]='h000005a0;  wr_data_rom[ 4212]='h0000116e;
    rd_cycle[ 4213] = 1'b0;  wr_cycle[ 4213] = 1'b1;  addr_rom[ 4213]='h00002ef0;  wr_data_rom[ 4213]='h00001862;
    rd_cycle[ 4214] = 1'b1;  wr_cycle[ 4214] = 1'b0;  addr_rom[ 4214]='h00000078;  wr_data_rom[ 4214]='h00000000;
    rd_cycle[ 4215] = 1'b1;  wr_cycle[ 4215] = 1'b0;  addr_rom[ 4215]='h0000272c;  wr_data_rom[ 4215]='h00000000;
    rd_cycle[ 4216] = 1'b1;  wr_cycle[ 4216] = 1'b0;  addr_rom[ 4216]='h000026a4;  wr_data_rom[ 4216]='h00000000;
    rd_cycle[ 4217] = 1'b1;  wr_cycle[ 4217] = 1'b0;  addr_rom[ 4217]='h00000c30;  wr_data_rom[ 4217]='h00000000;
    rd_cycle[ 4218] = 1'b1;  wr_cycle[ 4218] = 1'b0;  addr_rom[ 4218]='h00002e00;  wr_data_rom[ 4218]='h00000000;
    rd_cycle[ 4219] = 1'b1;  wr_cycle[ 4219] = 1'b0;  addr_rom[ 4219]='h00001258;  wr_data_rom[ 4219]='h00000000;
    rd_cycle[ 4220] = 1'b0;  wr_cycle[ 4220] = 1'b1;  addr_rom[ 4220]='h0000182c;  wr_data_rom[ 4220]='h000023c9;
    rd_cycle[ 4221] = 1'b0;  wr_cycle[ 4221] = 1'b1;  addr_rom[ 4221]='h00000730;  wr_data_rom[ 4221]='h00003c82;
    rd_cycle[ 4222] = 1'b0;  wr_cycle[ 4222] = 1'b1;  addr_rom[ 4222]='h00001600;  wr_data_rom[ 4222]='h00001acb;
    rd_cycle[ 4223] = 1'b0;  wr_cycle[ 4223] = 1'b1;  addr_rom[ 4223]='h00000188;  wr_data_rom[ 4223]='h00002a68;
    rd_cycle[ 4224] = 1'b0;  wr_cycle[ 4224] = 1'b1;  addr_rom[ 4224]='h0000168c;  wr_data_rom[ 4224]='h000039c5;
    rd_cycle[ 4225] = 1'b1;  wr_cycle[ 4225] = 1'b0;  addr_rom[ 4225]='h00001748;  wr_data_rom[ 4225]='h00000000;
    rd_cycle[ 4226] = 1'b1;  wr_cycle[ 4226] = 1'b0;  addr_rom[ 4226]='h00002900;  wr_data_rom[ 4226]='h00000000;
    rd_cycle[ 4227] = 1'b1;  wr_cycle[ 4227] = 1'b0;  addr_rom[ 4227]='h00002664;  wr_data_rom[ 4227]='h00000000;
    rd_cycle[ 4228] = 1'b1;  wr_cycle[ 4228] = 1'b0;  addr_rom[ 4228]='h00003b20;  wr_data_rom[ 4228]='h00000000;
    rd_cycle[ 4229] = 1'b0;  wr_cycle[ 4229] = 1'b1;  addr_rom[ 4229]='h00001820;  wr_data_rom[ 4229]='h00002033;
    rd_cycle[ 4230] = 1'b1;  wr_cycle[ 4230] = 1'b0;  addr_rom[ 4230]='h00002d88;  wr_data_rom[ 4230]='h00000000;
    rd_cycle[ 4231] = 1'b1;  wr_cycle[ 4231] = 1'b0;  addr_rom[ 4231]='h00003b68;  wr_data_rom[ 4231]='h00000000;
    rd_cycle[ 4232] = 1'b1;  wr_cycle[ 4232] = 1'b0;  addr_rom[ 4232]='h00003e60;  wr_data_rom[ 4232]='h00000000;
    rd_cycle[ 4233] = 1'b1;  wr_cycle[ 4233] = 1'b0;  addr_rom[ 4233]='h00003df0;  wr_data_rom[ 4233]='h00000000;
    rd_cycle[ 4234] = 1'b0;  wr_cycle[ 4234] = 1'b1;  addr_rom[ 4234]='h00003618;  wr_data_rom[ 4234]='h00003ab6;
    rd_cycle[ 4235] = 1'b0;  wr_cycle[ 4235] = 1'b1;  addr_rom[ 4235]='h00001424;  wr_data_rom[ 4235]='h000005fd;
    rd_cycle[ 4236] = 1'b1;  wr_cycle[ 4236] = 1'b0;  addr_rom[ 4236]='h000023e4;  wr_data_rom[ 4236]='h00000000;
    rd_cycle[ 4237] = 1'b1;  wr_cycle[ 4237] = 1'b0;  addr_rom[ 4237]='h00001d6c;  wr_data_rom[ 4237]='h00000000;
    rd_cycle[ 4238] = 1'b1;  wr_cycle[ 4238] = 1'b0;  addr_rom[ 4238]='h00002ec0;  wr_data_rom[ 4238]='h00000000;
    rd_cycle[ 4239] = 1'b1;  wr_cycle[ 4239] = 1'b0;  addr_rom[ 4239]='h0000029c;  wr_data_rom[ 4239]='h00000000;
    rd_cycle[ 4240] = 1'b0;  wr_cycle[ 4240] = 1'b1;  addr_rom[ 4240]='h00001a14;  wr_data_rom[ 4240]='h00001a03;
    rd_cycle[ 4241] = 1'b1;  wr_cycle[ 4241] = 1'b0;  addr_rom[ 4241]='h00002f68;  wr_data_rom[ 4241]='h00000000;
    rd_cycle[ 4242] = 1'b1;  wr_cycle[ 4242] = 1'b0;  addr_rom[ 4242]='h00001fc0;  wr_data_rom[ 4242]='h00000000;
    rd_cycle[ 4243] = 1'b0;  wr_cycle[ 4243] = 1'b1;  addr_rom[ 4243]='h00002784;  wr_data_rom[ 4243]='h00003ff0;
    rd_cycle[ 4244] = 1'b0;  wr_cycle[ 4244] = 1'b1;  addr_rom[ 4244]='h00001cdc;  wr_data_rom[ 4244]='h00001a69;
    rd_cycle[ 4245] = 1'b1;  wr_cycle[ 4245] = 1'b0;  addr_rom[ 4245]='h00002d54;  wr_data_rom[ 4245]='h00000000;
    rd_cycle[ 4246] = 1'b1;  wr_cycle[ 4246] = 1'b0;  addr_rom[ 4246]='h0000282c;  wr_data_rom[ 4246]='h00000000;
    rd_cycle[ 4247] = 1'b1;  wr_cycle[ 4247] = 1'b0;  addr_rom[ 4247]='h00002b7c;  wr_data_rom[ 4247]='h00000000;
    rd_cycle[ 4248] = 1'b1;  wr_cycle[ 4248] = 1'b0;  addr_rom[ 4248]='h00000430;  wr_data_rom[ 4248]='h00000000;
    rd_cycle[ 4249] = 1'b1;  wr_cycle[ 4249] = 1'b0;  addr_rom[ 4249]='h0000267c;  wr_data_rom[ 4249]='h00000000;
    rd_cycle[ 4250] = 1'b1;  wr_cycle[ 4250] = 1'b0;  addr_rom[ 4250]='h00002fc0;  wr_data_rom[ 4250]='h00000000;
    rd_cycle[ 4251] = 1'b1;  wr_cycle[ 4251] = 1'b0;  addr_rom[ 4251]='h00003d68;  wr_data_rom[ 4251]='h00000000;
    rd_cycle[ 4252] = 1'b1;  wr_cycle[ 4252] = 1'b0;  addr_rom[ 4252]='h00000bdc;  wr_data_rom[ 4252]='h00000000;
    rd_cycle[ 4253] = 1'b0;  wr_cycle[ 4253] = 1'b1;  addr_rom[ 4253]='h00000ed0;  wr_data_rom[ 4253]='h0000337b;
    rd_cycle[ 4254] = 1'b1;  wr_cycle[ 4254] = 1'b0;  addr_rom[ 4254]='h00003e38;  wr_data_rom[ 4254]='h00000000;
    rd_cycle[ 4255] = 1'b0;  wr_cycle[ 4255] = 1'b1;  addr_rom[ 4255]='h0000280c;  wr_data_rom[ 4255]='h0000210f;
    rd_cycle[ 4256] = 1'b0;  wr_cycle[ 4256] = 1'b1;  addr_rom[ 4256]='h00000704;  wr_data_rom[ 4256]='h00001226;
    rd_cycle[ 4257] = 1'b1;  wr_cycle[ 4257] = 1'b0;  addr_rom[ 4257]='h00000760;  wr_data_rom[ 4257]='h00000000;
    rd_cycle[ 4258] = 1'b0;  wr_cycle[ 4258] = 1'b1;  addr_rom[ 4258]='h000027b8;  wr_data_rom[ 4258]='h00003bef;
    rd_cycle[ 4259] = 1'b1;  wr_cycle[ 4259] = 1'b0;  addr_rom[ 4259]='h000003cc;  wr_data_rom[ 4259]='h00000000;
    rd_cycle[ 4260] = 1'b0;  wr_cycle[ 4260] = 1'b1;  addr_rom[ 4260]='h00001fd4;  wr_data_rom[ 4260]='h000038da;
    rd_cycle[ 4261] = 1'b1;  wr_cycle[ 4261] = 1'b0;  addr_rom[ 4261]='h00000fb4;  wr_data_rom[ 4261]='h00000000;
    rd_cycle[ 4262] = 1'b0;  wr_cycle[ 4262] = 1'b1;  addr_rom[ 4262]='h00000fdc;  wr_data_rom[ 4262]='h000033e1;
    rd_cycle[ 4263] = 1'b0;  wr_cycle[ 4263] = 1'b1;  addr_rom[ 4263]='h000028c0;  wr_data_rom[ 4263]='h00000225;
    rd_cycle[ 4264] = 1'b1;  wr_cycle[ 4264] = 1'b0;  addr_rom[ 4264]='h00000d78;  wr_data_rom[ 4264]='h00000000;
    rd_cycle[ 4265] = 1'b1;  wr_cycle[ 4265] = 1'b0;  addr_rom[ 4265]='h000030dc;  wr_data_rom[ 4265]='h00000000;
    rd_cycle[ 4266] = 1'b1;  wr_cycle[ 4266] = 1'b0;  addr_rom[ 4266]='h00000fc0;  wr_data_rom[ 4266]='h00000000;
    rd_cycle[ 4267] = 1'b1;  wr_cycle[ 4267] = 1'b0;  addr_rom[ 4267]='h00003850;  wr_data_rom[ 4267]='h00000000;
    rd_cycle[ 4268] = 1'b1;  wr_cycle[ 4268] = 1'b0;  addr_rom[ 4268]='h00003844;  wr_data_rom[ 4268]='h00000000;
    rd_cycle[ 4269] = 1'b0;  wr_cycle[ 4269] = 1'b1;  addr_rom[ 4269]='h000013d8;  wr_data_rom[ 4269]='h00003954;
    rd_cycle[ 4270] = 1'b0;  wr_cycle[ 4270] = 1'b1;  addr_rom[ 4270]='h00002d84;  wr_data_rom[ 4270]='h00003b40;
    rd_cycle[ 4271] = 1'b0;  wr_cycle[ 4271] = 1'b1;  addr_rom[ 4271]='h00002cc4;  wr_data_rom[ 4271]='h000033b5;
    rd_cycle[ 4272] = 1'b1;  wr_cycle[ 4272] = 1'b0;  addr_rom[ 4272]='h00000214;  wr_data_rom[ 4272]='h00000000;
    rd_cycle[ 4273] = 1'b0;  wr_cycle[ 4273] = 1'b1;  addr_rom[ 4273]='h0000028c;  wr_data_rom[ 4273]='h00003784;
    rd_cycle[ 4274] = 1'b0;  wr_cycle[ 4274] = 1'b1;  addr_rom[ 4274]='h00003b10;  wr_data_rom[ 4274]='h00001eba;
    rd_cycle[ 4275] = 1'b1;  wr_cycle[ 4275] = 1'b0;  addr_rom[ 4275]='h00003d88;  wr_data_rom[ 4275]='h00000000;
    rd_cycle[ 4276] = 1'b1;  wr_cycle[ 4276] = 1'b0;  addr_rom[ 4276]='h00000fd0;  wr_data_rom[ 4276]='h00000000;
    rd_cycle[ 4277] = 1'b1;  wr_cycle[ 4277] = 1'b0;  addr_rom[ 4277]='h00000dc0;  wr_data_rom[ 4277]='h00000000;
    rd_cycle[ 4278] = 1'b0;  wr_cycle[ 4278] = 1'b1;  addr_rom[ 4278]='h00000b00;  wr_data_rom[ 4278]='h000019cc;
    rd_cycle[ 4279] = 1'b0;  wr_cycle[ 4279] = 1'b1;  addr_rom[ 4279]='h00002298;  wr_data_rom[ 4279]='h00000b9d;
    rd_cycle[ 4280] = 1'b0;  wr_cycle[ 4280] = 1'b1;  addr_rom[ 4280]='h00001e14;  wr_data_rom[ 4280]='h00003b12;
    rd_cycle[ 4281] = 1'b0;  wr_cycle[ 4281] = 1'b1;  addr_rom[ 4281]='h00000770;  wr_data_rom[ 4281]='h000033b9;
    rd_cycle[ 4282] = 1'b1;  wr_cycle[ 4282] = 1'b0;  addr_rom[ 4282]='h00000e84;  wr_data_rom[ 4282]='h00000000;
    rd_cycle[ 4283] = 1'b1;  wr_cycle[ 4283] = 1'b0;  addr_rom[ 4283]='h00001ab8;  wr_data_rom[ 4283]='h00000000;
    rd_cycle[ 4284] = 1'b0;  wr_cycle[ 4284] = 1'b1;  addr_rom[ 4284]='h00002820;  wr_data_rom[ 4284]='h0000012c;
    rd_cycle[ 4285] = 1'b0;  wr_cycle[ 4285] = 1'b1;  addr_rom[ 4285]='h00003d4c;  wr_data_rom[ 4285]='h00002fbc;
    rd_cycle[ 4286] = 1'b0;  wr_cycle[ 4286] = 1'b1;  addr_rom[ 4286]='h00001c8c;  wr_data_rom[ 4286]='h00000b10;
    rd_cycle[ 4287] = 1'b0;  wr_cycle[ 4287] = 1'b1;  addr_rom[ 4287]='h00002e88;  wr_data_rom[ 4287]='h000038ea;
    rd_cycle[ 4288] = 1'b1;  wr_cycle[ 4288] = 1'b0;  addr_rom[ 4288]='h000016ac;  wr_data_rom[ 4288]='h00000000;
    rd_cycle[ 4289] = 1'b1;  wr_cycle[ 4289] = 1'b0;  addr_rom[ 4289]='h00000868;  wr_data_rom[ 4289]='h00000000;
    rd_cycle[ 4290] = 1'b0;  wr_cycle[ 4290] = 1'b1;  addr_rom[ 4290]='h0000013c;  wr_data_rom[ 4290]='h00002414;
    rd_cycle[ 4291] = 1'b0;  wr_cycle[ 4291] = 1'b1;  addr_rom[ 4291]='h00002f3c;  wr_data_rom[ 4291]='h00001307;
    rd_cycle[ 4292] = 1'b1;  wr_cycle[ 4292] = 1'b0;  addr_rom[ 4292]='h00002060;  wr_data_rom[ 4292]='h00000000;
    rd_cycle[ 4293] = 1'b0;  wr_cycle[ 4293] = 1'b1;  addr_rom[ 4293]='h0000187c;  wr_data_rom[ 4293]='h00001fbe;
    rd_cycle[ 4294] = 1'b0;  wr_cycle[ 4294] = 1'b1;  addr_rom[ 4294]='h00002b18;  wr_data_rom[ 4294]='h0000223d;
    rd_cycle[ 4295] = 1'b0;  wr_cycle[ 4295] = 1'b1;  addr_rom[ 4295]='h0000313c;  wr_data_rom[ 4295]='h00003bdb;
    rd_cycle[ 4296] = 1'b0;  wr_cycle[ 4296] = 1'b1;  addr_rom[ 4296]='h00000c10;  wr_data_rom[ 4296]='h000016fe;
    rd_cycle[ 4297] = 1'b1;  wr_cycle[ 4297] = 1'b0;  addr_rom[ 4297]='h00000e30;  wr_data_rom[ 4297]='h00000000;
    rd_cycle[ 4298] = 1'b1;  wr_cycle[ 4298] = 1'b0;  addr_rom[ 4298]='h00001fe4;  wr_data_rom[ 4298]='h00000000;
    rd_cycle[ 4299] = 1'b1;  wr_cycle[ 4299] = 1'b0;  addr_rom[ 4299]='h000010f4;  wr_data_rom[ 4299]='h00000000;
    rd_cycle[ 4300] = 1'b0;  wr_cycle[ 4300] = 1'b1;  addr_rom[ 4300]='h00000304;  wr_data_rom[ 4300]='h000023e0;
    rd_cycle[ 4301] = 1'b1;  wr_cycle[ 4301] = 1'b0;  addr_rom[ 4301]='h000004b0;  wr_data_rom[ 4301]='h00000000;
    rd_cycle[ 4302] = 1'b1;  wr_cycle[ 4302] = 1'b0;  addr_rom[ 4302]='h00002078;  wr_data_rom[ 4302]='h00000000;
    rd_cycle[ 4303] = 1'b0;  wr_cycle[ 4303] = 1'b1;  addr_rom[ 4303]='h000021d8;  wr_data_rom[ 4303]='h00000c37;
    rd_cycle[ 4304] = 1'b1;  wr_cycle[ 4304] = 1'b0;  addr_rom[ 4304]='h000012b0;  wr_data_rom[ 4304]='h00000000;
    rd_cycle[ 4305] = 1'b1;  wr_cycle[ 4305] = 1'b0;  addr_rom[ 4305]='h000036a0;  wr_data_rom[ 4305]='h00000000;
    rd_cycle[ 4306] = 1'b1;  wr_cycle[ 4306] = 1'b0;  addr_rom[ 4306]='h00003fc4;  wr_data_rom[ 4306]='h00000000;
    rd_cycle[ 4307] = 1'b0;  wr_cycle[ 4307] = 1'b1;  addr_rom[ 4307]='h00003b2c;  wr_data_rom[ 4307]='h00002664;
    rd_cycle[ 4308] = 1'b0;  wr_cycle[ 4308] = 1'b1;  addr_rom[ 4308]='h000009f0;  wr_data_rom[ 4308]='h000020d8;
    rd_cycle[ 4309] = 1'b1;  wr_cycle[ 4309] = 1'b0;  addr_rom[ 4309]='h00002ad8;  wr_data_rom[ 4309]='h00000000;
    rd_cycle[ 4310] = 1'b1;  wr_cycle[ 4310] = 1'b0;  addr_rom[ 4310]='h000010d8;  wr_data_rom[ 4310]='h00000000;
    rd_cycle[ 4311] = 1'b0;  wr_cycle[ 4311] = 1'b1;  addr_rom[ 4311]='h000019dc;  wr_data_rom[ 4311]='h00003625;
    rd_cycle[ 4312] = 1'b0;  wr_cycle[ 4312] = 1'b1;  addr_rom[ 4312]='h00001940;  wr_data_rom[ 4312]='h00003867;
    rd_cycle[ 4313] = 1'b0;  wr_cycle[ 4313] = 1'b1;  addr_rom[ 4313]='h00000d68;  wr_data_rom[ 4313]='h0000313f;
    rd_cycle[ 4314] = 1'b0;  wr_cycle[ 4314] = 1'b1;  addr_rom[ 4314]='h00000e98;  wr_data_rom[ 4314]='h000002b7;
    rd_cycle[ 4315] = 1'b1;  wr_cycle[ 4315] = 1'b0;  addr_rom[ 4315]='h00002004;  wr_data_rom[ 4315]='h00000000;
    rd_cycle[ 4316] = 1'b1;  wr_cycle[ 4316] = 1'b0;  addr_rom[ 4316]='h00000168;  wr_data_rom[ 4316]='h00000000;
    rd_cycle[ 4317] = 1'b1;  wr_cycle[ 4317] = 1'b0;  addr_rom[ 4317]='h000018a0;  wr_data_rom[ 4317]='h00000000;
    rd_cycle[ 4318] = 1'b0;  wr_cycle[ 4318] = 1'b1;  addr_rom[ 4318]='h000034d8;  wr_data_rom[ 4318]='h00003707;
    rd_cycle[ 4319] = 1'b0;  wr_cycle[ 4319] = 1'b1;  addr_rom[ 4319]='h00003b7c;  wr_data_rom[ 4319]='h00001839;
    rd_cycle[ 4320] = 1'b0;  wr_cycle[ 4320] = 1'b1;  addr_rom[ 4320]='h00000eb4;  wr_data_rom[ 4320]='h0000347b;
    rd_cycle[ 4321] = 1'b0;  wr_cycle[ 4321] = 1'b1;  addr_rom[ 4321]='h000031a0;  wr_data_rom[ 4321]='h00001993;
    rd_cycle[ 4322] = 1'b0;  wr_cycle[ 4322] = 1'b1;  addr_rom[ 4322]='h00001ad8;  wr_data_rom[ 4322]='h00003993;
    rd_cycle[ 4323] = 1'b0;  wr_cycle[ 4323] = 1'b1;  addr_rom[ 4323]='h000015fc;  wr_data_rom[ 4323]='h00003d31;
    rd_cycle[ 4324] = 1'b1;  wr_cycle[ 4324] = 1'b0;  addr_rom[ 4324]='h00003cd0;  wr_data_rom[ 4324]='h00000000;
    rd_cycle[ 4325] = 1'b0;  wr_cycle[ 4325] = 1'b1;  addr_rom[ 4325]='h00000e94;  wr_data_rom[ 4325]='h000019b3;
    rd_cycle[ 4326] = 1'b1;  wr_cycle[ 4326] = 1'b0;  addr_rom[ 4326]='h000021ac;  wr_data_rom[ 4326]='h00000000;
    rd_cycle[ 4327] = 1'b0;  wr_cycle[ 4327] = 1'b1;  addr_rom[ 4327]='h00002dcc;  wr_data_rom[ 4327]='h00002897;
    rd_cycle[ 4328] = 1'b1;  wr_cycle[ 4328] = 1'b0;  addr_rom[ 4328]='h000024e4;  wr_data_rom[ 4328]='h00000000;
    rd_cycle[ 4329] = 1'b0;  wr_cycle[ 4329] = 1'b1;  addr_rom[ 4329]='h000015dc;  wr_data_rom[ 4329]='h00001529;
    rd_cycle[ 4330] = 1'b1;  wr_cycle[ 4330] = 1'b0;  addr_rom[ 4330]='h0000142c;  wr_data_rom[ 4330]='h00000000;
    rd_cycle[ 4331] = 1'b1;  wr_cycle[ 4331] = 1'b0;  addr_rom[ 4331]='h000039c0;  wr_data_rom[ 4331]='h00000000;
    rd_cycle[ 4332] = 1'b0;  wr_cycle[ 4332] = 1'b1;  addr_rom[ 4332]='h000016ac;  wr_data_rom[ 4332]='h00000c1a;
    rd_cycle[ 4333] = 1'b0;  wr_cycle[ 4333] = 1'b1;  addr_rom[ 4333]='h00001694;  wr_data_rom[ 4333]='h00002331;
    rd_cycle[ 4334] = 1'b0;  wr_cycle[ 4334] = 1'b1;  addr_rom[ 4334]='h000007d8;  wr_data_rom[ 4334]='h000003f0;
    rd_cycle[ 4335] = 1'b1;  wr_cycle[ 4335] = 1'b0;  addr_rom[ 4335]='h000012bc;  wr_data_rom[ 4335]='h00000000;
    rd_cycle[ 4336] = 1'b1;  wr_cycle[ 4336] = 1'b0;  addr_rom[ 4336]='h00000318;  wr_data_rom[ 4336]='h00000000;
    rd_cycle[ 4337] = 1'b0;  wr_cycle[ 4337] = 1'b1;  addr_rom[ 4337]='h00001b60;  wr_data_rom[ 4337]='h00001e6d;
    rd_cycle[ 4338] = 1'b1;  wr_cycle[ 4338] = 1'b0;  addr_rom[ 4338]='h00001180;  wr_data_rom[ 4338]='h00000000;
    rd_cycle[ 4339] = 1'b0;  wr_cycle[ 4339] = 1'b1;  addr_rom[ 4339]='h00002dc8;  wr_data_rom[ 4339]='h00002ea0;
    rd_cycle[ 4340] = 1'b0;  wr_cycle[ 4340] = 1'b1;  addr_rom[ 4340]='h00003ee0;  wr_data_rom[ 4340]='h0000023c;
    rd_cycle[ 4341] = 1'b1;  wr_cycle[ 4341] = 1'b0;  addr_rom[ 4341]='h00002af4;  wr_data_rom[ 4341]='h00000000;
    rd_cycle[ 4342] = 1'b0;  wr_cycle[ 4342] = 1'b1;  addr_rom[ 4342]='h00000360;  wr_data_rom[ 4342]='h00003c09;
    rd_cycle[ 4343] = 1'b1;  wr_cycle[ 4343] = 1'b0;  addr_rom[ 4343]='h00002030;  wr_data_rom[ 4343]='h00000000;
    rd_cycle[ 4344] = 1'b1;  wr_cycle[ 4344] = 1'b0;  addr_rom[ 4344]='h0000222c;  wr_data_rom[ 4344]='h00000000;
    rd_cycle[ 4345] = 1'b1;  wr_cycle[ 4345] = 1'b0;  addr_rom[ 4345]='h000019e8;  wr_data_rom[ 4345]='h00000000;
    rd_cycle[ 4346] = 1'b0;  wr_cycle[ 4346] = 1'b1;  addr_rom[ 4346]='h00002d7c;  wr_data_rom[ 4346]='h00001520;
    rd_cycle[ 4347] = 1'b0;  wr_cycle[ 4347] = 1'b1;  addr_rom[ 4347]='h00003e90;  wr_data_rom[ 4347]='h00001471;
    rd_cycle[ 4348] = 1'b1;  wr_cycle[ 4348] = 1'b0;  addr_rom[ 4348]='h00003250;  wr_data_rom[ 4348]='h00000000;
    rd_cycle[ 4349] = 1'b0;  wr_cycle[ 4349] = 1'b1;  addr_rom[ 4349]='h00002d44;  wr_data_rom[ 4349]='h000002d0;
    rd_cycle[ 4350] = 1'b1;  wr_cycle[ 4350] = 1'b0;  addr_rom[ 4350]='h000014f4;  wr_data_rom[ 4350]='h00000000;
    rd_cycle[ 4351] = 1'b1;  wr_cycle[ 4351] = 1'b0;  addr_rom[ 4351]='h00001690;  wr_data_rom[ 4351]='h00000000;
    rd_cycle[ 4352] = 1'b1;  wr_cycle[ 4352] = 1'b0;  addr_rom[ 4352]='h00000c40;  wr_data_rom[ 4352]='h00000000;
    rd_cycle[ 4353] = 1'b1;  wr_cycle[ 4353] = 1'b0;  addr_rom[ 4353]='h00002b6c;  wr_data_rom[ 4353]='h00000000;
    rd_cycle[ 4354] = 1'b0;  wr_cycle[ 4354] = 1'b1;  addr_rom[ 4354]='h000002b8;  wr_data_rom[ 4354]='h00002d04;
    rd_cycle[ 4355] = 1'b1;  wr_cycle[ 4355] = 1'b0;  addr_rom[ 4355]='h00003954;  wr_data_rom[ 4355]='h00000000;
    rd_cycle[ 4356] = 1'b1;  wr_cycle[ 4356] = 1'b0;  addr_rom[ 4356]='h00001888;  wr_data_rom[ 4356]='h00000000;
    rd_cycle[ 4357] = 1'b0;  wr_cycle[ 4357] = 1'b1;  addr_rom[ 4357]='h00001128;  wr_data_rom[ 4357]='h00002b50;
    rd_cycle[ 4358] = 1'b1;  wr_cycle[ 4358] = 1'b0;  addr_rom[ 4358]='h0000245c;  wr_data_rom[ 4358]='h00000000;
    rd_cycle[ 4359] = 1'b0;  wr_cycle[ 4359] = 1'b1;  addr_rom[ 4359]='h0000103c;  wr_data_rom[ 4359]='h0000011b;
    rd_cycle[ 4360] = 1'b0;  wr_cycle[ 4360] = 1'b1;  addr_rom[ 4360]='h00002e20;  wr_data_rom[ 4360]='h000018e7;
    rd_cycle[ 4361] = 1'b1;  wr_cycle[ 4361] = 1'b0;  addr_rom[ 4361]='h000007ac;  wr_data_rom[ 4361]='h00000000;
    rd_cycle[ 4362] = 1'b0;  wr_cycle[ 4362] = 1'b1;  addr_rom[ 4362]='h00001fbc;  wr_data_rom[ 4362]='h00001c05;
    rd_cycle[ 4363] = 1'b1;  wr_cycle[ 4363] = 1'b0;  addr_rom[ 4363]='h000017ec;  wr_data_rom[ 4363]='h00000000;
    rd_cycle[ 4364] = 1'b0;  wr_cycle[ 4364] = 1'b1;  addr_rom[ 4364]='h00001218;  wr_data_rom[ 4364]='h00000094;
    rd_cycle[ 4365] = 1'b0;  wr_cycle[ 4365] = 1'b1;  addr_rom[ 4365]='h000012b0;  wr_data_rom[ 4365]='h00002562;
    rd_cycle[ 4366] = 1'b1;  wr_cycle[ 4366] = 1'b0;  addr_rom[ 4366]='h00003074;  wr_data_rom[ 4366]='h00000000;
    rd_cycle[ 4367] = 1'b0;  wr_cycle[ 4367] = 1'b1;  addr_rom[ 4367]='h00001a08;  wr_data_rom[ 4367]='h0000196b;
    rd_cycle[ 4368] = 1'b0;  wr_cycle[ 4368] = 1'b1;  addr_rom[ 4368]='h00002f7c;  wr_data_rom[ 4368]='h00000118;
    rd_cycle[ 4369] = 1'b1;  wr_cycle[ 4369] = 1'b0;  addr_rom[ 4369]='h00001f88;  wr_data_rom[ 4369]='h00000000;
    rd_cycle[ 4370] = 1'b1;  wr_cycle[ 4370] = 1'b0;  addr_rom[ 4370]='h00000a98;  wr_data_rom[ 4370]='h00000000;
    rd_cycle[ 4371] = 1'b1;  wr_cycle[ 4371] = 1'b0;  addr_rom[ 4371]='h00001428;  wr_data_rom[ 4371]='h00000000;
    rd_cycle[ 4372] = 1'b0;  wr_cycle[ 4372] = 1'b1;  addr_rom[ 4372]='h00001490;  wr_data_rom[ 4372]='h00003561;
    rd_cycle[ 4373] = 1'b0;  wr_cycle[ 4373] = 1'b1;  addr_rom[ 4373]='h00003f9c;  wr_data_rom[ 4373]='h00000fd0;
    rd_cycle[ 4374] = 1'b0;  wr_cycle[ 4374] = 1'b1;  addr_rom[ 4374]='h00003f38;  wr_data_rom[ 4374]='h00000cb0;
    rd_cycle[ 4375] = 1'b0;  wr_cycle[ 4375] = 1'b1;  addr_rom[ 4375]='h00003358;  wr_data_rom[ 4375]='h000035e4;
    rd_cycle[ 4376] = 1'b1;  wr_cycle[ 4376] = 1'b0;  addr_rom[ 4376]='h000038b0;  wr_data_rom[ 4376]='h00000000;
    rd_cycle[ 4377] = 1'b1;  wr_cycle[ 4377] = 1'b0;  addr_rom[ 4377]='h00001360;  wr_data_rom[ 4377]='h00000000;
    rd_cycle[ 4378] = 1'b1;  wr_cycle[ 4378] = 1'b0;  addr_rom[ 4378]='h00002818;  wr_data_rom[ 4378]='h00000000;
    rd_cycle[ 4379] = 1'b0;  wr_cycle[ 4379] = 1'b1;  addr_rom[ 4379]='h00001e64;  wr_data_rom[ 4379]='h0000397d;
    rd_cycle[ 4380] = 1'b1;  wr_cycle[ 4380] = 1'b0;  addr_rom[ 4380]='h00003a58;  wr_data_rom[ 4380]='h00000000;
    rd_cycle[ 4381] = 1'b0;  wr_cycle[ 4381] = 1'b1;  addr_rom[ 4381]='h00000b8c;  wr_data_rom[ 4381]='h00002348;
    rd_cycle[ 4382] = 1'b0;  wr_cycle[ 4382] = 1'b1;  addr_rom[ 4382]='h000003a0;  wr_data_rom[ 4382]='h00000a97;
    rd_cycle[ 4383] = 1'b1;  wr_cycle[ 4383] = 1'b0;  addr_rom[ 4383]='h000014e4;  wr_data_rom[ 4383]='h00000000;
    rd_cycle[ 4384] = 1'b0;  wr_cycle[ 4384] = 1'b1;  addr_rom[ 4384]='h00002504;  wr_data_rom[ 4384]='h00001ed7;
    rd_cycle[ 4385] = 1'b1;  wr_cycle[ 4385] = 1'b0;  addr_rom[ 4385]='h00003210;  wr_data_rom[ 4385]='h00000000;
    rd_cycle[ 4386] = 1'b0;  wr_cycle[ 4386] = 1'b1;  addr_rom[ 4386]='h000006fc;  wr_data_rom[ 4386]='h00002487;
    rd_cycle[ 4387] = 1'b0;  wr_cycle[ 4387] = 1'b1;  addr_rom[ 4387]='h000029f0;  wr_data_rom[ 4387]='h00001120;
    rd_cycle[ 4388] = 1'b0;  wr_cycle[ 4388] = 1'b1;  addr_rom[ 4388]='h000001c4;  wr_data_rom[ 4388]='h00003298;
    rd_cycle[ 4389] = 1'b1;  wr_cycle[ 4389] = 1'b0;  addr_rom[ 4389]='h00000a18;  wr_data_rom[ 4389]='h00000000;
    rd_cycle[ 4390] = 1'b0;  wr_cycle[ 4390] = 1'b1;  addr_rom[ 4390]='h00003c40;  wr_data_rom[ 4390]='h00001666;
    rd_cycle[ 4391] = 1'b0;  wr_cycle[ 4391] = 1'b1;  addr_rom[ 4391]='h00001f60;  wr_data_rom[ 4391]='h000010c0;
    rd_cycle[ 4392] = 1'b1;  wr_cycle[ 4392] = 1'b0;  addr_rom[ 4392]='h0000297c;  wr_data_rom[ 4392]='h00000000;
    rd_cycle[ 4393] = 1'b0;  wr_cycle[ 4393] = 1'b1;  addr_rom[ 4393]='h00001eec;  wr_data_rom[ 4393]='h00002cb3;
    rd_cycle[ 4394] = 1'b0;  wr_cycle[ 4394] = 1'b1;  addr_rom[ 4394]='h0000294c;  wr_data_rom[ 4394]='h00003dee;
    rd_cycle[ 4395] = 1'b0;  wr_cycle[ 4395] = 1'b1;  addr_rom[ 4395]='h00002d5c;  wr_data_rom[ 4395]='h0000018e;
    rd_cycle[ 4396] = 1'b1;  wr_cycle[ 4396] = 1'b0;  addr_rom[ 4396]='h00001380;  wr_data_rom[ 4396]='h00000000;
    rd_cycle[ 4397] = 1'b0;  wr_cycle[ 4397] = 1'b1;  addr_rom[ 4397]='h00003e70;  wr_data_rom[ 4397]='h00003371;
    rd_cycle[ 4398] = 1'b0;  wr_cycle[ 4398] = 1'b1;  addr_rom[ 4398]='h00002e00;  wr_data_rom[ 4398]='h00002d09;
    rd_cycle[ 4399] = 1'b1;  wr_cycle[ 4399] = 1'b0;  addr_rom[ 4399]='h000033d4;  wr_data_rom[ 4399]='h00000000;
    rd_cycle[ 4400] = 1'b1;  wr_cycle[ 4400] = 1'b0;  addr_rom[ 4400]='h00000704;  wr_data_rom[ 4400]='h00000000;
    rd_cycle[ 4401] = 1'b0;  wr_cycle[ 4401] = 1'b1;  addr_rom[ 4401]='h00002cf0;  wr_data_rom[ 4401]='h000026d7;
    rd_cycle[ 4402] = 1'b1;  wr_cycle[ 4402] = 1'b0;  addr_rom[ 4402]='h00003d54;  wr_data_rom[ 4402]='h00000000;
    rd_cycle[ 4403] = 1'b0;  wr_cycle[ 4403] = 1'b1;  addr_rom[ 4403]='h00002d74;  wr_data_rom[ 4403]='h00002858;
    rd_cycle[ 4404] = 1'b0;  wr_cycle[ 4404] = 1'b1;  addr_rom[ 4404]='h000020bc;  wr_data_rom[ 4404]='h00001927;
    rd_cycle[ 4405] = 1'b0;  wr_cycle[ 4405] = 1'b1;  addr_rom[ 4405]='h00001c5c;  wr_data_rom[ 4405]='h00000415;
    rd_cycle[ 4406] = 1'b0;  wr_cycle[ 4406] = 1'b1;  addr_rom[ 4406]='h00002750;  wr_data_rom[ 4406]='h00000b46;
    rd_cycle[ 4407] = 1'b1;  wr_cycle[ 4407] = 1'b0;  addr_rom[ 4407]='h0000371c;  wr_data_rom[ 4407]='h00000000;
    rd_cycle[ 4408] = 1'b1;  wr_cycle[ 4408] = 1'b0;  addr_rom[ 4408]='h000028cc;  wr_data_rom[ 4408]='h00000000;
    rd_cycle[ 4409] = 1'b1;  wr_cycle[ 4409] = 1'b0;  addr_rom[ 4409]='h00002c88;  wr_data_rom[ 4409]='h00000000;
    rd_cycle[ 4410] = 1'b0;  wr_cycle[ 4410] = 1'b1;  addr_rom[ 4410]='h000036e8;  wr_data_rom[ 4410]='h0000054b;
    rd_cycle[ 4411] = 1'b1;  wr_cycle[ 4411] = 1'b0;  addr_rom[ 4411]='h000022dc;  wr_data_rom[ 4411]='h00000000;
    rd_cycle[ 4412] = 1'b0;  wr_cycle[ 4412] = 1'b1;  addr_rom[ 4412]='h00000fec;  wr_data_rom[ 4412]='h000018de;
    rd_cycle[ 4413] = 1'b1;  wr_cycle[ 4413] = 1'b0;  addr_rom[ 4413]='h00000554;  wr_data_rom[ 4413]='h00000000;
    rd_cycle[ 4414] = 1'b1;  wr_cycle[ 4414] = 1'b0;  addr_rom[ 4414]='h00003d04;  wr_data_rom[ 4414]='h00000000;
    rd_cycle[ 4415] = 1'b1;  wr_cycle[ 4415] = 1'b0;  addr_rom[ 4415]='h00003f78;  wr_data_rom[ 4415]='h00000000;
    rd_cycle[ 4416] = 1'b1;  wr_cycle[ 4416] = 1'b0;  addr_rom[ 4416]='h00003b24;  wr_data_rom[ 4416]='h00000000;
    rd_cycle[ 4417] = 1'b0;  wr_cycle[ 4417] = 1'b1;  addr_rom[ 4417]='h000039e8;  wr_data_rom[ 4417]='h00001cf4;
    rd_cycle[ 4418] = 1'b1;  wr_cycle[ 4418] = 1'b0;  addr_rom[ 4418]='h000016a4;  wr_data_rom[ 4418]='h00000000;
    rd_cycle[ 4419] = 1'b0;  wr_cycle[ 4419] = 1'b1;  addr_rom[ 4419]='h00001348;  wr_data_rom[ 4419]='h00003cd0;
    rd_cycle[ 4420] = 1'b0;  wr_cycle[ 4420] = 1'b1;  addr_rom[ 4420]='h000000f0;  wr_data_rom[ 4420]='h00000656;
    rd_cycle[ 4421] = 1'b1;  wr_cycle[ 4421] = 1'b0;  addr_rom[ 4421]='h0000293c;  wr_data_rom[ 4421]='h00000000;
    rd_cycle[ 4422] = 1'b0;  wr_cycle[ 4422] = 1'b1;  addr_rom[ 4422]='h00000794;  wr_data_rom[ 4422]='h000009d9;
    rd_cycle[ 4423] = 1'b1;  wr_cycle[ 4423] = 1'b0;  addr_rom[ 4423]='h00003a38;  wr_data_rom[ 4423]='h00000000;
    rd_cycle[ 4424] = 1'b1;  wr_cycle[ 4424] = 1'b0;  addr_rom[ 4424]='h0000297c;  wr_data_rom[ 4424]='h00000000;
    rd_cycle[ 4425] = 1'b0;  wr_cycle[ 4425] = 1'b1;  addr_rom[ 4425]='h0000210c;  wr_data_rom[ 4425]='h00000ff2;
    rd_cycle[ 4426] = 1'b1;  wr_cycle[ 4426] = 1'b0;  addr_rom[ 4426]='h00003c48;  wr_data_rom[ 4426]='h00000000;
    rd_cycle[ 4427] = 1'b0;  wr_cycle[ 4427] = 1'b1;  addr_rom[ 4427]='h00002bd8;  wr_data_rom[ 4427]='h00000c90;
    rd_cycle[ 4428] = 1'b0;  wr_cycle[ 4428] = 1'b1;  addr_rom[ 4428]='h00002c64;  wr_data_rom[ 4428]='h000014a3;
    rd_cycle[ 4429] = 1'b0;  wr_cycle[ 4429] = 1'b1;  addr_rom[ 4429]='h000029ec;  wr_data_rom[ 4429]='h00002dad;
    rd_cycle[ 4430] = 1'b1;  wr_cycle[ 4430] = 1'b0;  addr_rom[ 4430]='h00002a48;  wr_data_rom[ 4430]='h00000000;
    rd_cycle[ 4431] = 1'b0;  wr_cycle[ 4431] = 1'b1;  addr_rom[ 4431]='h00002ea8;  wr_data_rom[ 4431]='h000002b2;
    rd_cycle[ 4432] = 1'b0;  wr_cycle[ 4432] = 1'b1;  addr_rom[ 4432]='h00000ad4;  wr_data_rom[ 4432]='h0000158c;
    rd_cycle[ 4433] = 1'b0;  wr_cycle[ 4433] = 1'b1;  addr_rom[ 4433]='h00003914;  wr_data_rom[ 4433]='h00000de3;
    rd_cycle[ 4434] = 1'b0;  wr_cycle[ 4434] = 1'b1;  addr_rom[ 4434]='h000007b0;  wr_data_rom[ 4434]='h00003150;
    rd_cycle[ 4435] = 1'b1;  wr_cycle[ 4435] = 1'b0;  addr_rom[ 4435]='h000038a8;  wr_data_rom[ 4435]='h00000000;
    rd_cycle[ 4436] = 1'b0;  wr_cycle[ 4436] = 1'b1;  addr_rom[ 4436]='h00002a5c;  wr_data_rom[ 4436]='h00000ccc;
    rd_cycle[ 4437] = 1'b1;  wr_cycle[ 4437] = 1'b0;  addr_rom[ 4437]='h00000cfc;  wr_data_rom[ 4437]='h00000000;
    rd_cycle[ 4438] = 1'b0;  wr_cycle[ 4438] = 1'b1;  addr_rom[ 4438]='h00003ef8;  wr_data_rom[ 4438]='h00000863;
    rd_cycle[ 4439] = 1'b0;  wr_cycle[ 4439] = 1'b1;  addr_rom[ 4439]='h00002dd0;  wr_data_rom[ 4439]='h00001b99;
    rd_cycle[ 4440] = 1'b1;  wr_cycle[ 4440] = 1'b0;  addr_rom[ 4440]='h00003adc;  wr_data_rom[ 4440]='h00000000;
    rd_cycle[ 4441] = 1'b1;  wr_cycle[ 4441] = 1'b0;  addr_rom[ 4441]='h000012f4;  wr_data_rom[ 4441]='h00000000;
    rd_cycle[ 4442] = 1'b1;  wr_cycle[ 4442] = 1'b0;  addr_rom[ 4442]='h00002570;  wr_data_rom[ 4442]='h00000000;
    rd_cycle[ 4443] = 1'b0;  wr_cycle[ 4443] = 1'b1;  addr_rom[ 4443]='h00002b98;  wr_data_rom[ 4443]='h00003c0b;
    rd_cycle[ 4444] = 1'b1;  wr_cycle[ 4444] = 1'b0;  addr_rom[ 4444]='h00001410;  wr_data_rom[ 4444]='h00000000;
    rd_cycle[ 4445] = 1'b0;  wr_cycle[ 4445] = 1'b1;  addr_rom[ 4445]='h00002f60;  wr_data_rom[ 4445]='h00000764;
    rd_cycle[ 4446] = 1'b0;  wr_cycle[ 4446] = 1'b1;  addr_rom[ 4446]='h000032cc;  wr_data_rom[ 4446]='h00002ec5;
    rd_cycle[ 4447] = 1'b0;  wr_cycle[ 4447] = 1'b1;  addr_rom[ 4447]='h00003268;  wr_data_rom[ 4447]='h0000073e;
    rd_cycle[ 4448] = 1'b0;  wr_cycle[ 4448] = 1'b1;  addr_rom[ 4448]='h00000214;  wr_data_rom[ 4448]='h000014db;
    rd_cycle[ 4449] = 1'b0;  wr_cycle[ 4449] = 1'b1;  addr_rom[ 4449]='h00002594;  wr_data_rom[ 4449]='h00000b50;
    rd_cycle[ 4450] = 1'b0;  wr_cycle[ 4450] = 1'b1;  addr_rom[ 4450]='h00001060;  wr_data_rom[ 4450]='h00003d0f;
    rd_cycle[ 4451] = 1'b1;  wr_cycle[ 4451] = 1'b0;  addr_rom[ 4451]='h0000184c;  wr_data_rom[ 4451]='h00000000;
    rd_cycle[ 4452] = 1'b0;  wr_cycle[ 4452] = 1'b1;  addr_rom[ 4452]='h000035b0;  wr_data_rom[ 4452]='h0000195c;
    rd_cycle[ 4453] = 1'b0;  wr_cycle[ 4453] = 1'b1;  addr_rom[ 4453]='h00002368;  wr_data_rom[ 4453]='h00001c65;
    rd_cycle[ 4454] = 1'b0;  wr_cycle[ 4454] = 1'b1;  addr_rom[ 4454]='h0000022c;  wr_data_rom[ 4454]='h000012e2;
    rd_cycle[ 4455] = 1'b0;  wr_cycle[ 4455] = 1'b1;  addr_rom[ 4455]='h00001924;  wr_data_rom[ 4455]='h00001ce3;
    rd_cycle[ 4456] = 1'b1;  wr_cycle[ 4456] = 1'b0;  addr_rom[ 4456]='h00000328;  wr_data_rom[ 4456]='h00000000;
    rd_cycle[ 4457] = 1'b0;  wr_cycle[ 4457] = 1'b1;  addr_rom[ 4457]='h00000fd8;  wr_data_rom[ 4457]='h00001f0d;
    rd_cycle[ 4458] = 1'b0;  wr_cycle[ 4458] = 1'b1;  addr_rom[ 4458]='h000031b8;  wr_data_rom[ 4458]='h000022e7;
    rd_cycle[ 4459] = 1'b1;  wr_cycle[ 4459] = 1'b0;  addr_rom[ 4459]='h000001d0;  wr_data_rom[ 4459]='h00000000;
    rd_cycle[ 4460] = 1'b1;  wr_cycle[ 4460] = 1'b0;  addr_rom[ 4460]='h00001c7c;  wr_data_rom[ 4460]='h00000000;
    rd_cycle[ 4461] = 1'b0;  wr_cycle[ 4461] = 1'b1;  addr_rom[ 4461]='h00003b30;  wr_data_rom[ 4461]='h00001f6a;
    rd_cycle[ 4462] = 1'b0;  wr_cycle[ 4462] = 1'b1;  addr_rom[ 4462]='h00001090;  wr_data_rom[ 4462]='h00002188;
    rd_cycle[ 4463] = 1'b1;  wr_cycle[ 4463] = 1'b0;  addr_rom[ 4463]='h000015e4;  wr_data_rom[ 4463]='h00000000;
    rd_cycle[ 4464] = 1'b1;  wr_cycle[ 4464] = 1'b0;  addr_rom[ 4464]='h00000a04;  wr_data_rom[ 4464]='h00000000;
    rd_cycle[ 4465] = 1'b0;  wr_cycle[ 4465] = 1'b1;  addr_rom[ 4465]='h000020c8;  wr_data_rom[ 4465]='h00000688;
    rd_cycle[ 4466] = 1'b0;  wr_cycle[ 4466] = 1'b1;  addr_rom[ 4466]='h00001f8c;  wr_data_rom[ 4466]='h00001d9d;
    rd_cycle[ 4467] = 1'b1;  wr_cycle[ 4467] = 1'b0;  addr_rom[ 4467]='h0000218c;  wr_data_rom[ 4467]='h00000000;
    rd_cycle[ 4468] = 1'b1;  wr_cycle[ 4468] = 1'b0;  addr_rom[ 4468]='h000034d4;  wr_data_rom[ 4468]='h00000000;
    rd_cycle[ 4469] = 1'b0;  wr_cycle[ 4469] = 1'b1;  addr_rom[ 4469]='h000021f0;  wr_data_rom[ 4469]='h00003af4;
    rd_cycle[ 4470] = 1'b1;  wr_cycle[ 4470] = 1'b0;  addr_rom[ 4470]='h0000205c;  wr_data_rom[ 4470]='h00000000;
    rd_cycle[ 4471] = 1'b0;  wr_cycle[ 4471] = 1'b1;  addr_rom[ 4471]='h0000032c;  wr_data_rom[ 4471]='h00000a0a;
    rd_cycle[ 4472] = 1'b1;  wr_cycle[ 4472] = 1'b0;  addr_rom[ 4472]='h000030bc;  wr_data_rom[ 4472]='h00000000;
    rd_cycle[ 4473] = 1'b0;  wr_cycle[ 4473] = 1'b1;  addr_rom[ 4473]='h00003f7c;  wr_data_rom[ 4473]='h00002583;
    rd_cycle[ 4474] = 1'b1;  wr_cycle[ 4474] = 1'b0;  addr_rom[ 4474]='h000038cc;  wr_data_rom[ 4474]='h00000000;
    rd_cycle[ 4475] = 1'b0;  wr_cycle[ 4475] = 1'b1;  addr_rom[ 4475]='h00000d48;  wr_data_rom[ 4475]='h00003841;
    rd_cycle[ 4476] = 1'b0;  wr_cycle[ 4476] = 1'b1;  addr_rom[ 4476]='h00001cec;  wr_data_rom[ 4476]='h000017e7;
    rd_cycle[ 4477] = 1'b0;  wr_cycle[ 4477] = 1'b1;  addr_rom[ 4477]='h00000698;  wr_data_rom[ 4477]='h00001a77;
    rd_cycle[ 4478] = 1'b0;  wr_cycle[ 4478] = 1'b1;  addr_rom[ 4478]='h00000968;  wr_data_rom[ 4478]='h00003753;
    rd_cycle[ 4479] = 1'b1;  wr_cycle[ 4479] = 1'b0;  addr_rom[ 4479]='h000007d4;  wr_data_rom[ 4479]='h00000000;
    rd_cycle[ 4480] = 1'b0;  wr_cycle[ 4480] = 1'b1;  addr_rom[ 4480]='h000013a4;  wr_data_rom[ 4480]='h000032c0;
    rd_cycle[ 4481] = 1'b0;  wr_cycle[ 4481] = 1'b1;  addr_rom[ 4481]='h000016c4;  wr_data_rom[ 4481]='h00003870;
    rd_cycle[ 4482] = 1'b1;  wr_cycle[ 4482] = 1'b0;  addr_rom[ 4482]='h00001bf8;  wr_data_rom[ 4482]='h00000000;
    rd_cycle[ 4483] = 1'b0;  wr_cycle[ 4483] = 1'b1;  addr_rom[ 4483]='h00001958;  wr_data_rom[ 4483]='h0000142b;
    rd_cycle[ 4484] = 1'b0;  wr_cycle[ 4484] = 1'b1;  addr_rom[ 4484]='h00002b7c;  wr_data_rom[ 4484]='h0000191c;
    rd_cycle[ 4485] = 1'b0;  wr_cycle[ 4485] = 1'b1;  addr_rom[ 4485]='h00003488;  wr_data_rom[ 4485]='h0000264f;
    rd_cycle[ 4486] = 1'b1;  wr_cycle[ 4486] = 1'b0;  addr_rom[ 4486]='h00001d84;  wr_data_rom[ 4486]='h00000000;
    rd_cycle[ 4487] = 1'b1;  wr_cycle[ 4487] = 1'b0;  addr_rom[ 4487]='h000015f4;  wr_data_rom[ 4487]='h00000000;
    rd_cycle[ 4488] = 1'b1;  wr_cycle[ 4488] = 1'b0;  addr_rom[ 4488]='h00000228;  wr_data_rom[ 4488]='h00000000;
    rd_cycle[ 4489] = 1'b1;  wr_cycle[ 4489] = 1'b0;  addr_rom[ 4489]='h000001b4;  wr_data_rom[ 4489]='h00000000;
    rd_cycle[ 4490] = 1'b1;  wr_cycle[ 4490] = 1'b0;  addr_rom[ 4490]='h00003714;  wr_data_rom[ 4490]='h00000000;
    rd_cycle[ 4491] = 1'b1;  wr_cycle[ 4491] = 1'b0;  addr_rom[ 4491]='h000015a0;  wr_data_rom[ 4491]='h00000000;
    rd_cycle[ 4492] = 1'b0;  wr_cycle[ 4492] = 1'b1;  addr_rom[ 4492]='h0000395c;  wr_data_rom[ 4492]='h00001e84;
    rd_cycle[ 4493] = 1'b0;  wr_cycle[ 4493] = 1'b1;  addr_rom[ 4493]='h000035a0;  wr_data_rom[ 4493]='h00000423;
    rd_cycle[ 4494] = 1'b1;  wr_cycle[ 4494] = 1'b0;  addr_rom[ 4494]='h000026f4;  wr_data_rom[ 4494]='h00000000;
    rd_cycle[ 4495] = 1'b0;  wr_cycle[ 4495] = 1'b1;  addr_rom[ 4495]='h00002570;  wr_data_rom[ 4495]='h00000563;
    rd_cycle[ 4496] = 1'b1;  wr_cycle[ 4496] = 1'b0;  addr_rom[ 4496]='h00001610;  wr_data_rom[ 4496]='h00000000;
    rd_cycle[ 4497] = 1'b1;  wr_cycle[ 4497] = 1'b0;  addr_rom[ 4497]='h00002228;  wr_data_rom[ 4497]='h00000000;
    rd_cycle[ 4498] = 1'b1;  wr_cycle[ 4498] = 1'b0;  addr_rom[ 4498]='h00001934;  wr_data_rom[ 4498]='h00000000;
    rd_cycle[ 4499] = 1'b1;  wr_cycle[ 4499] = 1'b0;  addr_rom[ 4499]='h00002238;  wr_data_rom[ 4499]='h00000000;
    rd_cycle[ 4500] = 1'b1;  wr_cycle[ 4500] = 1'b0;  addr_rom[ 4500]='h000014fc;  wr_data_rom[ 4500]='h00000000;
    rd_cycle[ 4501] = 1'b0;  wr_cycle[ 4501] = 1'b1;  addr_rom[ 4501]='h000038a4;  wr_data_rom[ 4501]='h00002a1d;
    rd_cycle[ 4502] = 1'b1;  wr_cycle[ 4502] = 1'b0;  addr_rom[ 4502]='h00002244;  wr_data_rom[ 4502]='h00000000;
    rd_cycle[ 4503] = 1'b0;  wr_cycle[ 4503] = 1'b1;  addr_rom[ 4503]='h00000088;  wr_data_rom[ 4503]='h00002e75;
    rd_cycle[ 4504] = 1'b1;  wr_cycle[ 4504] = 1'b0;  addr_rom[ 4504]='h0000341c;  wr_data_rom[ 4504]='h00000000;
    rd_cycle[ 4505] = 1'b0;  wr_cycle[ 4505] = 1'b1;  addr_rom[ 4505]='h00003944;  wr_data_rom[ 4505]='h00003925;
    rd_cycle[ 4506] = 1'b1;  wr_cycle[ 4506] = 1'b0;  addr_rom[ 4506]='h00001ce0;  wr_data_rom[ 4506]='h00000000;
    rd_cycle[ 4507] = 1'b0;  wr_cycle[ 4507] = 1'b1;  addr_rom[ 4507]='h00002e80;  wr_data_rom[ 4507]='h00001a1d;
    rd_cycle[ 4508] = 1'b1;  wr_cycle[ 4508] = 1'b0;  addr_rom[ 4508]='h0000148c;  wr_data_rom[ 4508]='h00000000;
    rd_cycle[ 4509] = 1'b0;  wr_cycle[ 4509] = 1'b1;  addr_rom[ 4509]='h00000f14;  wr_data_rom[ 4509]='h00002db4;
    rd_cycle[ 4510] = 1'b1;  wr_cycle[ 4510] = 1'b0;  addr_rom[ 4510]='h00001d3c;  wr_data_rom[ 4510]='h00000000;
    rd_cycle[ 4511] = 1'b1;  wr_cycle[ 4511] = 1'b0;  addr_rom[ 4511]='h00000dc0;  wr_data_rom[ 4511]='h00000000;
    rd_cycle[ 4512] = 1'b1;  wr_cycle[ 4512] = 1'b0;  addr_rom[ 4512]='h00003374;  wr_data_rom[ 4512]='h00000000;
    rd_cycle[ 4513] = 1'b0;  wr_cycle[ 4513] = 1'b1;  addr_rom[ 4513]='h00003ef4;  wr_data_rom[ 4513]='h00000904;
    rd_cycle[ 4514] = 1'b0;  wr_cycle[ 4514] = 1'b1;  addr_rom[ 4514]='h00000914;  wr_data_rom[ 4514]='h00003f8b;
    rd_cycle[ 4515] = 1'b0;  wr_cycle[ 4515] = 1'b1;  addr_rom[ 4515]='h0000241c;  wr_data_rom[ 4515]='h000021e1;
    rd_cycle[ 4516] = 1'b0;  wr_cycle[ 4516] = 1'b1;  addr_rom[ 4516]='h00001050;  wr_data_rom[ 4516]='h00003ad3;
    rd_cycle[ 4517] = 1'b1;  wr_cycle[ 4517] = 1'b0;  addr_rom[ 4517]='h0000049c;  wr_data_rom[ 4517]='h00000000;
    rd_cycle[ 4518] = 1'b0;  wr_cycle[ 4518] = 1'b1;  addr_rom[ 4518]='h00000650;  wr_data_rom[ 4518]='h00003b14;
    rd_cycle[ 4519] = 1'b0;  wr_cycle[ 4519] = 1'b1;  addr_rom[ 4519]='h00000738;  wr_data_rom[ 4519]='h00001048;
    rd_cycle[ 4520] = 1'b1;  wr_cycle[ 4520] = 1'b0;  addr_rom[ 4520]='h00002180;  wr_data_rom[ 4520]='h00000000;
    rd_cycle[ 4521] = 1'b0;  wr_cycle[ 4521] = 1'b1;  addr_rom[ 4521]='h00002cac;  wr_data_rom[ 4521]='h000008de;
    rd_cycle[ 4522] = 1'b0;  wr_cycle[ 4522] = 1'b1;  addr_rom[ 4522]='h0000090c;  wr_data_rom[ 4522]='h00000998;
    rd_cycle[ 4523] = 1'b1;  wr_cycle[ 4523] = 1'b0;  addr_rom[ 4523]='h00003dcc;  wr_data_rom[ 4523]='h00000000;
    rd_cycle[ 4524] = 1'b0;  wr_cycle[ 4524] = 1'b1;  addr_rom[ 4524]='h000018fc;  wr_data_rom[ 4524]='h000028ee;
    rd_cycle[ 4525] = 1'b1;  wr_cycle[ 4525] = 1'b0;  addr_rom[ 4525]='h000020c8;  wr_data_rom[ 4525]='h00000000;
    rd_cycle[ 4526] = 1'b0;  wr_cycle[ 4526] = 1'b1;  addr_rom[ 4526]='h000023f4;  wr_data_rom[ 4526]='h0000023b;
    rd_cycle[ 4527] = 1'b0;  wr_cycle[ 4527] = 1'b1;  addr_rom[ 4527]='h00000bf0;  wr_data_rom[ 4527]='h00003ed0;
    rd_cycle[ 4528] = 1'b1;  wr_cycle[ 4528] = 1'b0;  addr_rom[ 4528]='h00003280;  wr_data_rom[ 4528]='h00000000;
    rd_cycle[ 4529] = 1'b1;  wr_cycle[ 4529] = 1'b0;  addr_rom[ 4529]='h00002ec0;  wr_data_rom[ 4529]='h00000000;
    rd_cycle[ 4530] = 1'b1;  wr_cycle[ 4530] = 1'b0;  addr_rom[ 4530]='h00003bc4;  wr_data_rom[ 4530]='h00000000;
    rd_cycle[ 4531] = 1'b1;  wr_cycle[ 4531] = 1'b0;  addr_rom[ 4531]='h000005fc;  wr_data_rom[ 4531]='h00000000;
    rd_cycle[ 4532] = 1'b0;  wr_cycle[ 4532] = 1'b1;  addr_rom[ 4532]='h0000306c;  wr_data_rom[ 4532]='h0000131b;
    rd_cycle[ 4533] = 1'b1;  wr_cycle[ 4533] = 1'b0;  addr_rom[ 4533]='h000037f0;  wr_data_rom[ 4533]='h00000000;
    rd_cycle[ 4534] = 1'b1;  wr_cycle[ 4534] = 1'b0;  addr_rom[ 4534]='h00002490;  wr_data_rom[ 4534]='h00000000;
    rd_cycle[ 4535] = 1'b1;  wr_cycle[ 4535] = 1'b0;  addr_rom[ 4535]='h000007e4;  wr_data_rom[ 4535]='h00000000;
    rd_cycle[ 4536] = 1'b1;  wr_cycle[ 4536] = 1'b0;  addr_rom[ 4536]='h00002514;  wr_data_rom[ 4536]='h00000000;
    rd_cycle[ 4537] = 1'b0;  wr_cycle[ 4537] = 1'b1;  addr_rom[ 4537]='h00003fdc;  wr_data_rom[ 4537]='h00003f01;
    rd_cycle[ 4538] = 1'b0;  wr_cycle[ 4538] = 1'b1;  addr_rom[ 4538]='h000019a8;  wr_data_rom[ 4538]='h00000579;
    rd_cycle[ 4539] = 1'b0;  wr_cycle[ 4539] = 1'b1;  addr_rom[ 4539]='h00001038;  wr_data_rom[ 4539]='h000036d1;
    rd_cycle[ 4540] = 1'b0;  wr_cycle[ 4540] = 1'b1;  addr_rom[ 4540]='h00003fbc;  wr_data_rom[ 4540]='h0000329d;
    rd_cycle[ 4541] = 1'b0;  wr_cycle[ 4541] = 1'b1;  addr_rom[ 4541]='h00003414;  wr_data_rom[ 4541]='h000017df;
    rd_cycle[ 4542] = 1'b1;  wr_cycle[ 4542] = 1'b0;  addr_rom[ 4542]='h00002028;  wr_data_rom[ 4542]='h00000000;
    rd_cycle[ 4543] = 1'b0;  wr_cycle[ 4543] = 1'b1;  addr_rom[ 4543]='h00002f0c;  wr_data_rom[ 4543]='h00002adb;
    rd_cycle[ 4544] = 1'b1;  wr_cycle[ 4544] = 1'b0;  addr_rom[ 4544]='h00003548;  wr_data_rom[ 4544]='h00000000;
    rd_cycle[ 4545] = 1'b1;  wr_cycle[ 4545] = 1'b0;  addr_rom[ 4545]='h00002f94;  wr_data_rom[ 4545]='h00000000;
    rd_cycle[ 4546] = 1'b0;  wr_cycle[ 4546] = 1'b1;  addr_rom[ 4546]='h00002918;  wr_data_rom[ 4546]='h000005ab;
    rd_cycle[ 4547] = 1'b1;  wr_cycle[ 4547] = 1'b0;  addr_rom[ 4547]='h0000397c;  wr_data_rom[ 4547]='h00000000;
    rd_cycle[ 4548] = 1'b1;  wr_cycle[ 4548] = 1'b0;  addr_rom[ 4548]='h000038f4;  wr_data_rom[ 4548]='h00000000;
    rd_cycle[ 4549] = 1'b1;  wr_cycle[ 4549] = 1'b0;  addr_rom[ 4549]='h000014f0;  wr_data_rom[ 4549]='h00000000;
    rd_cycle[ 4550] = 1'b0;  wr_cycle[ 4550] = 1'b1;  addr_rom[ 4550]='h00003f74;  wr_data_rom[ 4550]='h000027ec;
    rd_cycle[ 4551] = 1'b1;  wr_cycle[ 4551] = 1'b0;  addr_rom[ 4551]='h00002650;  wr_data_rom[ 4551]='h00000000;
    rd_cycle[ 4552] = 1'b1;  wr_cycle[ 4552] = 1'b0;  addr_rom[ 4552]='h0000343c;  wr_data_rom[ 4552]='h00000000;
    rd_cycle[ 4553] = 1'b1;  wr_cycle[ 4553] = 1'b0;  addr_rom[ 4553]='h00002fd0;  wr_data_rom[ 4553]='h00000000;
    rd_cycle[ 4554] = 1'b0;  wr_cycle[ 4554] = 1'b1;  addr_rom[ 4554]='h00000630;  wr_data_rom[ 4554]='h00000eda;
    rd_cycle[ 4555] = 1'b0;  wr_cycle[ 4555] = 1'b1;  addr_rom[ 4555]='h00001ce4;  wr_data_rom[ 4555]='h00001fce;
    rd_cycle[ 4556] = 1'b1;  wr_cycle[ 4556] = 1'b0;  addr_rom[ 4556]='h00002d30;  wr_data_rom[ 4556]='h00000000;
    rd_cycle[ 4557] = 1'b1;  wr_cycle[ 4557] = 1'b0;  addr_rom[ 4557]='h00003218;  wr_data_rom[ 4557]='h00000000;
    rd_cycle[ 4558] = 1'b0;  wr_cycle[ 4558] = 1'b1;  addr_rom[ 4558]='h000001b0;  wr_data_rom[ 4558]='h000009a6;
    rd_cycle[ 4559] = 1'b1;  wr_cycle[ 4559] = 1'b0;  addr_rom[ 4559]='h00001adc;  wr_data_rom[ 4559]='h00000000;
    rd_cycle[ 4560] = 1'b0;  wr_cycle[ 4560] = 1'b1;  addr_rom[ 4560]='h00002114;  wr_data_rom[ 4560]='h00002049;
    rd_cycle[ 4561] = 1'b0;  wr_cycle[ 4561] = 1'b1;  addr_rom[ 4561]='h00003430;  wr_data_rom[ 4561]='h000031e0;
    rd_cycle[ 4562] = 1'b1;  wr_cycle[ 4562] = 1'b0;  addr_rom[ 4562]='h00001970;  wr_data_rom[ 4562]='h00000000;
    rd_cycle[ 4563] = 1'b1;  wr_cycle[ 4563] = 1'b0;  addr_rom[ 4563]='h00002020;  wr_data_rom[ 4563]='h00000000;
    rd_cycle[ 4564] = 1'b0;  wr_cycle[ 4564] = 1'b1;  addr_rom[ 4564]='h000001ec;  wr_data_rom[ 4564]='h00002ae7;
    rd_cycle[ 4565] = 1'b0;  wr_cycle[ 4565] = 1'b1;  addr_rom[ 4565]='h00003c54;  wr_data_rom[ 4565]='h0000209e;
    rd_cycle[ 4566] = 1'b0;  wr_cycle[ 4566] = 1'b1;  addr_rom[ 4566]='h0000085c;  wr_data_rom[ 4566]='h00000f80;
    rd_cycle[ 4567] = 1'b1;  wr_cycle[ 4567] = 1'b0;  addr_rom[ 4567]='h00000924;  wr_data_rom[ 4567]='h00000000;
    rd_cycle[ 4568] = 1'b1;  wr_cycle[ 4568] = 1'b0;  addr_rom[ 4568]='h000013e4;  wr_data_rom[ 4568]='h00000000;
    rd_cycle[ 4569] = 1'b1;  wr_cycle[ 4569] = 1'b0;  addr_rom[ 4569]='h00000b7c;  wr_data_rom[ 4569]='h00000000;
    rd_cycle[ 4570] = 1'b1;  wr_cycle[ 4570] = 1'b0;  addr_rom[ 4570]='h00002ed8;  wr_data_rom[ 4570]='h00000000;
    rd_cycle[ 4571] = 1'b0;  wr_cycle[ 4571] = 1'b1;  addr_rom[ 4571]='h00003844;  wr_data_rom[ 4571]='h00000aa0;
    rd_cycle[ 4572] = 1'b1;  wr_cycle[ 4572] = 1'b0;  addr_rom[ 4572]='h00000804;  wr_data_rom[ 4572]='h00000000;
    rd_cycle[ 4573] = 1'b0;  wr_cycle[ 4573] = 1'b1;  addr_rom[ 4573]='h00001e14;  wr_data_rom[ 4573]='h000015da;
    rd_cycle[ 4574] = 1'b1;  wr_cycle[ 4574] = 1'b0;  addr_rom[ 4574]='h0000355c;  wr_data_rom[ 4574]='h00000000;
    rd_cycle[ 4575] = 1'b1;  wr_cycle[ 4575] = 1'b0;  addr_rom[ 4575]='h00002a98;  wr_data_rom[ 4575]='h00000000;
    rd_cycle[ 4576] = 1'b0;  wr_cycle[ 4576] = 1'b1;  addr_rom[ 4576]='h00000f18;  wr_data_rom[ 4576]='h00002a5c;
    rd_cycle[ 4577] = 1'b1;  wr_cycle[ 4577] = 1'b0;  addr_rom[ 4577]='h00002504;  wr_data_rom[ 4577]='h00000000;
    rd_cycle[ 4578] = 1'b0;  wr_cycle[ 4578] = 1'b1;  addr_rom[ 4578]='h00002318;  wr_data_rom[ 4578]='h00001582;
    rd_cycle[ 4579] = 1'b1;  wr_cycle[ 4579] = 1'b0;  addr_rom[ 4579]='h000039a4;  wr_data_rom[ 4579]='h00000000;
    rd_cycle[ 4580] = 1'b1;  wr_cycle[ 4580] = 1'b0;  addr_rom[ 4580]='h00000088;  wr_data_rom[ 4580]='h00000000;
    rd_cycle[ 4581] = 1'b1;  wr_cycle[ 4581] = 1'b0;  addr_rom[ 4581]='h000035d4;  wr_data_rom[ 4581]='h00000000;
    rd_cycle[ 4582] = 1'b1;  wr_cycle[ 4582] = 1'b0;  addr_rom[ 4582]='h00001880;  wr_data_rom[ 4582]='h00000000;
    rd_cycle[ 4583] = 1'b1;  wr_cycle[ 4583] = 1'b0;  addr_rom[ 4583]='h00003424;  wr_data_rom[ 4583]='h00000000;
    rd_cycle[ 4584] = 1'b0;  wr_cycle[ 4584] = 1'b1;  addr_rom[ 4584]='h00003764;  wr_data_rom[ 4584]='h00001509;
    rd_cycle[ 4585] = 1'b1;  wr_cycle[ 4585] = 1'b0;  addr_rom[ 4585]='h0000081c;  wr_data_rom[ 4585]='h00000000;
    rd_cycle[ 4586] = 1'b0;  wr_cycle[ 4586] = 1'b1;  addr_rom[ 4586]='h00003c44;  wr_data_rom[ 4586]='h00002e27;
    rd_cycle[ 4587] = 1'b0;  wr_cycle[ 4587] = 1'b1;  addr_rom[ 4587]='h00002e68;  wr_data_rom[ 4587]='h00001d0b;
    rd_cycle[ 4588] = 1'b0;  wr_cycle[ 4588] = 1'b1;  addr_rom[ 4588]='h00003000;  wr_data_rom[ 4588]='h00002d44;
    rd_cycle[ 4589] = 1'b0;  wr_cycle[ 4589] = 1'b1;  addr_rom[ 4589]='h00003d94;  wr_data_rom[ 4589]='h0000117d;
    rd_cycle[ 4590] = 1'b1;  wr_cycle[ 4590] = 1'b0;  addr_rom[ 4590]='h00003a8c;  wr_data_rom[ 4590]='h00000000;
    rd_cycle[ 4591] = 1'b1;  wr_cycle[ 4591] = 1'b0;  addr_rom[ 4591]='h00001c90;  wr_data_rom[ 4591]='h00000000;
    rd_cycle[ 4592] = 1'b1;  wr_cycle[ 4592] = 1'b0;  addr_rom[ 4592]='h00001e6c;  wr_data_rom[ 4592]='h00000000;
    rd_cycle[ 4593] = 1'b1;  wr_cycle[ 4593] = 1'b0;  addr_rom[ 4593]='h00000ebc;  wr_data_rom[ 4593]='h00000000;
    rd_cycle[ 4594] = 1'b0;  wr_cycle[ 4594] = 1'b1;  addr_rom[ 4594]='h0000149c;  wr_data_rom[ 4594]='h00003d9c;
    rd_cycle[ 4595] = 1'b0;  wr_cycle[ 4595] = 1'b1;  addr_rom[ 4595]='h00001b7c;  wr_data_rom[ 4595]='h00002bc5;
    rd_cycle[ 4596] = 1'b1;  wr_cycle[ 4596] = 1'b0;  addr_rom[ 4596]='h00002bac;  wr_data_rom[ 4596]='h00000000;
    rd_cycle[ 4597] = 1'b0;  wr_cycle[ 4597] = 1'b1;  addr_rom[ 4597]='h00000b04;  wr_data_rom[ 4597]='h0000297e;
    rd_cycle[ 4598] = 1'b1;  wr_cycle[ 4598] = 1'b0;  addr_rom[ 4598]='h000030b0;  wr_data_rom[ 4598]='h00000000;
    rd_cycle[ 4599] = 1'b0;  wr_cycle[ 4599] = 1'b1;  addr_rom[ 4599]='h000009ac;  wr_data_rom[ 4599]='h000027a1;
    rd_cycle[ 4600] = 1'b1;  wr_cycle[ 4600] = 1'b0;  addr_rom[ 4600]='h00003c08;  wr_data_rom[ 4600]='h00000000;
    rd_cycle[ 4601] = 1'b1;  wr_cycle[ 4601] = 1'b0;  addr_rom[ 4601]='h00002f20;  wr_data_rom[ 4601]='h00000000;
    rd_cycle[ 4602] = 1'b0;  wr_cycle[ 4602] = 1'b1;  addr_rom[ 4602]='h0000373c;  wr_data_rom[ 4602]='h0000165c;
    rd_cycle[ 4603] = 1'b0;  wr_cycle[ 4603] = 1'b1;  addr_rom[ 4603]='h000036b4;  wr_data_rom[ 4603]='h000010de;
    rd_cycle[ 4604] = 1'b0;  wr_cycle[ 4604] = 1'b1;  addr_rom[ 4604]='h000014e4;  wr_data_rom[ 4604]='h0000047e;
    rd_cycle[ 4605] = 1'b0;  wr_cycle[ 4605] = 1'b1;  addr_rom[ 4605]='h00003fa4;  wr_data_rom[ 4605]='h00000933;
    rd_cycle[ 4606] = 1'b1;  wr_cycle[ 4606] = 1'b0;  addr_rom[ 4606]='h00003118;  wr_data_rom[ 4606]='h00000000;
    rd_cycle[ 4607] = 1'b0;  wr_cycle[ 4607] = 1'b1;  addr_rom[ 4607]='h00000674;  wr_data_rom[ 4607]='h00002409;
    rd_cycle[ 4608] = 1'b1;  wr_cycle[ 4608] = 1'b0;  addr_rom[ 4608]='h00003d58;  wr_data_rom[ 4608]='h00000000;
    rd_cycle[ 4609] = 1'b0;  wr_cycle[ 4609] = 1'b1;  addr_rom[ 4609]='h00002bd8;  wr_data_rom[ 4609]='h00000704;
    rd_cycle[ 4610] = 1'b0;  wr_cycle[ 4610] = 1'b1;  addr_rom[ 4610]='h00002e10;  wr_data_rom[ 4610]='h00003ad8;
    rd_cycle[ 4611] = 1'b1;  wr_cycle[ 4611] = 1'b0;  addr_rom[ 4611]='h00002338;  wr_data_rom[ 4611]='h00000000;
    rd_cycle[ 4612] = 1'b1;  wr_cycle[ 4612] = 1'b0;  addr_rom[ 4612]='h00000eb0;  wr_data_rom[ 4612]='h00000000;
    rd_cycle[ 4613] = 1'b0;  wr_cycle[ 4613] = 1'b1;  addr_rom[ 4613]='h0000324c;  wr_data_rom[ 4613]='h00002a1d;
    rd_cycle[ 4614] = 1'b1;  wr_cycle[ 4614] = 1'b0;  addr_rom[ 4614]='h00001bb4;  wr_data_rom[ 4614]='h00000000;
    rd_cycle[ 4615] = 1'b1;  wr_cycle[ 4615] = 1'b0;  addr_rom[ 4615]='h000008c0;  wr_data_rom[ 4615]='h00000000;
    rd_cycle[ 4616] = 1'b1;  wr_cycle[ 4616] = 1'b0;  addr_rom[ 4616]='h00003028;  wr_data_rom[ 4616]='h00000000;
    rd_cycle[ 4617] = 1'b1;  wr_cycle[ 4617] = 1'b0;  addr_rom[ 4617]='h00003588;  wr_data_rom[ 4617]='h00000000;
    rd_cycle[ 4618] = 1'b1;  wr_cycle[ 4618] = 1'b0;  addr_rom[ 4618]='h000011ac;  wr_data_rom[ 4618]='h00000000;
    rd_cycle[ 4619] = 1'b1;  wr_cycle[ 4619] = 1'b0;  addr_rom[ 4619]='h00001b00;  wr_data_rom[ 4619]='h00000000;
    rd_cycle[ 4620] = 1'b1;  wr_cycle[ 4620] = 1'b0;  addr_rom[ 4620]='h00001c70;  wr_data_rom[ 4620]='h00000000;
    rd_cycle[ 4621] = 1'b1;  wr_cycle[ 4621] = 1'b0;  addr_rom[ 4621]='h00003904;  wr_data_rom[ 4621]='h00000000;
    rd_cycle[ 4622] = 1'b0;  wr_cycle[ 4622] = 1'b1;  addr_rom[ 4622]='h00001ce8;  wr_data_rom[ 4622]='h00001217;
    rd_cycle[ 4623] = 1'b0;  wr_cycle[ 4623] = 1'b1;  addr_rom[ 4623]='h00003ec0;  wr_data_rom[ 4623]='h000022c5;
    rd_cycle[ 4624] = 1'b1;  wr_cycle[ 4624] = 1'b0;  addr_rom[ 4624]='h00001fd4;  wr_data_rom[ 4624]='h00000000;
    rd_cycle[ 4625] = 1'b0;  wr_cycle[ 4625] = 1'b1;  addr_rom[ 4625]='h0000046c;  wr_data_rom[ 4625]='h00002ad2;
    rd_cycle[ 4626] = 1'b0;  wr_cycle[ 4626] = 1'b1;  addr_rom[ 4626]='h00002088;  wr_data_rom[ 4626]='h00000ec1;
    rd_cycle[ 4627] = 1'b0;  wr_cycle[ 4627] = 1'b1;  addr_rom[ 4627]='h000025e8;  wr_data_rom[ 4627]='h00002121;
    rd_cycle[ 4628] = 1'b0;  wr_cycle[ 4628] = 1'b1;  addr_rom[ 4628]='h00000f70;  wr_data_rom[ 4628]='h00002f0a;
    rd_cycle[ 4629] = 1'b0;  wr_cycle[ 4629] = 1'b1;  addr_rom[ 4629]='h000028ac;  wr_data_rom[ 4629]='h00000a0e;
    rd_cycle[ 4630] = 1'b0;  wr_cycle[ 4630] = 1'b1;  addr_rom[ 4630]='h000015e0;  wr_data_rom[ 4630]='h00002708;
    rd_cycle[ 4631] = 1'b1;  wr_cycle[ 4631] = 1'b0;  addr_rom[ 4631]='h00000e84;  wr_data_rom[ 4631]='h00000000;
    rd_cycle[ 4632] = 1'b0;  wr_cycle[ 4632] = 1'b1;  addr_rom[ 4632]='h00000ed4;  wr_data_rom[ 4632]='h00001468;
    rd_cycle[ 4633] = 1'b0;  wr_cycle[ 4633] = 1'b1;  addr_rom[ 4633]='h000013a0;  wr_data_rom[ 4633]='h00003148;
    rd_cycle[ 4634] = 1'b1;  wr_cycle[ 4634] = 1'b0;  addr_rom[ 4634]='h00002294;  wr_data_rom[ 4634]='h00000000;
    rd_cycle[ 4635] = 1'b0;  wr_cycle[ 4635] = 1'b1;  addr_rom[ 4635]='h00001d6c;  wr_data_rom[ 4635]='h00002251;
    rd_cycle[ 4636] = 1'b1;  wr_cycle[ 4636] = 1'b0;  addr_rom[ 4636]='h000028e8;  wr_data_rom[ 4636]='h00000000;
    rd_cycle[ 4637] = 1'b0;  wr_cycle[ 4637] = 1'b1;  addr_rom[ 4637]='h00001874;  wr_data_rom[ 4637]='h00001d8e;
    rd_cycle[ 4638] = 1'b1;  wr_cycle[ 4638] = 1'b0;  addr_rom[ 4638]='h0000133c;  wr_data_rom[ 4638]='h00000000;
    rd_cycle[ 4639] = 1'b0;  wr_cycle[ 4639] = 1'b1;  addr_rom[ 4639]='h00003078;  wr_data_rom[ 4639]='h00003ea0;
    rd_cycle[ 4640] = 1'b1;  wr_cycle[ 4640] = 1'b0;  addr_rom[ 4640]='h000039a0;  wr_data_rom[ 4640]='h00000000;
    rd_cycle[ 4641] = 1'b0;  wr_cycle[ 4641] = 1'b1;  addr_rom[ 4641]='h000019e8;  wr_data_rom[ 4641]='h00001fca;
    rd_cycle[ 4642] = 1'b1;  wr_cycle[ 4642] = 1'b0;  addr_rom[ 4642]='h00003c50;  wr_data_rom[ 4642]='h00000000;
    rd_cycle[ 4643] = 1'b1;  wr_cycle[ 4643] = 1'b0;  addr_rom[ 4643]='h000001e4;  wr_data_rom[ 4643]='h00000000;
    rd_cycle[ 4644] = 1'b1;  wr_cycle[ 4644] = 1'b0;  addr_rom[ 4644]='h00001740;  wr_data_rom[ 4644]='h00000000;
    rd_cycle[ 4645] = 1'b1;  wr_cycle[ 4645] = 1'b0;  addr_rom[ 4645]='h00001d00;  wr_data_rom[ 4645]='h00000000;
    rd_cycle[ 4646] = 1'b1;  wr_cycle[ 4646] = 1'b0;  addr_rom[ 4646]='h00003e74;  wr_data_rom[ 4646]='h00000000;
    rd_cycle[ 4647] = 1'b0;  wr_cycle[ 4647] = 1'b1;  addr_rom[ 4647]='h00000c58;  wr_data_rom[ 4647]='h00001e7b;
    rd_cycle[ 4648] = 1'b0;  wr_cycle[ 4648] = 1'b1;  addr_rom[ 4648]='h000038cc;  wr_data_rom[ 4648]='h00003518;
    rd_cycle[ 4649] = 1'b1;  wr_cycle[ 4649] = 1'b0;  addr_rom[ 4649]='h00002000;  wr_data_rom[ 4649]='h00000000;
    rd_cycle[ 4650] = 1'b1;  wr_cycle[ 4650] = 1'b0;  addr_rom[ 4650]='h000034b8;  wr_data_rom[ 4650]='h00000000;
    rd_cycle[ 4651] = 1'b1;  wr_cycle[ 4651] = 1'b0;  addr_rom[ 4651]='h00003f68;  wr_data_rom[ 4651]='h00000000;
    rd_cycle[ 4652] = 1'b1;  wr_cycle[ 4652] = 1'b0;  addr_rom[ 4652]='h00000c44;  wr_data_rom[ 4652]='h00000000;
    rd_cycle[ 4653] = 1'b1;  wr_cycle[ 4653] = 1'b0;  addr_rom[ 4653]='h00001638;  wr_data_rom[ 4653]='h00000000;
    rd_cycle[ 4654] = 1'b1;  wr_cycle[ 4654] = 1'b0;  addr_rom[ 4654]='h00000478;  wr_data_rom[ 4654]='h00000000;
    rd_cycle[ 4655] = 1'b1;  wr_cycle[ 4655] = 1'b0;  addr_rom[ 4655]='h00002058;  wr_data_rom[ 4655]='h00000000;
    rd_cycle[ 4656] = 1'b0;  wr_cycle[ 4656] = 1'b1;  addr_rom[ 4656]='h00003e1c;  wr_data_rom[ 4656]='h00000007;
    rd_cycle[ 4657] = 1'b0;  wr_cycle[ 4657] = 1'b1;  addr_rom[ 4657]='h00001f98;  wr_data_rom[ 4657]='h000023e1;
    rd_cycle[ 4658] = 1'b1;  wr_cycle[ 4658] = 1'b0;  addr_rom[ 4658]='h00000f04;  wr_data_rom[ 4658]='h00000000;
    rd_cycle[ 4659] = 1'b1;  wr_cycle[ 4659] = 1'b0;  addr_rom[ 4659]='h00001510;  wr_data_rom[ 4659]='h00000000;
    rd_cycle[ 4660] = 1'b0;  wr_cycle[ 4660] = 1'b1;  addr_rom[ 4660]='h0000284c;  wr_data_rom[ 4660]='h000028cb;
    rd_cycle[ 4661] = 1'b0;  wr_cycle[ 4661] = 1'b1;  addr_rom[ 4661]='h00002670;  wr_data_rom[ 4661]='h000015f3;
    rd_cycle[ 4662] = 1'b0;  wr_cycle[ 4662] = 1'b1;  addr_rom[ 4662]='h00003e00;  wr_data_rom[ 4662]='h00000226;
    rd_cycle[ 4663] = 1'b0;  wr_cycle[ 4663] = 1'b1;  addr_rom[ 4663]='h00003460;  wr_data_rom[ 4663]='h00000169;
    rd_cycle[ 4664] = 1'b1;  wr_cycle[ 4664] = 1'b0;  addr_rom[ 4664]='h0000380c;  wr_data_rom[ 4664]='h00000000;
    rd_cycle[ 4665] = 1'b0;  wr_cycle[ 4665] = 1'b1;  addr_rom[ 4665]='h00003fa4;  wr_data_rom[ 4665]='h0000042b;
    rd_cycle[ 4666] = 1'b1;  wr_cycle[ 4666] = 1'b0;  addr_rom[ 4666]='h00003520;  wr_data_rom[ 4666]='h00000000;
    rd_cycle[ 4667] = 1'b1;  wr_cycle[ 4667] = 1'b0;  addr_rom[ 4667]='h00000bfc;  wr_data_rom[ 4667]='h00000000;
    rd_cycle[ 4668] = 1'b0;  wr_cycle[ 4668] = 1'b1;  addr_rom[ 4668]='h00001b14;  wr_data_rom[ 4668]='h00001f22;
    rd_cycle[ 4669] = 1'b0;  wr_cycle[ 4669] = 1'b1;  addr_rom[ 4669]='h00003130;  wr_data_rom[ 4669]='h000027d4;
    rd_cycle[ 4670] = 1'b0;  wr_cycle[ 4670] = 1'b1;  addr_rom[ 4670]='h00001760;  wr_data_rom[ 4670]='h0000376e;
    rd_cycle[ 4671] = 1'b1;  wr_cycle[ 4671] = 1'b0;  addr_rom[ 4671]='h00000ef8;  wr_data_rom[ 4671]='h00000000;
    rd_cycle[ 4672] = 1'b0;  wr_cycle[ 4672] = 1'b1;  addr_rom[ 4672]='h00002adc;  wr_data_rom[ 4672]='h00002d76;
    rd_cycle[ 4673] = 1'b0;  wr_cycle[ 4673] = 1'b1;  addr_rom[ 4673]='h00003aac;  wr_data_rom[ 4673]='h000007c3;
    rd_cycle[ 4674] = 1'b0;  wr_cycle[ 4674] = 1'b1;  addr_rom[ 4674]='h00001aa8;  wr_data_rom[ 4674]='h00000bd0;
    rd_cycle[ 4675] = 1'b1;  wr_cycle[ 4675] = 1'b0;  addr_rom[ 4675]='h000026d0;  wr_data_rom[ 4675]='h00000000;
    rd_cycle[ 4676] = 1'b0;  wr_cycle[ 4676] = 1'b1;  addr_rom[ 4676]='h00002364;  wr_data_rom[ 4676]='h00000825;
    rd_cycle[ 4677] = 1'b1;  wr_cycle[ 4677] = 1'b0;  addr_rom[ 4677]='h00001518;  wr_data_rom[ 4677]='h00000000;
    rd_cycle[ 4678] = 1'b0;  wr_cycle[ 4678] = 1'b1;  addr_rom[ 4678]='h00003d24;  wr_data_rom[ 4678]='h000007d1;
    rd_cycle[ 4679] = 1'b0;  wr_cycle[ 4679] = 1'b1;  addr_rom[ 4679]='h00000084;  wr_data_rom[ 4679]='h0000288b;
    rd_cycle[ 4680] = 1'b0;  wr_cycle[ 4680] = 1'b1;  addr_rom[ 4680]='h00002de4;  wr_data_rom[ 4680]='h00000b78;
    rd_cycle[ 4681] = 1'b0;  wr_cycle[ 4681] = 1'b1;  addr_rom[ 4681]='h000035c0;  wr_data_rom[ 4681]='h000019c4;
    rd_cycle[ 4682] = 1'b0;  wr_cycle[ 4682] = 1'b1;  addr_rom[ 4682]='h00001128;  wr_data_rom[ 4682]='h0000337e;
    rd_cycle[ 4683] = 1'b1;  wr_cycle[ 4683] = 1'b0;  addr_rom[ 4683]='h00000060;  wr_data_rom[ 4683]='h00000000;
    rd_cycle[ 4684] = 1'b1;  wr_cycle[ 4684] = 1'b0;  addr_rom[ 4684]='h00002454;  wr_data_rom[ 4684]='h00000000;
    rd_cycle[ 4685] = 1'b1;  wr_cycle[ 4685] = 1'b0;  addr_rom[ 4685]='h00003f28;  wr_data_rom[ 4685]='h00000000;
    rd_cycle[ 4686] = 1'b1;  wr_cycle[ 4686] = 1'b0;  addr_rom[ 4686]='h00000ca8;  wr_data_rom[ 4686]='h00000000;
    rd_cycle[ 4687] = 1'b1;  wr_cycle[ 4687] = 1'b0;  addr_rom[ 4687]='h00001e0c;  wr_data_rom[ 4687]='h00000000;
    rd_cycle[ 4688] = 1'b0;  wr_cycle[ 4688] = 1'b1;  addr_rom[ 4688]='h0000017c;  wr_data_rom[ 4688]='h000016ec;
    rd_cycle[ 4689] = 1'b0;  wr_cycle[ 4689] = 1'b1;  addr_rom[ 4689]='h00002f4c;  wr_data_rom[ 4689]='h00002eb4;
    rd_cycle[ 4690] = 1'b0;  wr_cycle[ 4690] = 1'b1;  addr_rom[ 4690]='h00003a8c;  wr_data_rom[ 4690]='h000022bb;
    rd_cycle[ 4691] = 1'b1;  wr_cycle[ 4691] = 1'b0;  addr_rom[ 4691]='h00003fec;  wr_data_rom[ 4691]='h00000000;
    rd_cycle[ 4692] = 1'b1;  wr_cycle[ 4692] = 1'b0;  addr_rom[ 4692]='h000011a0;  wr_data_rom[ 4692]='h00000000;
    rd_cycle[ 4693] = 1'b1;  wr_cycle[ 4693] = 1'b0;  addr_rom[ 4693]='h00001e5c;  wr_data_rom[ 4693]='h00000000;
    rd_cycle[ 4694] = 1'b0;  wr_cycle[ 4694] = 1'b1;  addr_rom[ 4694]='h00001e6c;  wr_data_rom[ 4694]='h00002fa8;
    rd_cycle[ 4695] = 1'b1;  wr_cycle[ 4695] = 1'b0;  addr_rom[ 4695]='h00002d10;  wr_data_rom[ 4695]='h00000000;
    rd_cycle[ 4696] = 1'b1;  wr_cycle[ 4696] = 1'b0;  addr_rom[ 4696]='h00002314;  wr_data_rom[ 4696]='h00000000;
    rd_cycle[ 4697] = 1'b1;  wr_cycle[ 4697] = 1'b0;  addr_rom[ 4697]='h00000228;  wr_data_rom[ 4697]='h00000000;
    rd_cycle[ 4698] = 1'b0;  wr_cycle[ 4698] = 1'b1;  addr_rom[ 4698]='h000027b8;  wr_data_rom[ 4698]='h00001e35;
    rd_cycle[ 4699] = 1'b1;  wr_cycle[ 4699] = 1'b0;  addr_rom[ 4699]='h00003e9c;  wr_data_rom[ 4699]='h00000000;
    rd_cycle[ 4700] = 1'b0;  wr_cycle[ 4700] = 1'b1;  addr_rom[ 4700]='h00003018;  wr_data_rom[ 4700]='h00001656;
    rd_cycle[ 4701] = 1'b1;  wr_cycle[ 4701] = 1'b0;  addr_rom[ 4701]='h00000c00;  wr_data_rom[ 4701]='h00000000;
    rd_cycle[ 4702] = 1'b0;  wr_cycle[ 4702] = 1'b1;  addr_rom[ 4702]='h00000a10;  wr_data_rom[ 4702]='h000018be;
    rd_cycle[ 4703] = 1'b0;  wr_cycle[ 4703] = 1'b1;  addr_rom[ 4703]='h000031d4;  wr_data_rom[ 4703]='h00003e9c;
    rd_cycle[ 4704] = 1'b0;  wr_cycle[ 4704] = 1'b1;  addr_rom[ 4704]='h000039d0;  wr_data_rom[ 4704]='h000029b6;
    rd_cycle[ 4705] = 1'b0;  wr_cycle[ 4705] = 1'b1;  addr_rom[ 4705]='h00000b7c;  wr_data_rom[ 4705]='h00003aa2;
    rd_cycle[ 4706] = 1'b1;  wr_cycle[ 4706] = 1'b0;  addr_rom[ 4706]='h00001ef4;  wr_data_rom[ 4706]='h00000000;
    rd_cycle[ 4707] = 1'b0;  wr_cycle[ 4707] = 1'b1;  addr_rom[ 4707]='h00000110;  wr_data_rom[ 4707]='h00001b85;
    rd_cycle[ 4708] = 1'b1;  wr_cycle[ 4708] = 1'b0;  addr_rom[ 4708]='h00002840;  wr_data_rom[ 4708]='h00000000;
    rd_cycle[ 4709] = 1'b1;  wr_cycle[ 4709] = 1'b0;  addr_rom[ 4709]='h00000e4c;  wr_data_rom[ 4709]='h00000000;
    rd_cycle[ 4710] = 1'b0;  wr_cycle[ 4710] = 1'b1;  addr_rom[ 4710]='h00000ba0;  wr_data_rom[ 4710]='h000032fc;
    rd_cycle[ 4711] = 1'b0;  wr_cycle[ 4711] = 1'b1;  addr_rom[ 4711]='h00000598;  wr_data_rom[ 4711]='h00003886;
    rd_cycle[ 4712] = 1'b0;  wr_cycle[ 4712] = 1'b1;  addr_rom[ 4712]='h00003524;  wr_data_rom[ 4712]='h000001f9;
    rd_cycle[ 4713] = 1'b0;  wr_cycle[ 4713] = 1'b1;  addr_rom[ 4713]='h000005d0;  wr_data_rom[ 4713]='h000013ca;
    rd_cycle[ 4714] = 1'b0;  wr_cycle[ 4714] = 1'b1;  addr_rom[ 4714]='h00003460;  wr_data_rom[ 4714]='h000024fe;
    rd_cycle[ 4715] = 1'b0;  wr_cycle[ 4715] = 1'b1;  addr_rom[ 4715]='h000033ec;  wr_data_rom[ 4715]='h000020bd;
    rd_cycle[ 4716] = 1'b0;  wr_cycle[ 4716] = 1'b1;  addr_rom[ 4716]='h000008f8;  wr_data_rom[ 4716]='h00001f5c;
    rd_cycle[ 4717] = 1'b0;  wr_cycle[ 4717] = 1'b1;  addr_rom[ 4717]='h00002754;  wr_data_rom[ 4717]='h00000b0a;
    rd_cycle[ 4718] = 1'b1;  wr_cycle[ 4718] = 1'b0;  addr_rom[ 4718]='h000024ac;  wr_data_rom[ 4718]='h00000000;
    rd_cycle[ 4719] = 1'b0;  wr_cycle[ 4719] = 1'b1;  addr_rom[ 4719]='h00000e08;  wr_data_rom[ 4719]='h00001fea;
    rd_cycle[ 4720] = 1'b0;  wr_cycle[ 4720] = 1'b1;  addr_rom[ 4720]='h00002474;  wr_data_rom[ 4720]='h00002a65;
    rd_cycle[ 4721] = 1'b1;  wr_cycle[ 4721] = 1'b0;  addr_rom[ 4721]='h000039c4;  wr_data_rom[ 4721]='h00000000;
    rd_cycle[ 4722] = 1'b0;  wr_cycle[ 4722] = 1'b1;  addr_rom[ 4722]='h00001e64;  wr_data_rom[ 4722]='h00000823;
    rd_cycle[ 4723] = 1'b1;  wr_cycle[ 4723] = 1'b0;  addr_rom[ 4723]='h000018e0;  wr_data_rom[ 4723]='h00000000;
    rd_cycle[ 4724] = 1'b0;  wr_cycle[ 4724] = 1'b1;  addr_rom[ 4724]='h00003d8c;  wr_data_rom[ 4724]='h000004cb;
    rd_cycle[ 4725] = 1'b0;  wr_cycle[ 4725] = 1'b1;  addr_rom[ 4725]='h00000580;  wr_data_rom[ 4725]='h00003e31;
    rd_cycle[ 4726] = 1'b0;  wr_cycle[ 4726] = 1'b1;  addr_rom[ 4726]='h000016f0;  wr_data_rom[ 4726]='h0000013d;
    rd_cycle[ 4727] = 1'b0;  wr_cycle[ 4727] = 1'b1;  addr_rom[ 4727]='h000034bc;  wr_data_rom[ 4727]='h00003d85;
    rd_cycle[ 4728] = 1'b1;  wr_cycle[ 4728] = 1'b0;  addr_rom[ 4728]='h0000122c;  wr_data_rom[ 4728]='h00000000;
    rd_cycle[ 4729] = 1'b1;  wr_cycle[ 4729] = 1'b0;  addr_rom[ 4729]='h00002f58;  wr_data_rom[ 4729]='h00000000;
    rd_cycle[ 4730] = 1'b0;  wr_cycle[ 4730] = 1'b1;  addr_rom[ 4730]='h00001df8;  wr_data_rom[ 4730]='h0000385f;
    rd_cycle[ 4731] = 1'b0;  wr_cycle[ 4731] = 1'b1;  addr_rom[ 4731]='h00002e04;  wr_data_rom[ 4731]='h00002fe3;
    rd_cycle[ 4732] = 1'b0;  wr_cycle[ 4732] = 1'b1;  addr_rom[ 4732]='h00001abc;  wr_data_rom[ 4732]='h000005ff;
    rd_cycle[ 4733] = 1'b0;  wr_cycle[ 4733] = 1'b1;  addr_rom[ 4733]='h00001520;  wr_data_rom[ 4733]='h0000242b;
    rd_cycle[ 4734] = 1'b0;  wr_cycle[ 4734] = 1'b1;  addr_rom[ 4734]='h000008bc;  wr_data_rom[ 4734]='h0000143d;
    rd_cycle[ 4735] = 1'b0;  wr_cycle[ 4735] = 1'b1;  addr_rom[ 4735]='h00000870;  wr_data_rom[ 4735]='h000009e6;
    rd_cycle[ 4736] = 1'b1;  wr_cycle[ 4736] = 1'b0;  addr_rom[ 4736]='h000032a4;  wr_data_rom[ 4736]='h00000000;
    rd_cycle[ 4737] = 1'b0;  wr_cycle[ 4737] = 1'b1;  addr_rom[ 4737]='h00003194;  wr_data_rom[ 4737]='h000030a5;
    rd_cycle[ 4738] = 1'b1;  wr_cycle[ 4738] = 1'b0;  addr_rom[ 4738]='h00002f1c;  wr_data_rom[ 4738]='h00000000;
    rd_cycle[ 4739] = 1'b1;  wr_cycle[ 4739] = 1'b0;  addr_rom[ 4739]='h00000268;  wr_data_rom[ 4739]='h00000000;
    rd_cycle[ 4740] = 1'b1;  wr_cycle[ 4740] = 1'b0;  addr_rom[ 4740]='h00001218;  wr_data_rom[ 4740]='h00000000;
    rd_cycle[ 4741] = 1'b0;  wr_cycle[ 4741] = 1'b1;  addr_rom[ 4741]='h00000b00;  wr_data_rom[ 4741]='h000033c4;
    rd_cycle[ 4742] = 1'b0;  wr_cycle[ 4742] = 1'b1;  addr_rom[ 4742]='h000017b8;  wr_data_rom[ 4742]='h000038ae;
    rd_cycle[ 4743] = 1'b1;  wr_cycle[ 4743] = 1'b0;  addr_rom[ 4743]='h000027e8;  wr_data_rom[ 4743]='h00000000;
    rd_cycle[ 4744] = 1'b1;  wr_cycle[ 4744] = 1'b0;  addr_rom[ 4744]='h000039f4;  wr_data_rom[ 4744]='h00000000;
    rd_cycle[ 4745] = 1'b1;  wr_cycle[ 4745] = 1'b0;  addr_rom[ 4745]='h000028bc;  wr_data_rom[ 4745]='h00000000;
    rd_cycle[ 4746] = 1'b0;  wr_cycle[ 4746] = 1'b1;  addr_rom[ 4746]='h00002f88;  wr_data_rom[ 4746]='h00000a22;
    rd_cycle[ 4747] = 1'b0;  wr_cycle[ 4747] = 1'b1;  addr_rom[ 4747]='h00003fc8;  wr_data_rom[ 4747]='h000034d3;
    rd_cycle[ 4748] = 1'b1;  wr_cycle[ 4748] = 1'b0;  addr_rom[ 4748]='h0000290c;  wr_data_rom[ 4748]='h00000000;
    rd_cycle[ 4749] = 1'b0;  wr_cycle[ 4749] = 1'b1;  addr_rom[ 4749]='h00002cc8;  wr_data_rom[ 4749]='h00003ecc;
    rd_cycle[ 4750] = 1'b0;  wr_cycle[ 4750] = 1'b1;  addr_rom[ 4750]='h00000fc0;  wr_data_rom[ 4750]='h0000385c;
    rd_cycle[ 4751] = 1'b0;  wr_cycle[ 4751] = 1'b1;  addr_rom[ 4751]='h000023b4;  wr_data_rom[ 4751]='h00002cda;
    rd_cycle[ 4752] = 1'b1;  wr_cycle[ 4752] = 1'b0;  addr_rom[ 4752]='h00003e4c;  wr_data_rom[ 4752]='h00000000;
    rd_cycle[ 4753] = 1'b0;  wr_cycle[ 4753] = 1'b1;  addr_rom[ 4753]='h00001554;  wr_data_rom[ 4753]='h00002296;
    rd_cycle[ 4754] = 1'b1;  wr_cycle[ 4754] = 1'b0;  addr_rom[ 4754]='h00000cd0;  wr_data_rom[ 4754]='h00000000;
    rd_cycle[ 4755] = 1'b1;  wr_cycle[ 4755] = 1'b0;  addr_rom[ 4755]='h00000304;  wr_data_rom[ 4755]='h00000000;
    rd_cycle[ 4756] = 1'b1;  wr_cycle[ 4756] = 1'b0;  addr_rom[ 4756]='h00001108;  wr_data_rom[ 4756]='h00000000;
    rd_cycle[ 4757] = 1'b1;  wr_cycle[ 4757] = 1'b0;  addr_rom[ 4757]='h0000214c;  wr_data_rom[ 4757]='h00000000;
    rd_cycle[ 4758] = 1'b0;  wr_cycle[ 4758] = 1'b1;  addr_rom[ 4758]='h00000c9c;  wr_data_rom[ 4758]='h0000149e;
    rd_cycle[ 4759] = 1'b0;  wr_cycle[ 4759] = 1'b1;  addr_rom[ 4759]='h00002290;  wr_data_rom[ 4759]='h000001c2;
    rd_cycle[ 4760] = 1'b0;  wr_cycle[ 4760] = 1'b1;  addr_rom[ 4760]='h00000e54;  wr_data_rom[ 4760]='h00003267;
    rd_cycle[ 4761] = 1'b1;  wr_cycle[ 4761] = 1'b0;  addr_rom[ 4761]='h00000724;  wr_data_rom[ 4761]='h00000000;
    rd_cycle[ 4762] = 1'b0;  wr_cycle[ 4762] = 1'b1;  addr_rom[ 4762]='h00001944;  wr_data_rom[ 4762]='h00003c5c;
    rd_cycle[ 4763] = 1'b1;  wr_cycle[ 4763] = 1'b0;  addr_rom[ 4763]='h000011b0;  wr_data_rom[ 4763]='h00000000;
    rd_cycle[ 4764] = 1'b1;  wr_cycle[ 4764] = 1'b0;  addr_rom[ 4764]='h00000354;  wr_data_rom[ 4764]='h00000000;
    rd_cycle[ 4765] = 1'b1;  wr_cycle[ 4765] = 1'b0;  addr_rom[ 4765]='h000024b8;  wr_data_rom[ 4765]='h00000000;
    rd_cycle[ 4766] = 1'b1;  wr_cycle[ 4766] = 1'b0;  addr_rom[ 4766]='h000037d8;  wr_data_rom[ 4766]='h00000000;
    rd_cycle[ 4767] = 1'b1;  wr_cycle[ 4767] = 1'b0;  addr_rom[ 4767]='h00002f4c;  wr_data_rom[ 4767]='h00000000;
    rd_cycle[ 4768] = 1'b0;  wr_cycle[ 4768] = 1'b1;  addr_rom[ 4768]='h00003c10;  wr_data_rom[ 4768]='h000014cd;
    rd_cycle[ 4769] = 1'b1;  wr_cycle[ 4769] = 1'b0;  addr_rom[ 4769]='h00003ebc;  wr_data_rom[ 4769]='h00000000;
    rd_cycle[ 4770] = 1'b0;  wr_cycle[ 4770] = 1'b1;  addr_rom[ 4770]='h00003a5c;  wr_data_rom[ 4770]='h00001a96;
    rd_cycle[ 4771] = 1'b0;  wr_cycle[ 4771] = 1'b1;  addr_rom[ 4771]='h000034dc;  wr_data_rom[ 4771]='h00002f5a;
    rd_cycle[ 4772] = 1'b1;  wr_cycle[ 4772] = 1'b0;  addr_rom[ 4772]='h00003970;  wr_data_rom[ 4772]='h00000000;
    rd_cycle[ 4773] = 1'b0;  wr_cycle[ 4773] = 1'b1;  addr_rom[ 4773]='h00003a60;  wr_data_rom[ 4773]='h000039ae;
    rd_cycle[ 4774] = 1'b1;  wr_cycle[ 4774] = 1'b0;  addr_rom[ 4774]='h00003004;  wr_data_rom[ 4774]='h00000000;
    rd_cycle[ 4775] = 1'b0;  wr_cycle[ 4775] = 1'b1;  addr_rom[ 4775]='h00002b20;  wr_data_rom[ 4775]='h000012dd;
    rd_cycle[ 4776] = 1'b0;  wr_cycle[ 4776] = 1'b1;  addr_rom[ 4776]='h00000e0c;  wr_data_rom[ 4776]='h00000eca;
    rd_cycle[ 4777] = 1'b0;  wr_cycle[ 4777] = 1'b1;  addr_rom[ 4777]='h00003bac;  wr_data_rom[ 4777]='h0000181a;
    rd_cycle[ 4778] = 1'b1;  wr_cycle[ 4778] = 1'b0;  addr_rom[ 4778]='h0000168c;  wr_data_rom[ 4778]='h00000000;
    rd_cycle[ 4779] = 1'b1;  wr_cycle[ 4779] = 1'b0;  addr_rom[ 4779]='h00002c74;  wr_data_rom[ 4779]='h00000000;
    rd_cycle[ 4780] = 1'b0;  wr_cycle[ 4780] = 1'b1;  addr_rom[ 4780]='h000011e8;  wr_data_rom[ 4780]='h00000b26;
    rd_cycle[ 4781] = 1'b0;  wr_cycle[ 4781] = 1'b1;  addr_rom[ 4781]='h00000ef0;  wr_data_rom[ 4781]='h000039de;
    rd_cycle[ 4782] = 1'b1;  wr_cycle[ 4782] = 1'b0;  addr_rom[ 4782]='h00000358;  wr_data_rom[ 4782]='h00000000;
    rd_cycle[ 4783] = 1'b0;  wr_cycle[ 4783] = 1'b1;  addr_rom[ 4783]='h0000257c;  wr_data_rom[ 4783]='h00001e56;
    rd_cycle[ 4784] = 1'b1;  wr_cycle[ 4784] = 1'b0;  addr_rom[ 4784]='h00000400;  wr_data_rom[ 4784]='h00000000;
    rd_cycle[ 4785] = 1'b1;  wr_cycle[ 4785] = 1'b0;  addr_rom[ 4785]='h00002d30;  wr_data_rom[ 4785]='h00000000;
    rd_cycle[ 4786] = 1'b0;  wr_cycle[ 4786] = 1'b1;  addr_rom[ 4786]='h00003ff0;  wr_data_rom[ 4786]='h00001f7f;
    rd_cycle[ 4787] = 1'b0;  wr_cycle[ 4787] = 1'b1;  addr_rom[ 4787]='h00003e50;  wr_data_rom[ 4787]='h00001c10;
    rd_cycle[ 4788] = 1'b0;  wr_cycle[ 4788] = 1'b1;  addr_rom[ 4788]='h000025f4;  wr_data_rom[ 4788]='h00001eb2;
    rd_cycle[ 4789] = 1'b1;  wr_cycle[ 4789] = 1'b0;  addr_rom[ 4789]='h00003018;  wr_data_rom[ 4789]='h00000000;
    rd_cycle[ 4790] = 1'b0;  wr_cycle[ 4790] = 1'b1;  addr_rom[ 4790]='h000013b0;  wr_data_rom[ 4790]='h00002f1a;
    rd_cycle[ 4791] = 1'b1;  wr_cycle[ 4791] = 1'b0;  addr_rom[ 4791]='h00001250;  wr_data_rom[ 4791]='h00000000;
    rd_cycle[ 4792] = 1'b1;  wr_cycle[ 4792] = 1'b0;  addr_rom[ 4792]='h00003ad8;  wr_data_rom[ 4792]='h00000000;
    rd_cycle[ 4793] = 1'b0;  wr_cycle[ 4793] = 1'b1;  addr_rom[ 4793]='h000015a0;  wr_data_rom[ 4793]='h00003b3d;
    rd_cycle[ 4794] = 1'b0;  wr_cycle[ 4794] = 1'b1;  addr_rom[ 4794]='h00003134;  wr_data_rom[ 4794]='h00001d1f;
    rd_cycle[ 4795] = 1'b1;  wr_cycle[ 4795] = 1'b0;  addr_rom[ 4795]='h000022a4;  wr_data_rom[ 4795]='h00000000;
    rd_cycle[ 4796] = 1'b1;  wr_cycle[ 4796] = 1'b0;  addr_rom[ 4796]='h00002dcc;  wr_data_rom[ 4796]='h00000000;
    rd_cycle[ 4797] = 1'b1;  wr_cycle[ 4797] = 1'b0;  addr_rom[ 4797]='h00000348;  wr_data_rom[ 4797]='h00000000;
    rd_cycle[ 4798] = 1'b0;  wr_cycle[ 4798] = 1'b1;  addr_rom[ 4798]='h00002474;  wr_data_rom[ 4798]='h00002a85;
    rd_cycle[ 4799] = 1'b0;  wr_cycle[ 4799] = 1'b1;  addr_rom[ 4799]='h00000700;  wr_data_rom[ 4799]='h00000bc8;
    rd_cycle[ 4800] = 1'b1;  wr_cycle[ 4800] = 1'b0;  addr_rom[ 4800]='h000022e0;  wr_data_rom[ 4800]='h00000000;
    rd_cycle[ 4801] = 1'b1;  wr_cycle[ 4801] = 1'b0;  addr_rom[ 4801]='h00000500;  wr_data_rom[ 4801]='h00000000;
    rd_cycle[ 4802] = 1'b1;  wr_cycle[ 4802] = 1'b0;  addr_rom[ 4802]='h00002080;  wr_data_rom[ 4802]='h00000000;
    rd_cycle[ 4803] = 1'b0;  wr_cycle[ 4803] = 1'b1;  addr_rom[ 4803]='h00003338;  wr_data_rom[ 4803]='h00003a8c;
    rd_cycle[ 4804] = 1'b0;  wr_cycle[ 4804] = 1'b1;  addr_rom[ 4804]='h00000e18;  wr_data_rom[ 4804]='h000003ff;
    rd_cycle[ 4805] = 1'b1;  wr_cycle[ 4805] = 1'b0;  addr_rom[ 4805]='h000003ec;  wr_data_rom[ 4805]='h00000000;
    rd_cycle[ 4806] = 1'b0;  wr_cycle[ 4806] = 1'b1;  addr_rom[ 4806]='h0000213c;  wr_data_rom[ 4806]='h00002f23;
    rd_cycle[ 4807] = 1'b0;  wr_cycle[ 4807] = 1'b1;  addr_rom[ 4807]='h00003d8c;  wr_data_rom[ 4807]='h000010ba;
    rd_cycle[ 4808] = 1'b0;  wr_cycle[ 4808] = 1'b1;  addr_rom[ 4808]='h00000f54;  wr_data_rom[ 4808]='h000005d9;
    rd_cycle[ 4809] = 1'b0;  wr_cycle[ 4809] = 1'b1;  addr_rom[ 4809]='h000001d0;  wr_data_rom[ 4809]='h000008fc;
    rd_cycle[ 4810] = 1'b0;  wr_cycle[ 4810] = 1'b1;  addr_rom[ 4810]='h00002fa4;  wr_data_rom[ 4810]='h00000a8c;
    rd_cycle[ 4811] = 1'b1;  wr_cycle[ 4811] = 1'b0;  addr_rom[ 4811]='h000034f8;  wr_data_rom[ 4811]='h00000000;
    rd_cycle[ 4812] = 1'b1;  wr_cycle[ 4812] = 1'b0;  addr_rom[ 4812]='h000008b0;  wr_data_rom[ 4812]='h00000000;
    rd_cycle[ 4813] = 1'b1;  wr_cycle[ 4813] = 1'b0;  addr_rom[ 4813]='h000032d8;  wr_data_rom[ 4813]='h00000000;
    rd_cycle[ 4814] = 1'b1;  wr_cycle[ 4814] = 1'b0;  addr_rom[ 4814]='h00000784;  wr_data_rom[ 4814]='h00000000;
    rd_cycle[ 4815] = 1'b1;  wr_cycle[ 4815] = 1'b0;  addr_rom[ 4815]='h000016a8;  wr_data_rom[ 4815]='h00000000;
    rd_cycle[ 4816] = 1'b1;  wr_cycle[ 4816] = 1'b0;  addr_rom[ 4816]='h000033c8;  wr_data_rom[ 4816]='h00000000;
    rd_cycle[ 4817] = 1'b1;  wr_cycle[ 4817] = 1'b0;  addr_rom[ 4817]='h00001704;  wr_data_rom[ 4817]='h00000000;
    rd_cycle[ 4818] = 1'b1;  wr_cycle[ 4818] = 1'b0;  addr_rom[ 4818]='h0000099c;  wr_data_rom[ 4818]='h00000000;
    rd_cycle[ 4819] = 1'b1;  wr_cycle[ 4819] = 1'b0;  addr_rom[ 4819]='h000037d0;  wr_data_rom[ 4819]='h00000000;
    rd_cycle[ 4820] = 1'b0;  wr_cycle[ 4820] = 1'b1;  addr_rom[ 4820]='h00001a90;  wr_data_rom[ 4820]='h0000397f;
    rd_cycle[ 4821] = 1'b0;  wr_cycle[ 4821] = 1'b1;  addr_rom[ 4821]='h00000014;  wr_data_rom[ 4821]='h000009dd;
    rd_cycle[ 4822] = 1'b1;  wr_cycle[ 4822] = 1'b0;  addr_rom[ 4822]='h00000a84;  wr_data_rom[ 4822]='h00000000;
    rd_cycle[ 4823] = 1'b1;  wr_cycle[ 4823] = 1'b0;  addr_rom[ 4823]='h0000173c;  wr_data_rom[ 4823]='h00000000;
    rd_cycle[ 4824] = 1'b0;  wr_cycle[ 4824] = 1'b1;  addr_rom[ 4824]='h000007b8;  wr_data_rom[ 4824]='h0000270e;
    rd_cycle[ 4825] = 1'b1;  wr_cycle[ 4825] = 1'b0;  addr_rom[ 4825]='h000000c0;  wr_data_rom[ 4825]='h00000000;
    rd_cycle[ 4826] = 1'b0;  wr_cycle[ 4826] = 1'b1;  addr_rom[ 4826]='h00000d8c;  wr_data_rom[ 4826]='h00002ac8;
    rd_cycle[ 4827] = 1'b1;  wr_cycle[ 4827] = 1'b0;  addr_rom[ 4827]='h00000a70;  wr_data_rom[ 4827]='h00000000;
    rd_cycle[ 4828] = 1'b1;  wr_cycle[ 4828] = 1'b0;  addr_rom[ 4828]='h00003d94;  wr_data_rom[ 4828]='h00000000;
    rd_cycle[ 4829] = 1'b1;  wr_cycle[ 4829] = 1'b0;  addr_rom[ 4829]='h0000198c;  wr_data_rom[ 4829]='h00000000;
    rd_cycle[ 4830] = 1'b1;  wr_cycle[ 4830] = 1'b0;  addr_rom[ 4830]='h00000914;  wr_data_rom[ 4830]='h00000000;
    rd_cycle[ 4831] = 1'b1;  wr_cycle[ 4831] = 1'b0;  addr_rom[ 4831]='h00003834;  wr_data_rom[ 4831]='h00000000;
    rd_cycle[ 4832] = 1'b1;  wr_cycle[ 4832] = 1'b0;  addr_rom[ 4832]='h00002250;  wr_data_rom[ 4832]='h00000000;
    rd_cycle[ 4833] = 1'b0;  wr_cycle[ 4833] = 1'b1;  addr_rom[ 4833]='h0000335c;  wr_data_rom[ 4833]='h0000303c;
    rd_cycle[ 4834] = 1'b0;  wr_cycle[ 4834] = 1'b1;  addr_rom[ 4834]='h0000327c;  wr_data_rom[ 4834]='h00000a02;
    rd_cycle[ 4835] = 1'b1;  wr_cycle[ 4835] = 1'b0;  addr_rom[ 4835]='h00000c54;  wr_data_rom[ 4835]='h00000000;
    rd_cycle[ 4836] = 1'b0;  wr_cycle[ 4836] = 1'b1;  addr_rom[ 4836]='h000025d4;  wr_data_rom[ 4836]='h000011e2;
    rd_cycle[ 4837] = 1'b1;  wr_cycle[ 4837] = 1'b0;  addr_rom[ 4837]='h00002280;  wr_data_rom[ 4837]='h00000000;
    rd_cycle[ 4838] = 1'b1;  wr_cycle[ 4838] = 1'b0;  addr_rom[ 4838]='h00003828;  wr_data_rom[ 4838]='h00000000;
    rd_cycle[ 4839] = 1'b0;  wr_cycle[ 4839] = 1'b1;  addr_rom[ 4839]='h00002658;  wr_data_rom[ 4839]='h00003200;
    rd_cycle[ 4840] = 1'b0;  wr_cycle[ 4840] = 1'b1;  addr_rom[ 4840]='h0000148c;  wr_data_rom[ 4840]='h00002500;
    rd_cycle[ 4841] = 1'b0;  wr_cycle[ 4841] = 1'b1;  addr_rom[ 4841]='h00002968;  wr_data_rom[ 4841]='h00003385;
    rd_cycle[ 4842] = 1'b1;  wr_cycle[ 4842] = 1'b0;  addr_rom[ 4842]='h00002da8;  wr_data_rom[ 4842]='h00000000;
    rd_cycle[ 4843] = 1'b0;  wr_cycle[ 4843] = 1'b1;  addr_rom[ 4843]='h000019cc;  wr_data_rom[ 4843]='h000034e0;
    rd_cycle[ 4844] = 1'b0;  wr_cycle[ 4844] = 1'b1;  addr_rom[ 4844]='h00001e50;  wr_data_rom[ 4844]='h0000362a;
    rd_cycle[ 4845] = 1'b1;  wr_cycle[ 4845] = 1'b0;  addr_rom[ 4845]='h0000074c;  wr_data_rom[ 4845]='h00000000;
    rd_cycle[ 4846] = 1'b0;  wr_cycle[ 4846] = 1'b1;  addr_rom[ 4846]='h00000c34;  wr_data_rom[ 4846]='h00000795;
    rd_cycle[ 4847] = 1'b1;  wr_cycle[ 4847] = 1'b0;  addr_rom[ 4847]='h00000f74;  wr_data_rom[ 4847]='h00000000;
    rd_cycle[ 4848] = 1'b0;  wr_cycle[ 4848] = 1'b1;  addr_rom[ 4848]='h00001968;  wr_data_rom[ 4848]='h00000efb;
    rd_cycle[ 4849] = 1'b1;  wr_cycle[ 4849] = 1'b0;  addr_rom[ 4849]='h000024ac;  wr_data_rom[ 4849]='h00000000;
    rd_cycle[ 4850] = 1'b0;  wr_cycle[ 4850] = 1'b1;  addr_rom[ 4850]='h00002824;  wr_data_rom[ 4850]='h0000031b;
    rd_cycle[ 4851] = 1'b0;  wr_cycle[ 4851] = 1'b1;  addr_rom[ 4851]='h000035f8;  wr_data_rom[ 4851]='h000037d4;
    rd_cycle[ 4852] = 1'b0;  wr_cycle[ 4852] = 1'b1;  addr_rom[ 4852]='h000036fc;  wr_data_rom[ 4852]='h00000414;
    rd_cycle[ 4853] = 1'b1;  wr_cycle[ 4853] = 1'b0;  addr_rom[ 4853]='h00001724;  wr_data_rom[ 4853]='h00000000;
    rd_cycle[ 4854] = 1'b0;  wr_cycle[ 4854] = 1'b1;  addr_rom[ 4854]='h00002cb0;  wr_data_rom[ 4854]='h00002331;
    rd_cycle[ 4855] = 1'b0;  wr_cycle[ 4855] = 1'b1;  addr_rom[ 4855]='h000006f4;  wr_data_rom[ 4855]='h0000109e;
    rd_cycle[ 4856] = 1'b0;  wr_cycle[ 4856] = 1'b1;  addr_rom[ 4856]='h00002844;  wr_data_rom[ 4856]='h000032b3;
    rd_cycle[ 4857] = 1'b0;  wr_cycle[ 4857] = 1'b1;  addr_rom[ 4857]='h00003954;  wr_data_rom[ 4857]='h00000f1e;
    rd_cycle[ 4858] = 1'b0;  wr_cycle[ 4858] = 1'b1;  addr_rom[ 4858]='h00000c60;  wr_data_rom[ 4858]='h000030ee;
    rd_cycle[ 4859] = 1'b1;  wr_cycle[ 4859] = 1'b0;  addr_rom[ 4859]='h00000828;  wr_data_rom[ 4859]='h00000000;
    rd_cycle[ 4860] = 1'b0;  wr_cycle[ 4860] = 1'b1;  addr_rom[ 4860]='h00000530;  wr_data_rom[ 4860]='h00000aee;
    rd_cycle[ 4861] = 1'b0;  wr_cycle[ 4861] = 1'b1;  addr_rom[ 4861]='h00000930;  wr_data_rom[ 4861]='h00003a6f;
    rd_cycle[ 4862] = 1'b0;  wr_cycle[ 4862] = 1'b1;  addr_rom[ 4862]='h0000025c;  wr_data_rom[ 4862]='h00001f54;
    rd_cycle[ 4863] = 1'b0;  wr_cycle[ 4863] = 1'b1;  addr_rom[ 4863]='h00002698;  wr_data_rom[ 4863]='h00003403;
    rd_cycle[ 4864] = 1'b1;  wr_cycle[ 4864] = 1'b0;  addr_rom[ 4864]='h00001340;  wr_data_rom[ 4864]='h00000000;
    rd_cycle[ 4865] = 1'b0;  wr_cycle[ 4865] = 1'b1;  addr_rom[ 4865]='h00003e54;  wr_data_rom[ 4865]='h000029e4;
    rd_cycle[ 4866] = 1'b0;  wr_cycle[ 4866] = 1'b1;  addr_rom[ 4866]='h00002410;  wr_data_rom[ 4866]='h00003ee2;
    rd_cycle[ 4867] = 1'b0;  wr_cycle[ 4867] = 1'b1;  addr_rom[ 4867]='h00001700;  wr_data_rom[ 4867]='h00003de1;
    rd_cycle[ 4868] = 1'b0;  wr_cycle[ 4868] = 1'b1;  addr_rom[ 4868]='h00000824;  wr_data_rom[ 4868]='h00000ad4;
    rd_cycle[ 4869] = 1'b0;  wr_cycle[ 4869] = 1'b1;  addr_rom[ 4869]='h00001910;  wr_data_rom[ 4869]='h0000074b;
    rd_cycle[ 4870] = 1'b0;  wr_cycle[ 4870] = 1'b1;  addr_rom[ 4870]='h00001c54;  wr_data_rom[ 4870]='h00001f6a;
    rd_cycle[ 4871] = 1'b0;  wr_cycle[ 4871] = 1'b1;  addr_rom[ 4871]='h00003b50;  wr_data_rom[ 4871]='h00002ae5;
    rd_cycle[ 4872] = 1'b1;  wr_cycle[ 4872] = 1'b0;  addr_rom[ 4872]='h00002a70;  wr_data_rom[ 4872]='h00000000;
    rd_cycle[ 4873] = 1'b0;  wr_cycle[ 4873] = 1'b1;  addr_rom[ 4873]='h000036ac;  wr_data_rom[ 4873]='h0000011b;
    rd_cycle[ 4874] = 1'b1;  wr_cycle[ 4874] = 1'b0;  addr_rom[ 4874]='h000000cc;  wr_data_rom[ 4874]='h00000000;
    rd_cycle[ 4875] = 1'b0;  wr_cycle[ 4875] = 1'b1;  addr_rom[ 4875]='h00001878;  wr_data_rom[ 4875]='h0000152d;
    rd_cycle[ 4876] = 1'b0;  wr_cycle[ 4876] = 1'b1;  addr_rom[ 4876]='h00002624;  wr_data_rom[ 4876]='h00001c17;
    rd_cycle[ 4877] = 1'b0;  wr_cycle[ 4877] = 1'b1;  addr_rom[ 4877]='h000027a8;  wr_data_rom[ 4877]='h0000311a;
    rd_cycle[ 4878] = 1'b1;  wr_cycle[ 4878] = 1'b0;  addr_rom[ 4878]='h00001d00;  wr_data_rom[ 4878]='h00000000;
    rd_cycle[ 4879] = 1'b1;  wr_cycle[ 4879] = 1'b0;  addr_rom[ 4879]='h0000274c;  wr_data_rom[ 4879]='h00000000;
    rd_cycle[ 4880] = 1'b1;  wr_cycle[ 4880] = 1'b0;  addr_rom[ 4880]='h00001000;  wr_data_rom[ 4880]='h00000000;
    rd_cycle[ 4881] = 1'b0;  wr_cycle[ 4881] = 1'b1;  addr_rom[ 4881]='h00003860;  wr_data_rom[ 4881]='h00003494;
    rd_cycle[ 4882] = 1'b0;  wr_cycle[ 4882] = 1'b1;  addr_rom[ 4882]='h00000b94;  wr_data_rom[ 4882]='h0000108a;
    rd_cycle[ 4883] = 1'b0;  wr_cycle[ 4883] = 1'b1;  addr_rom[ 4883]='h00003ee0;  wr_data_rom[ 4883]='h0000061a;
    rd_cycle[ 4884] = 1'b0;  wr_cycle[ 4884] = 1'b1;  addr_rom[ 4884]='h00001b74;  wr_data_rom[ 4884]='h000028c8;
    rd_cycle[ 4885] = 1'b1;  wr_cycle[ 4885] = 1'b0;  addr_rom[ 4885]='h00000af0;  wr_data_rom[ 4885]='h00000000;
    rd_cycle[ 4886] = 1'b0;  wr_cycle[ 4886] = 1'b1;  addr_rom[ 4886]='h00001b78;  wr_data_rom[ 4886]='h00002d28;
    rd_cycle[ 4887] = 1'b0;  wr_cycle[ 4887] = 1'b1;  addr_rom[ 4887]='h000006dc;  wr_data_rom[ 4887]='h00001946;
    rd_cycle[ 4888] = 1'b1;  wr_cycle[ 4888] = 1'b0;  addr_rom[ 4888]='h00002364;  wr_data_rom[ 4888]='h00000000;
    rd_cycle[ 4889] = 1'b0;  wr_cycle[ 4889] = 1'b1;  addr_rom[ 4889]='h00000730;  wr_data_rom[ 4889]='h0000342a;
    rd_cycle[ 4890] = 1'b1;  wr_cycle[ 4890] = 1'b0;  addr_rom[ 4890]='h00003708;  wr_data_rom[ 4890]='h00000000;
    rd_cycle[ 4891] = 1'b0;  wr_cycle[ 4891] = 1'b1;  addr_rom[ 4891]='h00003fc0;  wr_data_rom[ 4891]='h000021e2;
    rd_cycle[ 4892] = 1'b1;  wr_cycle[ 4892] = 1'b0;  addr_rom[ 4892]='h00002ffc;  wr_data_rom[ 4892]='h00000000;
    rd_cycle[ 4893] = 1'b1;  wr_cycle[ 4893] = 1'b0;  addr_rom[ 4893]='h00002d00;  wr_data_rom[ 4893]='h00000000;
    rd_cycle[ 4894] = 1'b0;  wr_cycle[ 4894] = 1'b1;  addr_rom[ 4894]='h00002d18;  wr_data_rom[ 4894]='h000015d7;
    rd_cycle[ 4895] = 1'b1;  wr_cycle[ 4895] = 1'b0;  addr_rom[ 4895]='h00002d54;  wr_data_rom[ 4895]='h00000000;
    rd_cycle[ 4896] = 1'b1;  wr_cycle[ 4896] = 1'b0;  addr_rom[ 4896]='h00002fe4;  wr_data_rom[ 4896]='h00000000;
    rd_cycle[ 4897] = 1'b0;  wr_cycle[ 4897] = 1'b1;  addr_rom[ 4897]='h00002028;  wr_data_rom[ 4897]='h0000078f;
    rd_cycle[ 4898] = 1'b0;  wr_cycle[ 4898] = 1'b1;  addr_rom[ 4898]='h00003ca8;  wr_data_rom[ 4898]='h00000921;
    rd_cycle[ 4899] = 1'b0;  wr_cycle[ 4899] = 1'b1;  addr_rom[ 4899]='h00003a30;  wr_data_rom[ 4899]='h00000fb4;
    rd_cycle[ 4900] = 1'b0;  wr_cycle[ 4900] = 1'b1;  addr_rom[ 4900]='h00001e90;  wr_data_rom[ 4900]='h0000049a;
    rd_cycle[ 4901] = 1'b1;  wr_cycle[ 4901] = 1'b0;  addr_rom[ 4901]='h00001b58;  wr_data_rom[ 4901]='h00000000;
    rd_cycle[ 4902] = 1'b1;  wr_cycle[ 4902] = 1'b0;  addr_rom[ 4902]='h00003c00;  wr_data_rom[ 4902]='h00000000;
    rd_cycle[ 4903] = 1'b1;  wr_cycle[ 4903] = 1'b0;  addr_rom[ 4903]='h00001610;  wr_data_rom[ 4903]='h00000000;
    rd_cycle[ 4904] = 1'b1;  wr_cycle[ 4904] = 1'b0;  addr_rom[ 4904]='h00003ccc;  wr_data_rom[ 4904]='h00000000;
    rd_cycle[ 4905] = 1'b0;  wr_cycle[ 4905] = 1'b1;  addr_rom[ 4905]='h000029d0;  wr_data_rom[ 4905]='h000033f8;
    rd_cycle[ 4906] = 1'b1;  wr_cycle[ 4906] = 1'b0;  addr_rom[ 4906]='h00001768;  wr_data_rom[ 4906]='h00000000;
    rd_cycle[ 4907] = 1'b0;  wr_cycle[ 4907] = 1'b1;  addr_rom[ 4907]='h00003b64;  wr_data_rom[ 4907]='h00001e1f;
    rd_cycle[ 4908] = 1'b0;  wr_cycle[ 4908] = 1'b1;  addr_rom[ 4908]='h000014c8;  wr_data_rom[ 4908]='h0000054c;
    rd_cycle[ 4909] = 1'b0;  wr_cycle[ 4909] = 1'b1;  addr_rom[ 4909]='h000030e4;  wr_data_rom[ 4909]='h00002082;
    rd_cycle[ 4910] = 1'b1;  wr_cycle[ 4910] = 1'b0;  addr_rom[ 4910]='h00002da8;  wr_data_rom[ 4910]='h00000000;
    rd_cycle[ 4911] = 1'b0;  wr_cycle[ 4911] = 1'b1;  addr_rom[ 4911]='h00002180;  wr_data_rom[ 4911]='h00003cb1;
    rd_cycle[ 4912] = 1'b0;  wr_cycle[ 4912] = 1'b1;  addr_rom[ 4912]='h00000894;  wr_data_rom[ 4912]='h00003fc8;
    rd_cycle[ 4913] = 1'b1;  wr_cycle[ 4913] = 1'b0;  addr_rom[ 4913]='h000012a0;  wr_data_rom[ 4913]='h00000000;
    rd_cycle[ 4914] = 1'b0;  wr_cycle[ 4914] = 1'b1;  addr_rom[ 4914]='h000004dc;  wr_data_rom[ 4914]='h00001e12;
    rd_cycle[ 4915] = 1'b0;  wr_cycle[ 4915] = 1'b1;  addr_rom[ 4915]='h00002938;  wr_data_rom[ 4915]='h000012ea;
    rd_cycle[ 4916] = 1'b1;  wr_cycle[ 4916] = 1'b0;  addr_rom[ 4916]='h000011f4;  wr_data_rom[ 4916]='h00000000;
    rd_cycle[ 4917] = 1'b1;  wr_cycle[ 4917] = 1'b0;  addr_rom[ 4917]='h00000910;  wr_data_rom[ 4917]='h00000000;
    rd_cycle[ 4918] = 1'b1;  wr_cycle[ 4918] = 1'b0;  addr_rom[ 4918]='h00002630;  wr_data_rom[ 4918]='h00000000;
    rd_cycle[ 4919] = 1'b0;  wr_cycle[ 4919] = 1'b1;  addr_rom[ 4919]='h00000eac;  wr_data_rom[ 4919]='h00001f29;
    rd_cycle[ 4920] = 1'b1;  wr_cycle[ 4920] = 1'b0;  addr_rom[ 4920]='h00002848;  wr_data_rom[ 4920]='h00000000;
    rd_cycle[ 4921] = 1'b0;  wr_cycle[ 4921] = 1'b1;  addr_rom[ 4921]='h00003014;  wr_data_rom[ 4921]='h000019ed;
    rd_cycle[ 4922] = 1'b0;  wr_cycle[ 4922] = 1'b1;  addr_rom[ 4922]='h00001d5c;  wr_data_rom[ 4922]='h00001b9c;
    rd_cycle[ 4923] = 1'b0;  wr_cycle[ 4923] = 1'b1;  addr_rom[ 4923]='h00001600;  wr_data_rom[ 4923]='h00002e63;
    rd_cycle[ 4924] = 1'b0;  wr_cycle[ 4924] = 1'b1;  addr_rom[ 4924]='h00003b6c;  wr_data_rom[ 4924]='h000015ca;
    rd_cycle[ 4925] = 1'b0;  wr_cycle[ 4925] = 1'b1;  addr_rom[ 4925]='h00003cac;  wr_data_rom[ 4925]='h00001e75;
    rd_cycle[ 4926] = 1'b1;  wr_cycle[ 4926] = 1'b0;  addr_rom[ 4926]='h00003794;  wr_data_rom[ 4926]='h00000000;
    rd_cycle[ 4927] = 1'b1;  wr_cycle[ 4927] = 1'b0;  addr_rom[ 4927]='h00002a08;  wr_data_rom[ 4927]='h00000000;
    rd_cycle[ 4928] = 1'b0;  wr_cycle[ 4928] = 1'b1;  addr_rom[ 4928]='h00000ee8;  wr_data_rom[ 4928]='h00000017;
    rd_cycle[ 4929] = 1'b0;  wr_cycle[ 4929] = 1'b1;  addr_rom[ 4929]='h000016a4;  wr_data_rom[ 4929]='h00001199;
    rd_cycle[ 4930] = 1'b1;  wr_cycle[ 4930] = 1'b0;  addr_rom[ 4930]='h00001d18;  wr_data_rom[ 4930]='h00000000;
    rd_cycle[ 4931] = 1'b1;  wr_cycle[ 4931] = 1'b0;  addr_rom[ 4931]='h00001f40;  wr_data_rom[ 4931]='h00000000;
    rd_cycle[ 4932] = 1'b1;  wr_cycle[ 4932] = 1'b0;  addr_rom[ 4932]='h00003004;  wr_data_rom[ 4932]='h00000000;
    rd_cycle[ 4933] = 1'b1;  wr_cycle[ 4933] = 1'b0;  addr_rom[ 4933]='h00001d34;  wr_data_rom[ 4933]='h00000000;
    rd_cycle[ 4934] = 1'b1;  wr_cycle[ 4934] = 1'b0;  addr_rom[ 4934]='h00000438;  wr_data_rom[ 4934]='h00000000;
    rd_cycle[ 4935] = 1'b1;  wr_cycle[ 4935] = 1'b0;  addr_rom[ 4935]='h00001810;  wr_data_rom[ 4935]='h00000000;
    rd_cycle[ 4936] = 1'b1;  wr_cycle[ 4936] = 1'b0;  addr_rom[ 4936]='h00001fb8;  wr_data_rom[ 4936]='h00000000;
    rd_cycle[ 4937] = 1'b1;  wr_cycle[ 4937] = 1'b0;  addr_rom[ 4937]='h00002210;  wr_data_rom[ 4937]='h00000000;
    rd_cycle[ 4938] = 1'b1;  wr_cycle[ 4938] = 1'b0;  addr_rom[ 4938]='h00000774;  wr_data_rom[ 4938]='h00000000;
    rd_cycle[ 4939] = 1'b0;  wr_cycle[ 4939] = 1'b1;  addr_rom[ 4939]='h00003074;  wr_data_rom[ 4939]='h000020b2;
    rd_cycle[ 4940] = 1'b0;  wr_cycle[ 4940] = 1'b1;  addr_rom[ 4940]='h00000910;  wr_data_rom[ 4940]='h00003747;
    rd_cycle[ 4941] = 1'b1;  wr_cycle[ 4941] = 1'b0;  addr_rom[ 4941]='h000021b4;  wr_data_rom[ 4941]='h00000000;
    rd_cycle[ 4942] = 1'b1;  wr_cycle[ 4942] = 1'b0;  addr_rom[ 4942]='h00002eac;  wr_data_rom[ 4942]='h00000000;
    rd_cycle[ 4943] = 1'b0;  wr_cycle[ 4943] = 1'b1;  addr_rom[ 4943]='h00001194;  wr_data_rom[ 4943]='h0000101a;
    rd_cycle[ 4944] = 1'b1;  wr_cycle[ 4944] = 1'b0;  addr_rom[ 4944]='h00000ee8;  wr_data_rom[ 4944]='h00000000;
    rd_cycle[ 4945] = 1'b1;  wr_cycle[ 4945] = 1'b0;  addr_rom[ 4945]='h000001fc;  wr_data_rom[ 4945]='h00000000;
    rd_cycle[ 4946] = 1'b0;  wr_cycle[ 4946] = 1'b1;  addr_rom[ 4946]='h00002d3c;  wr_data_rom[ 4946]='h00002d1a;
    rd_cycle[ 4947] = 1'b0;  wr_cycle[ 4947] = 1'b1;  addr_rom[ 4947]='h00002e70;  wr_data_rom[ 4947]='h00001d3c;
    rd_cycle[ 4948] = 1'b0;  wr_cycle[ 4948] = 1'b1;  addr_rom[ 4948]='h00003f24;  wr_data_rom[ 4948]='h00002eba;
    rd_cycle[ 4949] = 1'b0;  wr_cycle[ 4949] = 1'b1;  addr_rom[ 4949]='h000035c0;  wr_data_rom[ 4949]='h000039f4;
    rd_cycle[ 4950] = 1'b0;  wr_cycle[ 4950] = 1'b1;  addr_rom[ 4950]='h00002c2c;  wr_data_rom[ 4950]='h000009ee;
    rd_cycle[ 4951] = 1'b0;  wr_cycle[ 4951] = 1'b1;  addr_rom[ 4951]='h00003b08;  wr_data_rom[ 4951]='h000025b0;
    rd_cycle[ 4952] = 1'b0;  wr_cycle[ 4952] = 1'b1;  addr_rom[ 4952]='h0000046c;  wr_data_rom[ 4952]='h00000f26;
    rd_cycle[ 4953] = 1'b1;  wr_cycle[ 4953] = 1'b0;  addr_rom[ 4953]='h00003c14;  wr_data_rom[ 4953]='h00000000;
    rd_cycle[ 4954] = 1'b1;  wr_cycle[ 4954] = 1'b0;  addr_rom[ 4954]='h00000628;  wr_data_rom[ 4954]='h00000000;
    rd_cycle[ 4955] = 1'b0;  wr_cycle[ 4955] = 1'b1;  addr_rom[ 4955]='h00000ee8;  wr_data_rom[ 4955]='h00000abb;
    rd_cycle[ 4956] = 1'b1;  wr_cycle[ 4956] = 1'b0;  addr_rom[ 4956]='h00000ee0;  wr_data_rom[ 4956]='h00000000;
    rd_cycle[ 4957] = 1'b1;  wr_cycle[ 4957] = 1'b0;  addr_rom[ 4957]='h00001fc4;  wr_data_rom[ 4957]='h00000000;
    rd_cycle[ 4958] = 1'b1;  wr_cycle[ 4958] = 1'b0;  addr_rom[ 4958]='h000037e0;  wr_data_rom[ 4958]='h00000000;
    rd_cycle[ 4959] = 1'b0;  wr_cycle[ 4959] = 1'b1;  addr_rom[ 4959]='h00003198;  wr_data_rom[ 4959]='h00003a61;
    rd_cycle[ 4960] = 1'b1;  wr_cycle[ 4960] = 1'b0;  addr_rom[ 4960]='h00001724;  wr_data_rom[ 4960]='h00000000;
    rd_cycle[ 4961] = 1'b0;  wr_cycle[ 4961] = 1'b1;  addr_rom[ 4961]='h00003164;  wr_data_rom[ 4961]='h00002008;
    rd_cycle[ 4962] = 1'b1;  wr_cycle[ 4962] = 1'b0;  addr_rom[ 4962]='h00003928;  wr_data_rom[ 4962]='h00000000;
    rd_cycle[ 4963] = 1'b1;  wr_cycle[ 4963] = 1'b0;  addr_rom[ 4963]='h00002bf4;  wr_data_rom[ 4963]='h00000000;
    rd_cycle[ 4964] = 1'b0;  wr_cycle[ 4964] = 1'b1;  addr_rom[ 4964]='h000011f0;  wr_data_rom[ 4964]='h0000379b;
    rd_cycle[ 4965] = 1'b0;  wr_cycle[ 4965] = 1'b1;  addr_rom[ 4965]='h00002018;  wr_data_rom[ 4965]='h00003554;
    rd_cycle[ 4966] = 1'b1;  wr_cycle[ 4966] = 1'b0;  addr_rom[ 4966]='h0000066c;  wr_data_rom[ 4966]='h00000000;
    rd_cycle[ 4967] = 1'b1;  wr_cycle[ 4967] = 1'b0;  addr_rom[ 4967]='h00002910;  wr_data_rom[ 4967]='h00000000;
    rd_cycle[ 4968] = 1'b1;  wr_cycle[ 4968] = 1'b0;  addr_rom[ 4968]='h0000393c;  wr_data_rom[ 4968]='h00000000;
    rd_cycle[ 4969] = 1'b1;  wr_cycle[ 4969] = 1'b0;  addr_rom[ 4969]='h00003edc;  wr_data_rom[ 4969]='h00000000;
    rd_cycle[ 4970] = 1'b0;  wr_cycle[ 4970] = 1'b1;  addr_rom[ 4970]='h00002ec0;  wr_data_rom[ 4970]='h00002874;
    rd_cycle[ 4971] = 1'b1;  wr_cycle[ 4971] = 1'b0;  addr_rom[ 4971]='h00000840;  wr_data_rom[ 4971]='h00000000;
    rd_cycle[ 4972] = 1'b0;  wr_cycle[ 4972] = 1'b1;  addr_rom[ 4972]='h0000146c;  wr_data_rom[ 4972]='h00003b5a;
    rd_cycle[ 4973] = 1'b1;  wr_cycle[ 4973] = 1'b0;  addr_rom[ 4973]='h00001a58;  wr_data_rom[ 4973]='h00000000;
    rd_cycle[ 4974] = 1'b0;  wr_cycle[ 4974] = 1'b1;  addr_rom[ 4974]='h0000371c;  wr_data_rom[ 4974]='h000004d1;
    rd_cycle[ 4975] = 1'b0;  wr_cycle[ 4975] = 1'b1;  addr_rom[ 4975]='h0000047c;  wr_data_rom[ 4975]='h000013da;
    rd_cycle[ 4976] = 1'b0;  wr_cycle[ 4976] = 1'b1;  addr_rom[ 4976]='h000016e0;  wr_data_rom[ 4976]='h00003d06;
    rd_cycle[ 4977] = 1'b1;  wr_cycle[ 4977] = 1'b0;  addr_rom[ 4977]='h000017ac;  wr_data_rom[ 4977]='h00000000;
    rd_cycle[ 4978] = 1'b1;  wr_cycle[ 4978] = 1'b0;  addr_rom[ 4978]='h0000223c;  wr_data_rom[ 4978]='h00000000;
    rd_cycle[ 4979] = 1'b0;  wr_cycle[ 4979] = 1'b1;  addr_rom[ 4979]='h00001b7c;  wr_data_rom[ 4979]='h00003ec4;
    rd_cycle[ 4980] = 1'b1;  wr_cycle[ 4980] = 1'b0;  addr_rom[ 4980]='h00002bd4;  wr_data_rom[ 4980]='h00000000;
    rd_cycle[ 4981] = 1'b1;  wr_cycle[ 4981] = 1'b0;  addr_rom[ 4981]='h0000196c;  wr_data_rom[ 4981]='h00000000;
    rd_cycle[ 4982] = 1'b0;  wr_cycle[ 4982] = 1'b1;  addr_rom[ 4982]='h00000b98;  wr_data_rom[ 4982]='h00002133;
    rd_cycle[ 4983] = 1'b1;  wr_cycle[ 4983] = 1'b0;  addr_rom[ 4983]='h00001334;  wr_data_rom[ 4983]='h00000000;
    rd_cycle[ 4984] = 1'b1;  wr_cycle[ 4984] = 1'b0;  addr_rom[ 4984]='h000018ac;  wr_data_rom[ 4984]='h00000000;
    rd_cycle[ 4985] = 1'b0;  wr_cycle[ 4985] = 1'b1;  addr_rom[ 4985]='h000030b4;  wr_data_rom[ 4985]='h00002600;
    rd_cycle[ 4986] = 1'b1;  wr_cycle[ 4986] = 1'b0;  addr_rom[ 4986]='h00000944;  wr_data_rom[ 4986]='h00000000;
    rd_cycle[ 4987] = 1'b0;  wr_cycle[ 4987] = 1'b1;  addr_rom[ 4987]='h00001f70;  wr_data_rom[ 4987]='h00001f9b;
    rd_cycle[ 4988] = 1'b1;  wr_cycle[ 4988] = 1'b0;  addr_rom[ 4988]='h00001ee4;  wr_data_rom[ 4988]='h00000000;
    rd_cycle[ 4989] = 1'b1;  wr_cycle[ 4989] = 1'b0;  addr_rom[ 4989]='h00000598;  wr_data_rom[ 4989]='h00000000;
    rd_cycle[ 4990] = 1'b0;  wr_cycle[ 4990] = 1'b1;  addr_rom[ 4990]='h0000051c;  wr_data_rom[ 4990]='h000020db;
    rd_cycle[ 4991] = 1'b0;  wr_cycle[ 4991] = 1'b1;  addr_rom[ 4991]='h00000d58;  wr_data_rom[ 4991]='h000035f1;
    rd_cycle[ 4992] = 1'b1;  wr_cycle[ 4992] = 1'b0;  addr_rom[ 4992]='h00002bac;  wr_data_rom[ 4992]='h00000000;
    rd_cycle[ 4993] = 1'b0;  wr_cycle[ 4993] = 1'b1;  addr_rom[ 4993]='h000011c8;  wr_data_rom[ 4993]='h00001989;
    rd_cycle[ 4994] = 1'b0;  wr_cycle[ 4994] = 1'b1;  addr_rom[ 4994]='h00001510;  wr_data_rom[ 4994]='h00000e4f;
    rd_cycle[ 4995] = 1'b1;  wr_cycle[ 4995] = 1'b0;  addr_rom[ 4995]='h00002588;  wr_data_rom[ 4995]='h00000000;
    rd_cycle[ 4996] = 1'b0;  wr_cycle[ 4996] = 1'b1;  addr_rom[ 4996]='h000030f4;  wr_data_rom[ 4996]='h000032d9;
    rd_cycle[ 4997] = 1'b0;  wr_cycle[ 4997] = 1'b1;  addr_rom[ 4997]='h000032ac;  wr_data_rom[ 4997]='h000010f9;
    rd_cycle[ 4998] = 1'b0;  wr_cycle[ 4998] = 1'b1;  addr_rom[ 4998]='h000014c8;  wr_data_rom[ 4998]='h000035c1;
    rd_cycle[ 4999] = 1'b1;  wr_cycle[ 4999] = 1'b0;  addr_rom[ 4999]='h000038d8;  wr_data_rom[ 4999]='h00000000;
    rd_cycle[ 5000] = 1'b0;  wr_cycle[ 5000] = 1'b1;  addr_rom[ 5000]='h00001800;  wr_data_rom[ 5000]='h0000259c;
    rd_cycle[ 5001] = 1'b1;  wr_cycle[ 5001] = 1'b0;  addr_rom[ 5001]='h000003b4;  wr_data_rom[ 5001]='h00000000;
    rd_cycle[ 5002] = 1'b1;  wr_cycle[ 5002] = 1'b0;  addr_rom[ 5002]='h000024e4;  wr_data_rom[ 5002]='h00000000;
    rd_cycle[ 5003] = 1'b1;  wr_cycle[ 5003] = 1'b0;  addr_rom[ 5003]='h0000355c;  wr_data_rom[ 5003]='h00000000;
    rd_cycle[ 5004] = 1'b0;  wr_cycle[ 5004] = 1'b1;  addr_rom[ 5004]='h000008e8;  wr_data_rom[ 5004]='h00002d83;
    rd_cycle[ 5005] = 1'b0;  wr_cycle[ 5005] = 1'b1;  addr_rom[ 5005]='h000036e4;  wr_data_rom[ 5005]='h00003c4e;
    rd_cycle[ 5006] = 1'b0;  wr_cycle[ 5006] = 1'b1;  addr_rom[ 5006]='h0000324c;  wr_data_rom[ 5006]='h0000146a;
    rd_cycle[ 5007] = 1'b1;  wr_cycle[ 5007] = 1'b0;  addr_rom[ 5007]='h00001870;  wr_data_rom[ 5007]='h00000000;
    rd_cycle[ 5008] = 1'b1;  wr_cycle[ 5008] = 1'b0;  addr_rom[ 5008]='h000033f0;  wr_data_rom[ 5008]='h00000000;
    rd_cycle[ 5009] = 1'b0;  wr_cycle[ 5009] = 1'b1;  addr_rom[ 5009]='h0000065c;  wr_data_rom[ 5009]='h00002d34;
    rd_cycle[ 5010] = 1'b0;  wr_cycle[ 5010] = 1'b1;  addr_rom[ 5010]='h00000648;  wr_data_rom[ 5010]='h00000c7e;
    rd_cycle[ 5011] = 1'b1;  wr_cycle[ 5011] = 1'b0;  addr_rom[ 5011]='h00000530;  wr_data_rom[ 5011]='h00000000;
    rd_cycle[ 5012] = 1'b1;  wr_cycle[ 5012] = 1'b0;  addr_rom[ 5012]='h00000414;  wr_data_rom[ 5012]='h00000000;
    rd_cycle[ 5013] = 1'b0;  wr_cycle[ 5013] = 1'b1;  addr_rom[ 5013]='h00000e58;  wr_data_rom[ 5013]='h00001fed;
    rd_cycle[ 5014] = 1'b0;  wr_cycle[ 5014] = 1'b1;  addr_rom[ 5014]='h00001158;  wr_data_rom[ 5014]='h00001a56;
    rd_cycle[ 5015] = 1'b1;  wr_cycle[ 5015] = 1'b0;  addr_rom[ 5015]='h00002074;  wr_data_rom[ 5015]='h00000000;
    rd_cycle[ 5016] = 1'b0;  wr_cycle[ 5016] = 1'b1;  addr_rom[ 5016]='h0000397c;  wr_data_rom[ 5016]='h0000128f;
    rd_cycle[ 5017] = 1'b0;  wr_cycle[ 5017] = 1'b1;  addr_rom[ 5017]='h00003370;  wr_data_rom[ 5017]='h000001e2;
    rd_cycle[ 5018] = 1'b1;  wr_cycle[ 5018] = 1'b0;  addr_rom[ 5018]='h00000000;  wr_data_rom[ 5018]='h00000000;
    rd_cycle[ 5019] = 1'b1;  wr_cycle[ 5019] = 1'b0;  addr_rom[ 5019]='h00000444;  wr_data_rom[ 5019]='h00000000;
    rd_cycle[ 5020] = 1'b0;  wr_cycle[ 5020] = 1'b1;  addr_rom[ 5020]='h00000fa0;  wr_data_rom[ 5020]='h00000d26;
    rd_cycle[ 5021] = 1'b1;  wr_cycle[ 5021] = 1'b0;  addr_rom[ 5021]='h0000379c;  wr_data_rom[ 5021]='h00000000;
    rd_cycle[ 5022] = 1'b1;  wr_cycle[ 5022] = 1'b0;  addr_rom[ 5022]='h00000168;  wr_data_rom[ 5022]='h00000000;
    rd_cycle[ 5023] = 1'b0;  wr_cycle[ 5023] = 1'b1;  addr_rom[ 5023]='h00000b18;  wr_data_rom[ 5023]='h00001eb5;
    rd_cycle[ 5024] = 1'b1;  wr_cycle[ 5024] = 1'b0;  addr_rom[ 5024]='h00003770;  wr_data_rom[ 5024]='h00000000;
    rd_cycle[ 5025] = 1'b0;  wr_cycle[ 5025] = 1'b1;  addr_rom[ 5025]='h00003e20;  wr_data_rom[ 5025]='h00002def;
    rd_cycle[ 5026] = 1'b0;  wr_cycle[ 5026] = 1'b1;  addr_rom[ 5026]='h0000290c;  wr_data_rom[ 5026]='h000017c9;
    rd_cycle[ 5027] = 1'b1;  wr_cycle[ 5027] = 1'b0;  addr_rom[ 5027]='h000012bc;  wr_data_rom[ 5027]='h00000000;
    rd_cycle[ 5028] = 1'b1;  wr_cycle[ 5028] = 1'b0;  addr_rom[ 5028]='h0000221c;  wr_data_rom[ 5028]='h00000000;
    rd_cycle[ 5029] = 1'b1;  wr_cycle[ 5029] = 1'b0;  addr_rom[ 5029]='h00001ad0;  wr_data_rom[ 5029]='h00000000;
    rd_cycle[ 5030] = 1'b0;  wr_cycle[ 5030] = 1'b1;  addr_rom[ 5030]='h00000180;  wr_data_rom[ 5030]='h00003cf6;
    rd_cycle[ 5031] = 1'b1;  wr_cycle[ 5031] = 1'b0;  addr_rom[ 5031]='h00000ae4;  wr_data_rom[ 5031]='h00000000;
    rd_cycle[ 5032] = 1'b0;  wr_cycle[ 5032] = 1'b1;  addr_rom[ 5032]='h00002fd4;  wr_data_rom[ 5032]='h00002bb2;
    rd_cycle[ 5033] = 1'b0;  wr_cycle[ 5033] = 1'b1;  addr_rom[ 5033]='h00001f1c;  wr_data_rom[ 5033]='h00003714;
    rd_cycle[ 5034] = 1'b0;  wr_cycle[ 5034] = 1'b1;  addr_rom[ 5034]='h00003eec;  wr_data_rom[ 5034]='h00001af0;
    rd_cycle[ 5035] = 1'b0;  wr_cycle[ 5035] = 1'b1;  addr_rom[ 5035]='h000002c8;  wr_data_rom[ 5035]='h0000090c;
    rd_cycle[ 5036] = 1'b0;  wr_cycle[ 5036] = 1'b1;  addr_rom[ 5036]='h00003200;  wr_data_rom[ 5036]='h00001bfd;
    rd_cycle[ 5037] = 1'b0;  wr_cycle[ 5037] = 1'b1;  addr_rom[ 5037]='h00002a98;  wr_data_rom[ 5037]='h00000350;
    rd_cycle[ 5038] = 1'b1;  wr_cycle[ 5038] = 1'b0;  addr_rom[ 5038]='h00001b90;  wr_data_rom[ 5038]='h00000000;
    rd_cycle[ 5039] = 1'b1;  wr_cycle[ 5039] = 1'b0;  addr_rom[ 5039]='h00003c18;  wr_data_rom[ 5039]='h00000000;
    rd_cycle[ 5040] = 1'b0;  wr_cycle[ 5040] = 1'b1;  addr_rom[ 5040]='h00000d78;  wr_data_rom[ 5040]='h00001551;
    rd_cycle[ 5041] = 1'b0;  wr_cycle[ 5041] = 1'b1;  addr_rom[ 5041]='h00003a10;  wr_data_rom[ 5041]='h00002c24;
    rd_cycle[ 5042] = 1'b1;  wr_cycle[ 5042] = 1'b0;  addr_rom[ 5042]='h000001a8;  wr_data_rom[ 5042]='h00000000;
    rd_cycle[ 5043] = 1'b1;  wr_cycle[ 5043] = 1'b0;  addr_rom[ 5043]='h000036e0;  wr_data_rom[ 5043]='h00000000;
    rd_cycle[ 5044] = 1'b0;  wr_cycle[ 5044] = 1'b1;  addr_rom[ 5044]='h00002604;  wr_data_rom[ 5044]='h0000313e;
    rd_cycle[ 5045] = 1'b0;  wr_cycle[ 5045] = 1'b1;  addr_rom[ 5045]='h0000368c;  wr_data_rom[ 5045]='h000033d0;
    rd_cycle[ 5046] = 1'b0;  wr_cycle[ 5046] = 1'b1;  addr_rom[ 5046]='h00001900;  wr_data_rom[ 5046]='h00003189;
    rd_cycle[ 5047] = 1'b0;  wr_cycle[ 5047] = 1'b1;  addr_rom[ 5047]='h00003640;  wr_data_rom[ 5047]='h0000063b;
    rd_cycle[ 5048] = 1'b0;  wr_cycle[ 5048] = 1'b1;  addr_rom[ 5048]='h00003b14;  wr_data_rom[ 5048]='h00002cd9;
    rd_cycle[ 5049] = 1'b0;  wr_cycle[ 5049] = 1'b1;  addr_rom[ 5049]='h00000634;  wr_data_rom[ 5049]='h00000249;
    rd_cycle[ 5050] = 1'b0;  wr_cycle[ 5050] = 1'b1;  addr_rom[ 5050]='h00000f0c;  wr_data_rom[ 5050]='h000035da;
    rd_cycle[ 5051] = 1'b1;  wr_cycle[ 5051] = 1'b0;  addr_rom[ 5051]='h00000364;  wr_data_rom[ 5051]='h00000000;
    rd_cycle[ 5052] = 1'b0;  wr_cycle[ 5052] = 1'b1;  addr_rom[ 5052]='h0000036c;  wr_data_rom[ 5052]='h00000b5f;
    rd_cycle[ 5053] = 1'b1;  wr_cycle[ 5053] = 1'b0;  addr_rom[ 5053]='h00002f98;  wr_data_rom[ 5053]='h00000000;
    rd_cycle[ 5054] = 1'b0;  wr_cycle[ 5054] = 1'b1;  addr_rom[ 5054]='h00002854;  wr_data_rom[ 5054]='h00000106;
    rd_cycle[ 5055] = 1'b1;  wr_cycle[ 5055] = 1'b0;  addr_rom[ 5055]='h0000279c;  wr_data_rom[ 5055]='h00000000;
    rd_cycle[ 5056] = 1'b1;  wr_cycle[ 5056] = 1'b0;  addr_rom[ 5056]='h000033c4;  wr_data_rom[ 5056]='h00000000;
    rd_cycle[ 5057] = 1'b1;  wr_cycle[ 5057] = 1'b0;  addr_rom[ 5057]='h00002514;  wr_data_rom[ 5057]='h00000000;
    rd_cycle[ 5058] = 1'b0;  wr_cycle[ 5058] = 1'b1;  addr_rom[ 5058]='h00002cd0;  wr_data_rom[ 5058]='h0000040d;
    rd_cycle[ 5059] = 1'b1;  wr_cycle[ 5059] = 1'b0;  addr_rom[ 5059]='h0000104c;  wr_data_rom[ 5059]='h00000000;
    rd_cycle[ 5060] = 1'b0;  wr_cycle[ 5060] = 1'b1;  addr_rom[ 5060]='h000009c8;  wr_data_rom[ 5060]='h0000024f;
    rd_cycle[ 5061] = 1'b1;  wr_cycle[ 5061] = 1'b0;  addr_rom[ 5061]='h00000e0c;  wr_data_rom[ 5061]='h00000000;
    rd_cycle[ 5062] = 1'b1;  wr_cycle[ 5062] = 1'b0;  addr_rom[ 5062]='h00000dcc;  wr_data_rom[ 5062]='h00000000;
    rd_cycle[ 5063] = 1'b1;  wr_cycle[ 5063] = 1'b0;  addr_rom[ 5063]='h000035b8;  wr_data_rom[ 5063]='h00000000;
    rd_cycle[ 5064] = 1'b1;  wr_cycle[ 5064] = 1'b0;  addr_rom[ 5064]='h000028c8;  wr_data_rom[ 5064]='h00000000;
    rd_cycle[ 5065] = 1'b0;  wr_cycle[ 5065] = 1'b1;  addr_rom[ 5065]='h00000bc0;  wr_data_rom[ 5065]='h000011a4;
    rd_cycle[ 5066] = 1'b0;  wr_cycle[ 5066] = 1'b1;  addr_rom[ 5066]='h00001db0;  wr_data_rom[ 5066]='h000035a3;
    rd_cycle[ 5067] = 1'b0;  wr_cycle[ 5067] = 1'b1;  addr_rom[ 5067]='h00003ba0;  wr_data_rom[ 5067]='h000031e6;
    rd_cycle[ 5068] = 1'b0;  wr_cycle[ 5068] = 1'b1;  addr_rom[ 5068]='h000015c4;  wr_data_rom[ 5068]='h000020c0;
    rd_cycle[ 5069] = 1'b1;  wr_cycle[ 5069] = 1'b0;  addr_rom[ 5069]='h00000078;  wr_data_rom[ 5069]='h00000000;
    rd_cycle[ 5070] = 1'b0;  wr_cycle[ 5070] = 1'b1;  addr_rom[ 5070]='h00002d80;  wr_data_rom[ 5070]='h000018c6;
    rd_cycle[ 5071] = 1'b0;  wr_cycle[ 5071] = 1'b1;  addr_rom[ 5071]='h00002a98;  wr_data_rom[ 5071]='h00002836;
    rd_cycle[ 5072] = 1'b0;  wr_cycle[ 5072] = 1'b1;  addr_rom[ 5072]='h00001d2c;  wr_data_rom[ 5072]='h00001566;
    rd_cycle[ 5073] = 1'b1;  wr_cycle[ 5073] = 1'b0;  addr_rom[ 5073]='h00003c08;  wr_data_rom[ 5073]='h00000000;
    rd_cycle[ 5074] = 1'b1;  wr_cycle[ 5074] = 1'b0;  addr_rom[ 5074]='h0000194c;  wr_data_rom[ 5074]='h00000000;
    rd_cycle[ 5075] = 1'b1;  wr_cycle[ 5075] = 1'b0;  addr_rom[ 5075]='h00003f40;  wr_data_rom[ 5075]='h00000000;
    rd_cycle[ 5076] = 1'b1;  wr_cycle[ 5076] = 1'b0;  addr_rom[ 5076]='h00002f3c;  wr_data_rom[ 5076]='h00000000;
    rd_cycle[ 5077] = 1'b0;  wr_cycle[ 5077] = 1'b1;  addr_rom[ 5077]='h00003c68;  wr_data_rom[ 5077]='h00003c1c;
    rd_cycle[ 5078] = 1'b0;  wr_cycle[ 5078] = 1'b1;  addr_rom[ 5078]='h00002d44;  wr_data_rom[ 5078]='h000002b1;
    rd_cycle[ 5079] = 1'b0;  wr_cycle[ 5079] = 1'b1;  addr_rom[ 5079]='h00003ed0;  wr_data_rom[ 5079]='h00002005;
    rd_cycle[ 5080] = 1'b1;  wr_cycle[ 5080] = 1'b0;  addr_rom[ 5080]='h00001638;  wr_data_rom[ 5080]='h00000000;
    rd_cycle[ 5081] = 1'b0;  wr_cycle[ 5081] = 1'b1;  addr_rom[ 5081]='h00002af8;  wr_data_rom[ 5081]='h00000ed6;
    rd_cycle[ 5082] = 1'b1;  wr_cycle[ 5082] = 1'b0;  addr_rom[ 5082]='h000021d4;  wr_data_rom[ 5082]='h00000000;
    rd_cycle[ 5083] = 1'b1;  wr_cycle[ 5083] = 1'b0;  addr_rom[ 5083]='h0000340c;  wr_data_rom[ 5083]='h00000000;
    rd_cycle[ 5084] = 1'b0;  wr_cycle[ 5084] = 1'b1;  addr_rom[ 5084]='h00002af8;  wr_data_rom[ 5084]='h0000345f;
    rd_cycle[ 5085] = 1'b0;  wr_cycle[ 5085] = 1'b1;  addr_rom[ 5085]='h00003eec;  wr_data_rom[ 5085]='h00003491;
    rd_cycle[ 5086] = 1'b1;  wr_cycle[ 5086] = 1'b0;  addr_rom[ 5086]='h00000d44;  wr_data_rom[ 5086]='h00000000;
    rd_cycle[ 5087] = 1'b1;  wr_cycle[ 5087] = 1'b0;  addr_rom[ 5087]='h00000b20;  wr_data_rom[ 5087]='h00000000;
    rd_cycle[ 5088] = 1'b1;  wr_cycle[ 5088] = 1'b0;  addr_rom[ 5088]='h0000060c;  wr_data_rom[ 5088]='h00000000;
    rd_cycle[ 5089] = 1'b1;  wr_cycle[ 5089] = 1'b0;  addr_rom[ 5089]='h00002bfc;  wr_data_rom[ 5089]='h00000000;
    rd_cycle[ 5090] = 1'b1;  wr_cycle[ 5090] = 1'b0;  addr_rom[ 5090]='h00001c94;  wr_data_rom[ 5090]='h00000000;
    rd_cycle[ 5091] = 1'b1;  wr_cycle[ 5091] = 1'b0;  addr_rom[ 5091]='h000004c8;  wr_data_rom[ 5091]='h00000000;
    rd_cycle[ 5092] = 1'b0;  wr_cycle[ 5092] = 1'b1;  addr_rom[ 5092]='h00003814;  wr_data_rom[ 5092]='h00001893;
    rd_cycle[ 5093] = 1'b1;  wr_cycle[ 5093] = 1'b0;  addr_rom[ 5093]='h00002df0;  wr_data_rom[ 5093]='h00000000;
    rd_cycle[ 5094] = 1'b1;  wr_cycle[ 5094] = 1'b0;  addr_rom[ 5094]='h0000086c;  wr_data_rom[ 5094]='h00000000;
    rd_cycle[ 5095] = 1'b0;  wr_cycle[ 5095] = 1'b1;  addr_rom[ 5095]='h000017f4;  wr_data_rom[ 5095]='h00001f61;
    rd_cycle[ 5096] = 1'b1;  wr_cycle[ 5096] = 1'b0;  addr_rom[ 5096]='h00003d20;  wr_data_rom[ 5096]='h00000000;
    rd_cycle[ 5097] = 1'b1;  wr_cycle[ 5097] = 1'b0;  addr_rom[ 5097]='h00000fd4;  wr_data_rom[ 5097]='h00000000;
    rd_cycle[ 5098] = 1'b0;  wr_cycle[ 5098] = 1'b1;  addr_rom[ 5098]='h0000044c;  wr_data_rom[ 5098]='h00000c5b;
    rd_cycle[ 5099] = 1'b0;  wr_cycle[ 5099] = 1'b1;  addr_rom[ 5099]='h00002034;  wr_data_rom[ 5099]='h00003953;
    rd_cycle[ 5100] = 1'b0;  wr_cycle[ 5100] = 1'b1;  addr_rom[ 5100]='h00000804;  wr_data_rom[ 5100]='h000011b4;
    rd_cycle[ 5101] = 1'b0;  wr_cycle[ 5101] = 1'b1;  addr_rom[ 5101]='h00001a48;  wr_data_rom[ 5101]='h000027cf;
    rd_cycle[ 5102] = 1'b0;  wr_cycle[ 5102] = 1'b1;  addr_rom[ 5102]='h00003db4;  wr_data_rom[ 5102]='h00001ae6;
    rd_cycle[ 5103] = 1'b0;  wr_cycle[ 5103] = 1'b1;  addr_rom[ 5103]='h0000124c;  wr_data_rom[ 5103]='h00003ed4;
    rd_cycle[ 5104] = 1'b0;  wr_cycle[ 5104] = 1'b1;  addr_rom[ 5104]='h00003464;  wr_data_rom[ 5104]='h00001d15;
    rd_cycle[ 5105] = 1'b0;  wr_cycle[ 5105] = 1'b1;  addr_rom[ 5105]='h000004b4;  wr_data_rom[ 5105]='h00003b56;
    rd_cycle[ 5106] = 1'b1;  wr_cycle[ 5106] = 1'b0;  addr_rom[ 5106]='h00002aa8;  wr_data_rom[ 5106]='h00000000;
    rd_cycle[ 5107] = 1'b1;  wr_cycle[ 5107] = 1'b0;  addr_rom[ 5107]='h00001cf0;  wr_data_rom[ 5107]='h00000000;
    rd_cycle[ 5108] = 1'b1;  wr_cycle[ 5108] = 1'b0;  addr_rom[ 5108]='h000027a8;  wr_data_rom[ 5108]='h00000000;
    rd_cycle[ 5109] = 1'b0;  wr_cycle[ 5109] = 1'b1;  addr_rom[ 5109]='h000014d8;  wr_data_rom[ 5109]='h00000671;
    rd_cycle[ 5110] = 1'b0;  wr_cycle[ 5110] = 1'b1;  addr_rom[ 5110]='h00002718;  wr_data_rom[ 5110]='h00003ecd;
    rd_cycle[ 5111] = 1'b1;  wr_cycle[ 5111] = 1'b0;  addr_rom[ 5111]='h0000140c;  wr_data_rom[ 5111]='h00000000;
    rd_cycle[ 5112] = 1'b0;  wr_cycle[ 5112] = 1'b1;  addr_rom[ 5112]='h00000c0c;  wr_data_rom[ 5112]='h000010c6;
    rd_cycle[ 5113] = 1'b1;  wr_cycle[ 5113] = 1'b0;  addr_rom[ 5113]='h00003a64;  wr_data_rom[ 5113]='h00000000;
    rd_cycle[ 5114] = 1'b1;  wr_cycle[ 5114] = 1'b0;  addr_rom[ 5114]='h000002c4;  wr_data_rom[ 5114]='h00000000;
    rd_cycle[ 5115] = 1'b1;  wr_cycle[ 5115] = 1'b0;  addr_rom[ 5115]='h00001e68;  wr_data_rom[ 5115]='h00000000;
    rd_cycle[ 5116] = 1'b1;  wr_cycle[ 5116] = 1'b0;  addr_rom[ 5116]='h000014f0;  wr_data_rom[ 5116]='h00000000;
    rd_cycle[ 5117] = 1'b0;  wr_cycle[ 5117] = 1'b1;  addr_rom[ 5117]='h00000abc;  wr_data_rom[ 5117]='h0000207f;
    rd_cycle[ 5118] = 1'b1;  wr_cycle[ 5118] = 1'b0;  addr_rom[ 5118]='h00000428;  wr_data_rom[ 5118]='h00000000;
    rd_cycle[ 5119] = 1'b0;  wr_cycle[ 5119] = 1'b1;  addr_rom[ 5119]='h00002218;  wr_data_rom[ 5119]='h00001b34;
    rd_cycle[ 5120] = 1'b1;  wr_cycle[ 5120] = 1'b0;  addr_rom[ 5120]='h000000ec;  wr_data_rom[ 5120]='h00000000;
    rd_cycle[ 5121] = 1'b1;  wr_cycle[ 5121] = 1'b0;  addr_rom[ 5121]='h00001b30;  wr_data_rom[ 5121]='h00000000;
    rd_cycle[ 5122] = 1'b0;  wr_cycle[ 5122] = 1'b1;  addr_rom[ 5122]='h00003468;  wr_data_rom[ 5122]='h00003ea7;
    rd_cycle[ 5123] = 1'b0;  wr_cycle[ 5123] = 1'b1;  addr_rom[ 5123]='h00002e14;  wr_data_rom[ 5123]='h0000046b;
    rd_cycle[ 5124] = 1'b0;  wr_cycle[ 5124] = 1'b1;  addr_rom[ 5124]='h00002070;  wr_data_rom[ 5124]='h00001857;
    rd_cycle[ 5125] = 1'b1;  wr_cycle[ 5125] = 1'b0;  addr_rom[ 5125]='h00003914;  wr_data_rom[ 5125]='h00000000;
    rd_cycle[ 5126] = 1'b0;  wr_cycle[ 5126] = 1'b1;  addr_rom[ 5126]='h00003aac;  wr_data_rom[ 5126]='h000037c0;
    rd_cycle[ 5127] = 1'b1;  wr_cycle[ 5127] = 1'b0;  addr_rom[ 5127]='h000034f4;  wr_data_rom[ 5127]='h00000000;
    rd_cycle[ 5128] = 1'b1;  wr_cycle[ 5128] = 1'b0;  addr_rom[ 5128]='h000002ec;  wr_data_rom[ 5128]='h00000000;
    rd_cycle[ 5129] = 1'b0;  wr_cycle[ 5129] = 1'b1;  addr_rom[ 5129]='h0000114c;  wr_data_rom[ 5129]='h00002c7e;
    rd_cycle[ 5130] = 1'b1;  wr_cycle[ 5130] = 1'b0;  addr_rom[ 5130]='h000011b0;  wr_data_rom[ 5130]='h00000000;
    rd_cycle[ 5131] = 1'b0;  wr_cycle[ 5131] = 1'b1;  addr_rom[ 5131]='h00000050;  wr_data_rom[ 5131]='h0000346c;
    rd_cycle[ 5132] = 1'b0;  wr_cycle[ 5132] = 1'b1;  addr_rom[ 5132]='h00000f4c;  wr_data_rom[ 5132]='h00003df5;
    rd_cycle[ 5133] = 1'b1;  wr_cycle[ 5133] = 1'b0;  addr_rom[ 5133]='h00003a10;  wr_data_rom[ 5133]='h00000000;
    rd_cycle[ 5134] = 1'b1;  wr_cycle[ 5134] = 1'b0;  addr_rom[ 5134]='h00003b98;  wr_data_rom[ 5134]='h00000000;
    rd_cycle[ 5135] = 1'b0;  wr_cycle[ 5135] = 1'b1;  addr_rom[ 5135]='h00001574;  wr_data_rom[ 5135]='h00001fa6;
    rd_cycle[ 5136] = 1'b0;  wr_cycle[ 5136] = 1'b1;  addr_rom[ 5136]='h0000143c;  wr_data_rom[ 5136]='h00000230;
    rd_cycle[ 5137] = 1'b0;  wr_cycle[ 5137] = 1'b1;  addr_rom[ 5137]='h00001fec;  wr_data_rom[ 5137]='h0000315e;
    rd_cycle[ 5138] = 1'b1;  wr_cycle[ 5138] = 1'b0;  addr_rom[ 5138]='h000004bc;  wr_data_rom[ 5138]='h00000000;
    rd_cycle[ 5139] = 1'b0;  wr_cycle[ 5139] = 1'b1;  addr_rom[ 5139]='h00002898;  wr_data_rom[ 5139]='h00001a12;
    rd_cycle[ 5140] = 1'b0;  wr_cycle[ 5140] = 1'b1;  addr_rom[ 5140]='h00000f00;  wr_data_rom[ 5140]='h000005fc;
    rd_cycle[ 5141] = 1'b0;  wr_cycle[ 5141] = 1'b1;  addr_rom[ 5141]='h000023dc;  wr_data_rom[ 5141]='h00000229;
    rd_cycle[ 5142] = 1'b0;  wr_cycle[ 5142] = 1'b1;  addr_rom[ 5142]='h000024ec;  wr_data_rom[ 5142]='h0000017f;
    rd_cycle[ 5143] = 1'b1;  wr_cycle[ 5143] = 1'b0;  addr_rom[ 5143]='h0000112c;  wr_data_rom[ 5143]='h00000000;
    rd_cycle[ 5144] = 1'b1;  wr_cycle[ 5144] = 1'b0;  addr_rom[ 5144]='h000006a0;  wr_data_rom[ 5144]='h00000000;
    rd_cycle[ 5145] = 1'b1;  wr_cycle[ 5145] = 1'b0;  addr_rom[ 5145]='h00001648;  wr_data_rom[ 5145]='h00000000;
    rd_cycle[ 5146] = 1'b1;  wr_cycle[ 5146] = 1'b0;  addr_rom[ 5146]='h000019f4;  wr_data_rom[ 5146]='h00000000;
    rd_cycle[ 5147] = 1'b1;  wr_cycle[ 5147] = 1'b0;  addr_rom[ 5147]='h00003970;  wr_data_rom[ 5147]='h00000000;
    rd_cycle[ 5148] = 1'b1;  wr_cycle[ 5148] = 1'b0;  addr_rom[ 5148]='h00003478;  wr_data_rom[ 5148]='h00000000;
    rd_cycle[ 5149] = 1'b0;  wr_cycle[ 5149] = 1'b1;  addr_rom[ 5149]='h00001b90;  wr_data_rom[ 5149]='h00000cd1;
    rd_cycle[ 5150] = 1'b0;  wr_cycle[ 5150] = 1'b1;  addr_rom[ 5150]='h00000b50;  wr_data_rom[ 5150]='h000027b9;
    rd_cycle[ 5151] = 1'b1;  wr_cycle[ 5151] = 1'b0;  addr_rom[ 5151]='h00003860;  wr_data_rom[ 5151]='h00000000;
    rd_cycle[ 5152] = 1'b0;  wr_cycle[ 5152] = 1'b1;  addr_rom[ 5152]='h00000cd4;  wr_data_rom[ 5152]='h000036ae;
    rd_cycle[ 5153] = 1'b0;  wr_cycle[ 5153] = 1'b1;  addr_rom[ 5153]='h00001e94;  wr_data_rom[ 5153]='h00000851;
    rd_cycle[ 5154] = 1'b0;  wr_cycle[ 5154] = 1'b1;  addr_rom[ 5154]='h00000db4;  wr_data_rom[ 5154]='h00000d4e;
    rd_cycle[ 5155] = 1'b0;  wr_cycle[ 5155] = 1'b1;  addr_rom[ 5155]='h0000318c;  wr_data_rom[ 5155]='h00001865;
    rd_cycle[ 5156] = 1'b0;  wr_cycle[ 5156] = 1'b1;  addr_rom[ 5156]='h000004c8;  wr_data_rom[ 5156]='h00001113;
    rd_cycle[ 5157] = 1'b0;  wr_cycle[ 5157] = 1'b1;  addr_rom[ 5157]='h00002ab0;  wr_data_rom[ 5157]='h00000432;
    rd_cycle[ 5158] = 1'b0;  wr_cycle[ 5158] = 1'b1;  addr_rom[ 5158]='h00001288;  wr_data_rom[ 5158]='h00001e3e;
    rd_cycle[ 5159] = 1'b0;  wr_cycle[ 5159] = 1'b1;  addr_rom[ 5159]='h00000b40;  wr_data_rom[ 5159]='h0000030a;
    rd_cycle[ 5160] = 1'b0;  wr_cycle[ 5160] = 1'b1;  addr_rom[ 5160]='h00000cb0;  wr_data_rom[ 5160]='h000025ea;
    rd_cycle[ 5161] = 1'b1;  wr_cycle[ 5161] = 1'b0;  addr_rom[ 5161]='h00003e5c;  wr_data_rom[ 5161]='h00000000;
    rd_cycle[ 5162] = 1'b0;  wr_cycle[ 5162] = 1'b1;  addr_rom[ 5162]='h00000b4c;  wr_data_rom[ 5162]='h00001c5a;
    rd_cycle[ 5163] = 1'b1;  wr_cycle[ 5163] = 1'b0;  addr_rom[ 5163]='h00002adc;  wr_data_rom[ 5163]='h00000000;
    rd_cycle[ 5164] = 1'b0;  wr_cycle[ 5164] = 1'b1;  addr_rom[ 5164]='h00001990;  wr_data_rom[ 5164]='h00002ee6;
    rd_cycle[ 5165] = 1'b0;  wr_cycle[ 5165] = 1'b1;  addr_rom[ 5165]='h00001f1c;  wr_data_rom[ 5165]='h00003e86;
    rd_cycle[ 5166] = 1'b1;  wr_cycle[ 5166] = 1'b0;  addr_rom[ 5166]='h00003174;  wr_data_rom[ 5166]='h00000000;
    rd_cycle[ 5167] = 1'b0;  wr_cycle[ 5167] = 1'b1;  addr_rom[ 5167]='h00002e94;  wr_data_rom[ 5167]='h00000de8;
    rd_cycle[ 5168] = 1'b0;  wr_cycle[ 5168] = 1'b1;  addr_rom[ 5168]='h00000ee8;  wr_data_rom[ 5168]='h000028e8;
    rd_cycle[ 5169] = 1'b0;  wr_cycle[ 5169] = 1'b1;  addr_rom[ 5169]='h00002a28;  wr_data_rom[ 5169]='h00002597;
    rd_cycle[ 5170] = 1'b0;  wr_cycle[ 5170] = 1'b1;  addr_rom[ 5170]='h00002cb0;  wr_data_rom[ 5170]='h00002fdf;
    rd_cycle[ 5171] = 1'b1;  wr_cycle[ 5171] = 1'b0;  addr_rom[ 5171]='h00003ad4;  wr_data_rom[ 5171]='h00000000;
    rd_cycle[ 5172] = 1'b0;  wr_cycle[ 5172] = 1'b1;  addr_rom[ 5172]='h00002d94;  wr_data_rom[ 5172]='h00003c88;
    rd_cycle[ 5173] = 1'b0;  wr_cycle[ 5173] = 1'b1;  addr_rom[ 5173]='h000014ac;  wr_data_rom[ 5173]='h00000d22;
    rd_cycle[ 5174] = 1'b0;  wr_cycle[ 5174] = 1'b1;  addr_rom[ 5174]='h00001828;  wr_data_rom[ 5174]='h00003b41;
    rd_cycle[ 5175] = 1'b1;  wr_cycle[ 5175] = 1'b0;  addr_rom[ 5175]='h000020dc;  wr_data_rom[ 5175]='h00000000;
    rd_cycle[ 5176] = 1'b0;  wr_cycle[ 5176] = 1'b1;  addr_rom[ 5176]='h000009a8;  wr_data_rom[ 5176]='h00000c26;
    rd_cycle[ 5177] = 1'b0;  wr_cycle[ 5177] = 1'b1;  addr_rom[ 5177]='h00000358;  wr_data_rom[ 5177]='h000007fd;
    rd_cycle[ 5178] = 1'b0;  wr_cycle[ 5178] = 1'b1;  addr_rom[ 5178]='h00002c14;  wr_data_rom[ 5178]='h00002590;
    rd_cycle[ 5179] = 1'b0;  wr_cycle[ 5179] = 1'b1;  addr_rom[ 5179]='h000013f4;  wr_data_rom[ 5179]='h000000a8;
    rd_cycle[ 5180] = 1'b0;  wr_cycle[ 5180] = 1'b1;  addr_rom[ 5180]='h000024a8;  wr_data_rom[ 5180]='h00002c75;
    rd_cycle[ 5181] = 1'b0;  wr_cycle[ 5181] = 1'b1;  addr_rom[ 5181]='h00000538;  wr_data_rom[ 5181]='h00002f2b;
    rd_cycle[ 5182] = 1'b1;  wr_cycle[ 5182] = 1'b0;  addr_rom[ 5182]='h00001118;  wr_data_rom[ 5182]='h00000000;
    rd_cycle[ 5183] = 1'b0;  wr_cycle[ 5183] = 1'b1;  addr_rom[ 5183]='h000004b8;  wr_data_rom[ 5183]='h00001da9;
    rd_cycle[ 5184] = 1'b0;  wr_cycle[ 5184] = 1'b1;  addr_rom[ 5184]='h00003608;  wr_data_rom[ 5184]='h00001fb5;
    rd_cycle[ 5185] = 1'b1;  wr_cycle[ 5185] = 1'b0;  addr_rom[ 5185]='h00003304;  wr_data_rom[ 5185]='h00000000;
    rd_cycle[ 5186] = 1'b0;  wr_cycle[ 5186] = 1'b1;  addr_rom[ 5186]='h00003bb4;  wr_data_rom[ 5186]='h00003c0e;
    rd_cycle[ 5187] = 1'b0;  wr_cycle[ 5187] = 1'b1;  addr_rom[ 5187]='h0000179c;  wr_data_rom[ 5187]='h000020ce;
    rd_cycle[ 5188] = 1'b0;  wr_cycle[ 5188] = 1'b1;  addr_rom[ 5188]='h00003344;  wr_data_rom[ 5188]='h00002caf;
    rd_cycle[ 5189] = 1'b0;  wr_cycle[ 5189] = 1'b1;  addr_rom[ 5189]='h000033e4;  wr_data_rom[ 5189]='h00000aa2;
    rd_cycle[ 5190] = 1'b0;  wr_cycle[ 5190] = 1'b1;  addr_rom[ 5190]='h00001258;  wr_data_rom[ 5190]='h0000312d;
    rd_cycle[ 5191] = 1'b0;  wr_cycle[ 5191] = 1'b1;  addr_rom[ 5191]='h000034f0;  wr_data_rom[ 5191]='h000001ed;
    rd_cycle[ 5192] = 1'b1;  wr_cycle[ 5192] = 1'b0;  addr_rom[ 5192]='h0000123c;  wr_data_rom[ 5192]='h00000000;
    rd_cycle[ 5193] = 1'b0;  wr_cycle[ 5193] = 1'b1;  addr_rom[ 5193]='h00001250;  wr_data_rom[ 5193]='h000018f2;
    rd_cycle[ 5194] = 1'b1;  wr_cycle[ 5194] = 1'b0;  addr_rom[ 5194]='h0000241c;  wr_data_rom[ 5194]='h00000000;
    rd_cycle[ 5195] = 1'b1;  wr_cycle[ 5195] = 1'b0;  addr_rom[ 5195]='h00002abc;  wr_data_rom[ 5195]='h00000000;
    rd_cycle[ 5196] = 1'b0;  wr_cycle[ 5196] = 1'b1;  addr_rom[ 5196]='h000000a8;  wr_data_rom[ 5196]='h000009a1;
    rd_cycle[ 5197] = 1'b0;  wr_cycle[ 5197] = 1'b1;  addr_rom[ 5197]='h000035ac;  wr_data_rom[ 5197]='h00003cf3;
    rd_cycle[ 5198] = 1'b1;  wr_cycle[ 5198] = 1'b0;  addr_rom[ 5198]='h0000325c;  wr_data_rom[ 5198]='h00000000;
    rd_cycle[ 5199] = 1'b1;  wr_cycle[ 5199] = 1'b0;  addr_rom[ 5199]='h0000237c;  wr_data_rom[ 5199]='h00000000;
    rd_cycle[ 5200] = 1'b1;  wr_cycle[ 5200] = 1'b0;  addr_rom[ 5200]='h000039a8;  wr_data_rom[ 5200]='h00000000;
    rd_cycle[ 5201] = 1'b0;  wr_cycle[ 5201] = 1'b1;  addr_rom[ 5201]='h00000220;  wr_data_rom[ 5201]='h00001cfb;
    rd_cycle[ 5202] = 1'b0;  wr_cycle[ 5202] = 1'b1;  addr_rom[ 5202]='h0000394c;  wr_data_rom[ 5202]='h000005fe;
    rd_cycle[ 5203] = 1'b1;  wr_cycle[ 5203] = 1'b0;  addr_rom[ 5203]='h00000954;  wr_data_rom[ 5203]='h00000000;
    rd_cycle[ 5204] = 1'b0;  wr_cycle[ 5204] = 1'b1;  addr_rom[ 5204]='h0000158c;  wr_data_rom[ 5204]='h000004c8;
    rd_cycle[ 5205] = 1'b0;  wr_cycle[ 5205] = 1'b1;  addr_rom[ 5205]='h000015e0;  wr_data_rom[ 5205]='h0000073d;
    rd_cycle[ 5206] = 1'b1;  wr_cycle[ 5206] = 1'b0;  addr_rom[ 5206]='h00001238;  wr_data_rom[ 5206]='h00000000;
    rd_cycle[ 5207] = 1'b0;  wr_cycle[ 5207] = 1'b1;  addr_rom[ 5207]='h000026d0;  wr_data_rom[ 5207]='h000037e9;
    rd_cycle[ 5208] = 1'b0;  wr_cycle[ 5208] = 1'b1;  addr_rom[ 5208]='h00001b88;  wr_data_rom[ 5208]='h00002f3f;
    rd_cycle[ 5209] = 1'b0;  wr_cycle[ 5209] = 1'b1;  addr_rom[ 5209]='h00002120;  wr_data_rom[ 5209]='h00000965;
    rd_cycle[ 5210] = 1'b0;  wr_cycle[ 5210] = 1'b1;  addr_rom[ 5210]='h00001bd8;  wr_data_rom[ 5210]='h000013ef;
    rd_cycle[ 5211] = 1'b1;  wr_cycle[ 5211] = 1'b0;  addr_rom[ 5211]='h000003b8;  wr_data_rom[ 5211]='h00000000;
    rd_cycle[ 5212] = 1'b0;  wr_cycle[ 5212] = 1'b1;  addr_rom[ 5212]='h000011b0;  wr_data_rom[ 5212]='h00003d8d;
    rd_cycle[ 5213] = 1'b0;  wr_cycle[ 5213] = 1'b1;  addr_rom[ 5213]='h00003530;  wr_data_rom[ 5213]='h00003800;
    rd_cycle[ 5214] = 1'b0;  wr_cycle[ 5214] = 1'b1;  addr_rom[ 5214]='h00003b74;  wr_data_rom[ 5214]='h00001cfa;
    rd_cycle[ 5215] = 1'b0;  wr_cycle[ 5215] = 1'b1;  addr_rom[ 5215]='h00000930;  wr_data_rom[ 5215]='h0000307a;
    rd_cycle[ 5216] = 1'b0;  wr_cycle[ 5216] = 1'b1;  addr_rom[ 5216]='h00003bd0;  wr_data_rom[ 5216]='h000024aa;
    rd_cycle[ 5217] = 1'b1;  wr_cycle[ 5217] = 1'b0;  addr_rom[ 5217]='h00001f94;  wr_data_rom[ 5217]='h00000000;
    rd_cycle[ 5218] = 1'b1;  wr_cycle[ 5218] = 1'b0;  addr_rom[ 5218]='h00003980;  wr_data_rom[ 5218]='h00000000;
    rd_cycle[ 5219] = 1'b0;  wr_cycle[ 5219] = 1'b1;  addr_rom[ 5219]='h00000ae8;  wr_data_rom[ 5219]='h0000353f;
    rd_cycle[ 5220] = 1'b0;  wr_cycle[ 5220] = 1'b1;  addr_rom[ 5220]='h00001680;  wr_data_rom[ 5220]='h00000c3c;
    rd_cycle[ 5221] = 1'b1;  wr_cycle[ 5221] = 1'b0;  addr_rom[ 5221]='h00003080;  wr_data_rom[ 5221]='h00000000;
    rd_cycle[ 5222] = 1'b1;  wr_cycle[ 5222] = 1'b0;  addr_rom[ 5222]='h0000317c;  wr_data_rom[ 5222]='h00000000;
    rd_cycle[ 5223] = 1'b0;  wr_cycle[ 5223] = 1'b1;  addr_rom[ 5223]='h00002f28;  wr_data_rom[ 5223]='h00003662;
    rd_cycle[ 5224] = 1'b1;  wr_cycle[ 5224] = 1'b0;  addr_rom[ 5224]='h0000039c;  wr_data_rom[ 5224]='h00000000;
    rd_cycle[ 5225] = 1'b0;  wr_cycle[ 5225] = 1'b1;  addr_rom[ 5225]='h00001e90;  wr_data_rom[ 5225]='h00001785;
    rd_cycle[ 5226] = 1'b0;  wr_cycle[ 5226] = 1'b1;  addr_rom[ 5226]='h0000146c;  wr_data_rom[ 5226]='h00000a83;
    rd_cycle[ 5227] = 1'b1;  wr_cycle[ 5227] = 1'b0;  addr_rom[ 5227]='h00002ee0;  wr_data_rom[ 5227]='h00000000;
    rd_cycle[ 5228] = 1'b0;  wr_cycle[ 5228] = 1'b1;  addr_rom[ 5228]='h00002d58;  wr_data_rom[ 5228]='h00003d18;
    rd_cycle[ 5229] = 1'b1;  wr_cycle[ 5229] = 1'b0;  addr_rom[ 5229]='h00003e9c;  wr_data_rom[ 5229]='h00000000;
    rd_cycle[ 5230] = 1'b1;  wr_cycle[ 5230] = 1'b0;  addr_rom[ 5230]='h00002bd0;  wr_data_rom[ 5230]='h00000000;
    rd_cycle[ 5231] = 1'b0;  wr_cycle[ 5231] = 1'b1;  addr_rom[ 5231]='h00002290;  wr_data_rom[ 5231]='h00002262;
    rd_cycle[ 5232] = 1'b1;  wr_cycle[ 5232] = 1'b0;  addr_rom[ 5232]='h00003df0;  wr_data_rom[ 5232]='h00000000;
    rd_cycle[ 5233] = 1'b1;  wr_cycle[ 5233] = 1'b0;  addr_rom[ 5233]='h000006f8;  wr_data_rom[ 5233]='h00000000;
    rd_cycle[ 5234] = 1'b1;  wr_cycle[ 5234] = 1'b0;  addr_rom[ 5234]='h000005cc;  wr_data_rom[ 5234]='h00000000;
    rd_cycle[ 5235] = 1'b0;  wr_cycle[ 5235] = 1'b1;  addr_rom[ 5235]='h000005c4;  wr_data_rom[ 5235]='h00000d14;
    rd_cycle[ 5236] = 1'b1;  wr_cycle[ 5236] = 1'b0;  addr_rom[ 5236]='h000010f8;  wr_data_rom[ 5236]='h00000000;
    rd_cycle[ 5237] = 1'b0;  wr_cycle[ 5237] = 1'b1;  addr_rom[ 5237]='h0000102c;  wr_data_rom[ 5237]='h00003fc6;
    rd_cycle[ 5238] = 1'b0;  wr_cycle[ 5238] = 1'b1;  addr_rom[ 5238]='h00001a70;  wr_data_rom[ 5238]='h00001dae;
    rd_cycle[ 5239] = 1'b0;  wr_cycle[ 5239] = 1'b1;  addr_rom[ 5239]='h00003a70;  wr_data_rom[ 5239]='h0000031a;
    rd_cycle[ 5240] = 1'b1;  wr_cycle[ 5240] = 1'b0;  addr_rom[ 5240]='h00002ea8;  wr_data_rom[ 5240]='h00000000;
    rd_cycle[ 5241] = 1'b0;  wr_cycle[ 5241] = 1'b1;  addr_rom[ 5241]='h000037ac;  wr_data_rom[ 5241]='h00001e9e;
    rd_cycle[ 5242] = 1'b1;  wr_cycle[ 5242] = 1'b0;  addr_rom[ 5242]='h00003924;  wr_data_rom[ 5242]='h00000000;
    rd_cycle[ 5243] = 1'b1;  wr_cycle[ 5243] = 1'b0;  addr_rom[ 5243]='h00003f7c;  wr_data_rom[ 5243]='h00000000;
    rd_cycle[ 5244] = 1'b0;  wr_cycle[ 5244] = 1'b1;  addr_rom[ 5244]='h000016bc;  wr_data_rom[ 5244]='h00003665;
    rd_cycle[ 5245] = 1'b1;  wr_cycle[ 5245] = 1'b0;  addr_rom[ 5245]='h00002f98;  wr_data_rom[ 5245]='h00000000;
    rd_cycle[ 5246] = 1'b1;  wr_cycle[ 5246] = 1'b0;  addr_rom[ 5246]='h00000c9c;  wr_data_rom[ 5246]='h00000000;
    rd_cycle[ 5247] = 1'b0;  wr_cycle[ 5247] = 1'b1;  addr_rom[ 5247]='h00003d2c;  wr_data_rom[ 5247]='h000018ae;
    rd_cycle[ 5248] = 1'b1;  wr_cycle[ 5248] = 1'b0;  addr_rom[ 5248]='h00000738;  wr_data_rom[ 5248]='h00000000;
    rd_cycle[ 5249] = 1'b1;  wr_cycle[ 5249] = 1'b0;  addr_rom[ 5249]='h00001800;  wr_data_rom[ 5249]='h00000000;
    rd_cycle[ 5250] = 1'b0;  wr_cycle[ 5250] = 1'b1;  addr_rom[ 5250]='h000031fc;  wr_data_rom[ 5250]='h000035a4;
    rd_cycle[ 5251] = 1'b0;  wr_cycle[ 5251] = 1'b1;  addr_rom[ 5251]='h00000180;  wr_data_rom[ 5251]='h000021d7;
    rd_cycle[ 5252] = 1'b1;  wr_cycle[ 5252] = 1'b0;  addr_rom[ 5252]='h00000b64;  wr_data_rom[ 5252]='h00000000;
    rd_cycle[ 5253] = 1'b1;  wr_cycle[ 5253] = 1'b0;  addr_rom[ 5253]='h0000259c;  wr_data_rom[ 5253]='h00000000;
    rd_cycle[ 5254] = 1'b1;  wr_cycle[ 5254] = 1'b0;  addr_rom[ 5254]='h00003238;  wr_data_rom[ 5254]='h00000000;
    rd_cycle[ 5255] = 1'b0;  wr_cycle[ 5255] = 1'b1;  addr_rom[ 5255]='h00000ca8;  wr_data_rom[ 5255]='h00000d77;
    rd_cycle[ 5256] = 1'b0;  wr_cycle[ 5256] = 1'b1;  addr_rom[ 5256]='h000022e4;  wr_data_rom[ 5256]='h00003d35;
    rd_cycle[ 5257] = 1'b0;  wr_cycle[ 5257] = 1'b1;  addr_rom[ 5257]='h00002ff8;  wr_data_rom[ 5257]='h0000072f;
    rd_cycle[ 5258] = 1'b0;  wr_cycle[ 5258] = 1'b1;  addr_rom[ 5258]='h000001a8;  wr_data_rom[ 5258]='h000035a7;
    rd_cycle[ 5259] = 1'b1;  wr_cycle[ 5259] = 1'b0;  addr_rom[ 5259]='h00001eac;  wr_data_rom[ 5259]='h00000000;
    rd_cycle[ 5260] = 1'b1;  wr_cycle[ 5260] = 1'b0;  addr_rom[ 5260]='h00003908;  wr_data_rom[ 5260]='h00000000;
    rd_cycle[ 5261] = 1'b1;  wr_cycle[ 5261] = 1'b0;  addr_rom[ 5261]='h00002190;  wr_data_rom[ 5261]='h00000000;
    rd_cycle[ 5262] = 1'b0;  wr_cycle[ 5262] = 1'b1;  addr_rom[ 5262]='h00002df0;  wr_data_rom[ 5262]='h000025cf;
    rd_cycle[ 5263] = 1'b0;  wr_cycle[ 5263] = 1'b1;  addr_rom[ 5263]='h00000bec;  wr_data_rom[ 5263]='h00002853;
    rd_cycle[ 5264] = 1'b1;  wr_cycle[ 5264] = 1'b0;  addr_rom[ 5264]='h000025b8;  wr_data_rom[ 5264]='h00000000;
    rd_cycle[ 5265] = 1'b0;  wr_cycle[ 5265] = 1'b1;  addr_rom[ 5265]='h000000cc;  wr_data_rom[ 5265]='h0000102f;
    rd_cycle[ 5266] = 1'b1;  wr_cycle[ 5266] = 1'b0;  addr_rom[ 5266]='h000014e8;  wr_data_rom[ 5266]='h00000000;
    rd_cycle[ 5267] = 1'b0;  wr_cycle[ 5267] = 1'b1;  addr_rom[ 5267]='h000033c0;  wr_data_rom[ 5267]='h00000cb1;
    rd_cycle[ 5268] = 1'b0;  wr_cycle[ 5268] = 1'b1;  addr_rom[ 5268]='h0000387c;  wr_data_rom[ 5268]='h00000a47;
    rd_cycle[ 5269] = 1'b1;  wr_cycle[ 5269] = 1'b0;  addr_rom[ 5269]='h00002968;  wr_data_rom[ 5269]='h00000000;
    rd_cycle[ 5270] = 1'b1;  wr_cycle[ 5270] = 1'b0;  addr_rom[ 5270]='h000003a0;  wr_data_rom[ 5270]='h00000000;
    rd_cycle[ 5271] = 1'b1;  wr_cycle[ 5271] = 1'b0;  addr_rom[ 5271]='h00002f28;  wr_data_rom[ 5271]='h00000000;
    rd_cycle[ 5272] = 1'b0;  wr_cycle[ 5272] = 1'b1;  addr_rom[ 5272]='h00001a74;  wr_data_rom[ 5272]='h000013f8;
    rd_cycle[ 5273] = 1'b1;  wr_cycle[ 5273] = 1'b0;  addr_rom[ 5273]='h000012f4;  wr_data_rom[ 5273]='h00000000;
    rd_cycle[ 5274] = 1'b0;  wr_cycle[ 5274] = 1'b1;  addr_rom[ 5274]='h00002b00;  wr_data_rom[ 5274]='h0000160c;
    rd_cycle[ 5275] = 1'b1;  wr_cycle[ 5275] = 1'b0;  addr_rom[ 5275]='h00001c2c;  wr_data_rom[ 5275]='h00000000;
    rd_cycle[ 5276] = 1'b1;  wr_cycle[ 5276] = 1'b0;  addr_rom[ 5276]='h00002dcc;  wr_data_rom[ 5276]='h00000000;
    rd_cycle[ 5277] = 1'b1;  wr_cycle[ 5277] = 1'b0;  addr_rom[ 5277]='h000030cc;  wr_data_rom[ 5277]='h00000000;
    rd_cycle[ 5278] = 1'b0;  wr_cycle[ 5278] = 1'b1;  addr_rom[ 5278]='h00002e28;  wr_data_rom[ 5278]='h00002346;
    rd_cycle[ 5279] = 1'b1;  wr_cycle[ 5279] = 1'b0;  addr_rom[ 5279]='h00000728;  wr_data_rom[ 5279]='h00000000;
    rd_cycle[ 5280] = 1'b0;  wr_cycle[ 5280] = 1'b1;  addr_rom[ 5280]='h00000c80;  wr_data_rom[ 5280]='h00003f64;
    rd_cycle[ 5281] = 1'b1;  wr_cycle[ 5281] = 1'b0;  addr_rom[ 5281]='h00001b1c;  wr_data_rom[ 5281]='h00000000;
    rd_cycle[ 5282] = 1'b1;  wr_cycle[ 5282] = 1'b0;  addr_rom[ 5282]='h000000c4;  wr_data_rom[ 5282]='h00000000;
    rd_cycle[ 5283] = 1'b0;  wr_cycle[ 5283] = 1'b1;  addr_rom[ 5283]='h00000aa0;  wr_data_rom[ 5283]='h00001d91;
    rd_cycle[ 5284] = 1'b0;  wr_cycle[ 5284] = 1'b1;  addr_rom[ 5284]='h000003e8;  wr_data_rom[ 5284]='h000008d4;
    rd_cycle[ 5285] = 1'b1;  wr_cycle[ 5285] = 1'b0;  addr_rom[ 5285]='h00001268;  wr_data_rom[ 5285]='h00000000;
    rd_cycle[ 5286] = 1'b1;  wr_cycle[ 5286] = 1'b0;  addr_rom[ 5286]='h00000c18;  wr_data_rom[ 5286]='h00000000;
    rd_cycle[ 5287] = 1'b0;  wr_cycle[ 5287] = 1'b1;  addr_rom[ 5287]='h00000a50;  wr_data_rom[ 5287]='h00002524;
    rd_cycle[ 5288] = 1'b1;  wr_cycle[ 5288] = 1'b0;  addr_rom[ 5288]='h00000f14;  wr_data_rom[ 5288]='h00000000;
    rd_cycle[ 5289] = 1'b0;  wr_cycle[ 5289] = 1'b1;  addr_rom[ 5289]='h00000c44;  wr_data_rom[ 5289]='h000033cb;
    rd_cycle[ 5290] = 1'b1;  wr_cycle[ 5290] = 1'b0;  addr_rom[ 5290]='h00000b28;  wr_data_rom[ 5290]='h00000000;
    rd_cycle[ 5291] = 1'b0;  wr_cycle[ 5291] = 1'b1;  addr_rom[ 5291]='h00000edc;  wr_data_rom[ 5291]='h0000256d;
    rd_cycle[ 5292] = 1'b0;  wr_cycle[ 5292] = 1'b1;  addr_rom[ 5292]='h00001658;  wr_data_rom[ 5292]='h000009f1;
    rd_cycle[ 5293] = 1'b1;  wr_cycle[ 5293] = 1'b0;  addr_rom[ 5293]='h00001408;  wr_data_rom[ 5293]='h00000000;
    rd_cycle[ 5294] = 1'b0;  wr_cycle[ 5294] = 1'b1;  addr_rom[ 5294]='h00003f68;  wr_data_rom[ 5294]='h00003580;
    rd_cycle[ 5295] = 1'b1;  wr_cycle[ 5295] = 1'b0;  addr_rom[ 5295]='h00002e74;  wr_data_rom[ 5295]='h00000000;
    rd_cycle[ 5296] = 1'b0;  wr_cycle[ 5296] = 1'b1;  addr_rom[ 5296]='h00003024;  wr_data_rom[ 5296]='h00002ff4;
    rd_cycle[ 5297] = 1'b0;  wr_cycle[ 5297] = 1'b1;  addr_rom[ 5297]='h00003df0;  wr_data_rom[ 5297]='h000010da;
    rd_cycle[ 5298] = 1'b1;  wr_cycle[ 5298] = 1'b0;  addr_rom[ 5298]='h000000c4;  wr_data_rom[ 5298]='h00000000;
    rd_cycle[ 5299] = 1'b0;  wr_cycle[ 5299] = 1'b1;  addr_rom[ 5299]='h0000343c;  wr_data_rom[ 5299]='h00002832;
    rd_cycle[ 5300] = 1'b0;  wr_cycle[ 5300] = 1'b1;  addr_rom[ 5300]='h00002dfc;  wr_data_rom[ 5300]='h000010d6;
    rd_cycle[ 5301] = 1'b1;  wr_cycle[ 5301] = 1'b0;  addr_rom[ 5301]='h00001c04;  wr_data_rom[ 5301]='h00000000;
    rd_cycle[ 5302] = 1'b0;  wr_cycle[ 5302] = 1'b1;  addr_rom[ 5302]='h00000cc0;  wr_data_rom[ 5302]='h0000209b;
    rd_cycle[ 5303] = 1'b1;  wr_cycle[ 5303] = 1'b0;  addr_rom[ 5303]='h000037fc;  wr_data_rom[ 5303]='h00000000;
    rd_cycle[ 5304] = 1'b0;  wr_cycle[ 5304] = 1'b1;  addr_rom[ 5304]='h00003b20;  wr_data_rom[ 5304]='h00002cd8;
    rd_cycle[ 5305] = 1'b1;  wr_cycle[ 5305] = 1'b0;  addr_rom[ 5305]='h00003c3c;  wr_data_rom[ 5305]='h00000000;
    rd_cycle[ 5306] = 1'b0;  wr_cycle[ 5306] = 1'b1;  addr_rom[ 5306]='h00002de4;  wr_data_rom[ 5306]='h0000276d;
    rd_cycle[ 5307] = 1'b0;  wr_cycle[ 5307] = 1'b1;  addr_rom[ 5307]='h00002160;  wr_data_rom[ 5307]='h000021d5;
    rd_cycle[ 5308] = 1'b0;  wr_cycle[ 5308] = 1'b1;  addr_rom[ 5308]='h0000091c;  wr_data_rom[ 5308]='h00001a33;
    rd_cycle[ 5309] = 1'b0;  wr_cycle[ 5309] = 1'b1;  addr_rom[ 5309]='h00001400;  wr_data_rom[ 5309]='h000038ea;
    rd_cycle[ 5310] = 1'b0;  wr_cycle[ 5310] = 1'b1;  addr_rom[ 5310]='h00002638;  wr_data_rom[ 5310]='h00003b4c;
    rd_cycle[ 5311] = 1'b0;  wr_cycle[ 5311] = 1'b1;  addr_rom[ 5311]='h00002f40;  wr_data_rom[ 5311]='h00001b73;
    rd_cycle[ 5312] = 1'b0;  wr_cycle[ 5312] = 1'b1;  addr_rom[ 5312]='h00003990;  wr_data_rom[ 5312]='h0000185f;
    rd_cycle[ 5313] = 1'b1;  wr_cycle[ 5313] = 1'b0;  addr_rom[ 5313]='h000014f4;  wr_data_rom[ 5313]='h00000000;
    rd_cycle[ 5314] = 1'b1;  wr_cycle[ 5314] = 1'b0;  addr_rom[ 5314]='h00002690;  wr_data_rom[ 5314]='h00000000;
    rd_cycle[ 5315] = 1'b1;  wr_cycle[ 5315] = 1'b0;  addr_rom[ 5315]='h00000cbc;  wr_data_rom[ 5315]='h00000000;
    rd_cycle[ 5316] = 1'b1;  wr_cycle[ 5316] = 1'b0;  addr_rom[ 5316]='h0000028c;  wr_data_rom[ 5316]='h00000000;
    rd_cycle[ 5317] = 1'b0;  wr_cycle[ 5317] = 1'b1;  addr_rom[ 5317]='h00002018;  wr_data_rom[ 5317]='h00001337;
    rd_cycle[ 5318] = 1'b0;  wr_cycle[ 5318] = 1'b1;  addr_rom[ 5318]='h00003b1c;  wr_data_rom[ 5318]='h00000d5f;
    rd_cycle[ 5319] = 1'b0;  wr_cycle[ 5319] = 1'b1;  addr_rom[ 5319]='h00001870;  wr_data_rom[ 5319]='h00000e62;
    rd_cycle[ 5320] = 1'b1;  wr_cycle[ 5320] = 1'b0;  addr_rom[ 5320]='h00001500;  wr_data_rom[ 5320]='h00000000;
    rd_cycle[ 5321] = 1'b0;  wr_cycle[ 5321] = 1'b1;  addr_rom[ 5321]='h00001cd8;  wr_data_rom[ 5321]='h000014f4;
    rd_cycle[ 5322] = 1'b0;  wr_cycle[ 5322] = 1'b1;  addr_rom[ 5322]='h0000336c;  wr_data_rom[ 5322]='h00003f0f;
    rd_cycle[ 5323] = 1'b0;  wr_cycle[ 5323] = 1'b1;  addr_rom[ 5323]='h0000309c;  wr_data_rom[ 5323]='h00003594;
    rd_cycle[ 5324] = 1'b1;  wr_cycle[ 5324] = 1'b0;  addr_rom[ 5324]='h000007e0;  wr_data_rom[ 5324]='h00000000;
    rd_cycle[ 5325] = 1'b1;  wr_cycle[ 5325] = 1'b0;  addr_rom[ 5325]='h000018ac;  wr_data_rom[ 5325]='h00000000;
    rd_cycle[ 5326] = 1'b0;  wr_cycle[ 5326] = 1'b1;  addr_rom[ 5326]='h00003cc4;  wr_data_rom[ 5326]='h00002d7f;
    rd_cycle[ 5327] = 1'b1;  wr_cycle[ 5327] = 1'b0;  addr_rom[ 5327]='h000006c4;  wr_data_rom[ 5327]='h00000000;
    rd_cycle[ 5328] = 1'b1;  wr_cycle[ 5328] = 1'b0;  addr_rom[ 5328]='h00002ce4;  wr_data_rom[ 5328]='h00000000;
    rd_cycle[ 5329] = 1'b0;  wr_cycle[ 5329] = 1'b1;  addr_rom[ 5329]='h00001c58;  wr_data_rom[ 5329]='h00001eb9;
    rd_cycle[ 5330] = 1'b1;  wr_cycle[ 5330] = 1'b0;  addr_rom[ 5330]='h000039a4;  wr_data_rom[ 5330]='h00000000;
    rd_cycle[ 5331] = 1'b0;  wr_cycle[ 5331] = 1'b1;  addr_rom[ 5331]='h00003e34;  wr_data_rom[ 5331]='h0000208f;
    rd_cycle[ 5332] = 1'b1;  wr_cycle[ 5332] = 1'b0;  addr_rom[ 5332]='h00001c28;  wr_data_rom[ 5332]='h00000000;
    rd_cycle[ 5333] = 1'b0;  wr_cycle[ 5333] = 1'b1;  addr_rom[ 5333]='h00003e34;  wr_data_rom[ 5333]='h0000150d;
    rd_cycle[ 5334] = 1'b0;  wr_cycle[ 5334] = 1'b1;  addr_rom[ 5334]='h00003c10;  wr_data_rom[ 5334]='h00000684;
    rd_cycle[ 5335] = 1'b0;  wr_cycle[ 5335] = 1'b1;  addr_rom[ 5335]='h00001480;  wr_data_rom[ 5335]='h00003ee7;
    rd_cycle[ 5336] = 1'b1;  wr_cycle[ 5336] = 1'b0;  addr_rom[ 5336]='h00002918;  wr_data_rom[ 5336]='h00000000;
    rd_cycle[ 5337] = 1'b0;  wr_cycle[ 5337] = 1'b1;  addr_rom[ 5337]='h0000382c;  wr_data_rom[ 5337]='h000007f3;
    rd_cycle[ 5338] = 1'b0;  wr_cycle[ 5338] = 1'b1;  addr_rom[ 5338]='h00000d80;  wr_data_rom[ 5338]='h000034fe;
    rd_cycle[ 5339] = 1'b0;  wr_cycle[ 5339] = 1'b1;  addr_rom[ 5339]='h0000384c;  wr_data_rom[ 5339]='h00002e35;
    rd_cycle[ 5340] = 1'b0;  wr_cycle[ 5340] = 1'b1;  addr_rom[ 5340]='h0000064c;  wr_data_rom[ 5340]='h00003918;
    rd_cycle[ 5341] = 1'b1;  wr_cycle[ 5341] = 1'b0;  addr_rom[ 5341]='h00002df0;  wr_data_rom[ 5341]='h00000000;
    rd_cycle[ 5342] = 1'b0;  wr_cycle[ 5342] = 1'b1;  addr_rom[ 5342]='h000027d4;  wr_data_rom[ 5342]='h000029e1;
    rd_cycle[ 5343] = 1'b1;  wr_cycle[ 5343] = 1'b0;  addr_rom[ 5343]='h000028ec;  wr_data_rom[ 5343]='h00000000;
    rd_cycle[ 5344] = 1'b1;  wr_cycle[ 5344] = 1'b0;  addr_rom[ 5344]='h000002a4;  wr_data_rom[ 5344]='h00000000;
    rd_cycle[ 5345] = 1'b1;  wr_cycle[ 5345] = 1'b0;  addr_rom[ 5345]='h00000f50;  wr_data_rom[ 5345]='h00000000;
    rd_cycle[ 5346] = 1'b1;  wr_cycle[ 5346] = 1'b0;  addr_rom[ 5346]='h00000390;  wr_data_rom[ 5346]='h00000000;
    rd_cycle[ 5347] = 1'b0;  wr_cycle[ 5347] = 1'b1;  addr_rom[ 5347]='h00002cb4;  wr_data_rom[ 5347]='h00003001;
    rd_cycle[ 5348] = 1'b1;  wr_cycle[ 5348] = 1'b0;  addr_rom[ 5348]='h000016a8;  wr_data_rom[ 5348]='h00000000;
    rd_cycle[ 5349] = 1'b0;  wr_cycle[ 5349] = 1'b1;  addr_rom[ 5349]='h0000116c;  wr_data_rom[ 5349]='h00003d65;
    rd_cycle[ 5350] = 1'b1;  wr_cycle[ 5350] = 1'b0;  addr_rom[ 5350]='h00003804;  wr_data_rom[ 5350]='h00000000;
    rd_cycle[ 5351] = 1'b1;  wr_cycle[ 5351] = 1'b0;  addr_rom[ 5351]='h00001aa4;  wr_data_rom[ 5351]='h00000000;
    rd_cycle[ 5352] = 1'b1;  wr_cycle[ 5352] = 1'b0;  addr_rom[ 5352]='h000010a4;  wr_data_rom[ 5352]='h00000000;
    rd_cycle[ 5353] = 1'b1;  wr_cycle[ 5353] = 1'b0;  addr_rom[ 5353]='h00000968;  wr_data_rom[ 5353]='h00000000;
    rd_cycle[ 5354] = 1'b1;  wr_cycle[ 5354] = 1'b0;  addr_rom[ 5354]='h000007b4;  wr_data_rom[ 5354]='h00000000;
    rd_cycle[ 5355] = 1'b1;  wr_cycle[ 5355] = 1'b0;  addr_rom[ 5355]='h00002db0;  wr_data_rom[ 5355]='h00000000;
    rd_cycle[ 5356] = 1'b0;  wr_cycle[ 5356] = 1'b1;  addr_rom[ 5356]='h00000a2c;  wr_data_rom[ 5356]='h00003d11;
    rd_cycle[ 5357] = 1'b0;  wr_cycle[ 5357] = 1'b1;  addr_rom[ 5357]='h00002c68;  wr_data_rom[ 5357]='h000025f9;
    rd_cycle[ 5358] = 1'b1;  wr_cycle[ 5358] = 1'b0;  addr_rom[ 5358]='h00002fd8;  wr_data_rom[ 5358]='h00000000;
    rd_cycle[ 5359] = 1'b0;  wr_cycle[ 5359] = 1'b1;  addr_rom[ 5359]='h00003c50;  wr_data_rom[ 5359]='h00002108;
    rd_cycle[ 5360] = 1'b0;  wr_cycle[ 5360] = 1'b1;  addr_rom[ 5360]='h00003894;  wr_data_rom[ 5360]='h00002448;
    rd_cycle[ 5361] = 1'b1;  wr_cycle[ 5361] = 1'b0;  addr_rom[ 5361]='h00001578;  wr_data_rom[ 5361]='h00000000;
    rd_cycle[ 5362] = 1'b0;  wr_cycle[ 5362] = 1'b1;  addr_rom[ 5362]='h0000124c;  wr_data_rom[ 5362]='h000031bc;
    rd_cycle[ 5363] = 1'b1;  wr_cycle[ 5363] = 1'b0;  addr_rom[ 5363]='h00002abc;  wr_data_rom[ 5363]='h00000000;
    rd_cycle[ 5364] = 1'b0;  wr_cycle[ 5364] = 1'b1;  addr_rom[ 5364]='h0000211c;  wr_data_rom[ 5364]='h000019ac;
    rd_cycle[ 5365] = 1'b1;  wr_cycle[ 5365] = 1'b0;  addr_rom[ 5365]='h00001a78;  wr_data_rom[ 5365]='h00000000;
    rd_cycle[ 5366] = 1'b0;  wr_cycle[ 5366] = 1'b1;  addr_rom[ 5366]='h00000910;  wr_data_rom[ 5366]='h00000da9;
    rd_cycle[ 5367] = 1'b1;  wr_cycle[ 5367] = 1'b0;  addr_rom[ 5367]='h000006f0;  wr_data_rom[ 5367]='h00000000;
    rd_cycle[ 5368] = 1'b1;  wr_cycle[ 5368] = 1'b0;  addr_rom[ 5368]='h000026c0;  wr_data_rom[ 5368]='h00000000;
    rd_cycle[ 5369] = 1'b1;  wr_cycle[ 5369] = 1'b0;  addr_rom[ 5369]='h0000110c;  wr_data_rom[ 5369]='h00000000;
    rd_cycle[ 5370] = 1'b0;  wr_cycle[ 5370] = 1'b1;  addr_rom[ 5370]='h00000d2c;  wr_data_rom[ 5370]='h000000ea;
    rd_cycle[ 5371] = 1'b1;  wr_cycle[ 5371] = 1'b0;  addr_rom[ 5371]='h000009c4;  wr_data_rom[ 5371]='h00000000;
    rd_cycle[ 5372] = 1'b0;  wr_cycle[ 5372] = 1'b1;  addr_rom[ 5372]='h00002234;  wr_data_rom[ 5372]='h00001acf;
    rd_cycle[ 5373] = 1'b1;  wr_cycle[ 5373] = 1'b0;  addr_rom[ 5373]='h00002e04;  wr_data_rom[ 5373]='h00000000;
    rd_cycle[ 5374] = 1'b1;  wr_cycle[ 5374] = 1'b0;  addr_rom[ 5374]='h000019e8;  wr_data_rom[ 5374]='h00000000;
    rd_cycle[ 5375] = 1'b0;  wr_cycle[ 5375] = 1'b1;  addr_rom[ 5375]='h0000138c;  wr_data_rom[ 5375]='h000030a5;
    rd_cycle[ 5376] = 1'b1;  wr_cycle[ 5376] = 1'b0;  addr_rom[ 5376]='h00001a78;  wr_data_rom[ 5376]='h00000000;
    rd_cycle[ 5377] = 1'b1;  wr_cycle[ 5377] = 1'b0;  addr_rom[ 5377]='h00003e64;  wr_data_rom[ 5377]='h00000000;
    rd_cycle[ 5378] = 1'b1;  wr_cycle[ 5378] = 1'b0;  addr_rom[ 5378]='h0000166c;  wr_data_rom[ 5378]='h00000000;
    rd_cycle[ 5379] = 1'b1;  wr_cycle[ 5379] = 1'b0;  addr_rom[ 5379]='h00003a54;  wr_data_rom[ 5379]='h00000000;
    rd_cycle[ 5380] = 1'b1;  wr_cycle[ 5380] = 1'b0;  addr_rom[ 5380]='h00003d0c;  wr_data_rom[ 5380]='h00000000;
    rd_cycle[ 5381] = 1'b0;  wr_cycle[ 5381] = 1'b1;  addr_rom[ 5381]='h000033fc;  wr_data_rom[ 5381]='h0000128f;
    rd_cycle[ 5382] = 1'b1;  wr_cycle[ 5382] = 1'b0;  addr_rom[ 5382]='h000027dc;  wr_data_rom[ 5382]='h00000000;
    rd_cycle[ 5383] = 1'b1;  wr_cycle[ 5383] = 1'b0;  addr_rom[ 5383]='h00000ea0;  wr_data_rom[ 5383]='h00000000;
    rd_cycle[ 5384] = 1'b0;  wr_cycle[ 5384] = 1'b1;  addr_rom[ 5384]='h00000538;  wr_data_rom[ 5384]='h00001a86;
    rd_cycle[ 5385] = 1'b1;  wr_cycle[ 5385] = 1'b0;  addr_rom[ 5385]='h000016f0;  wr_data_rom[ 5385]='h00000000;
    rd_cycle[ 5386] = 1'b0;  wr_cycle[ 5386] = 1'b1;  addr_rom[ 5386]='h00000144;  wr_data_rom[ 5386]='h00001c3a;
    rd_cycle[ 5387] = 1'b1;  wr_cycle[ 5387] = 1'b0;  addr_rom[ 5387]='h0000089c;  wr_data_rom[ 5387]='h00000000;
    rd_cycle[ 5388] = 1'b1;  wr_cycle[ 5388] = 1'b0;  addr_rom[ 5388]='h00000590;  wr_data_rom[ 5388]='h00000000;
    rd_cycle[ 5389] = 1'b0;  wr_cycle[ 5389] = 1'b1;  addr_rom[ 5389]='h00003be0;  wr_data_rom[ 5389]='h000035a4;
    rd_cycle[ 5390] = 1'b0;  wr_cycle[ 5390] = 1'b1;  addr_rom[ 5390]='h00003da4;  wr_data_rom[ 5390]='h0000138e;
    rd_cycle[ 5391] = 1'b0;  wr_cycle[ 5391] = 1'b1;  addr_rom[ 5391]='h00002d68;  wr_data_rom[ 5391]='h00002c2d;
    rd_cycle[ 5392] = 1'b1;  wr_cycle[ 5392] = 1'b0;  addr_rom[ 5392]='h00000f68;  wr_data_rom[ 5392]='h00000000;
    rd_cycle[ 5393] = 1'b0;  wr_cycle[ 5393] = 1'b1;  addr_rom[ 5393]='h00000e90;  wr_data_rom[ 5393]='h0000059b;
    rd_cycle[ 5394] = 1'b0;  wr_cycle[ 5394] = 1'b1;  addr_rom[ 5394]='h00001698;  wr_data_rom[ 5394]='h00002763;
    rd_cycle[ 5395] = 1'b1;  wr_cycle[ 5395] = 1'b0;  addr_rom[ 5395]='h000014a0;  wr_data_rom[ 5395]='h00000000;
    rd_cycle[ 5396] = 1'b0;  wr_cycle[ 5396] = 1'b1;  addr_rom[ 5396]='h0000353c;  wr_data_rom[ 5396]='h00001115;
    rd_cycle[ 5397] = 1'b0;  wr_cycle[ 5397] = 1'b1;  addr_rom[ 5397]='h000033cc;  wr_data_rom[ 5397]='h000036cb;
    rd_cycle[ 5398] = 1'b0;  wr_cycle[ 5398] = 1'b1;  addr_rom[ 5398]='h00002094;  wr_data_rom[ 5398]='h00000965;
    rd_cycle[ 5399] = 1'b0;  wr_cycle[ 5399] = 1'b1;  addr_rom[ 5399]='h00000090;  wr_data_rom[ 5399]='h00001a94;
    rd_cycle[ 5400] = 1'b1;  wr_cycle[ 5400] = 1'b0;  addr_rom[ 5400]='h000013e4;  wr_data_rom[ 5400]='h00000000;
    rd_cycle[ 5401] = 1'b0;  wr_cycle[ 5401] = 1'b1;  addr_rom[ 5401]='h000038cc;  wr_data_rom[ 5401]='h00001aad;
    rd_cycle[ 5402] = 1'b1;  wr_cycle[ 5402] = 1'b0;  addr_rom[ 5402]='h00001838;  wr_data_rom[ 5402]='h00000000;
    rd_cycle[ 5403] = 1'b0;  wr_cycle[ 5403] = 1'b1;  addr_rom[ 5403]='h000026f8;  wr_data_rom[ 5403]='h00002953;
    rd_cycle[ 5404] = 1'b0;  wr_cycle[ 5404] = 1'b1;  addr_rom[ 5404]='h00003e24;  wr_data_rom[ 5404]='h000015a5;
    rd_cycle[ 5405] = 1'b1;  wr_cycle[ 5405] = 1'b0;  addr_rom[ 5405]='h000027f8;  wr_data_rom[ 5405]='h00000000;
    rd_cycle[ 5406] = 1'b0;  wr_cycle[ 5406] = 1'b1;  addr_rom[ 5406]='h0000122c;  wr_data_rom[ 5406]='h00001c6a;
    rd_cycle[ 5407] = 1'b0;  wr_cycle[ 5407] = 1'b1;  addr_rom[ 5407]='h000023e8;  wr_data_rom[ 5407]='h00002047;
    rd_cycle[ 5408] = 1'b0;  wr_cycle[ 5408] = 1'b1;  addr_rom[ 5408]='h000001fc;  wr_data_rom[ 5408]='h000038e4;
    rd_cycle[ 5409] = 1'b1;  wr_cycle[ 5409] = 1'b0;  addr_rom[ 5409]='h00002568;  wr_data_rom[ 5409]='h00000000;
    rd_cycle[ 5410] = 1'b1;  wr_cycle[ 5410] = 1'b0;  addr_rom[ 5410]='h00000b30;  wr_data_rom[ 5410]='h00000000;
    rd_cycle[ 5411] = 1'b0;  wr_cycle[ 5411] = 1'b1;  addr_rom[ 5411]='h00003468;  wr_data_rom[ 5411]='h000001ed;
    rd_cycle[ 5412] = 1'b0;  wr_cycle[ 5412] = 1'b1;  addr_rom[ 5412]='h00001978;  wr_data_rom[ 5412]='h000019bc;
    rd_cycle[ 5413] = 1'b1;  wr_cycle[ 5413] = 1'b0;  addr_rom[ 5413]='h0000117c;  wr_data_rom[ 5413]='h00000000;
    rd_cycle[ 5414] = 1'b0;  wr_cycle[ 5414] = 1'b1;  addr_rom[ 5414]='h00002c00;  wr_data_rom[ 5414]='h000039d1;
    rd_cycle[ 5415] = 1'b1;  wr_cycle[ 5415] = 1'b0;  addr_rom[ 5415]='h00002b44;  wr_data_rom[ 5415]='h00000000;
    rd_cycle[ 5416] = 1'b0;  wr_cycle[ 5416] = 1'b1;  addr_rom[ 5416]='h00001df0;  wr_data_rom[ 5416]='h00003f1b;
    rd_cycle[ 5417] = 1'b0;  wr_cycle[ 5417] = 1'b1;  addr_rom[ 5417]='h00000170;  wr_data_rom[ 5417]='h00001893;
    rd_cycle[ 5418] = 1'b0;  wr_cycle[ 5418] = 1'b1;  addr_rom[ 5418]='h00001790;  wr_data_rom[ 5418]='h00002114;
    rd_cycle[ 5419] = 1'b1;  wr_cycle[ 5419] = 1'b0;  addr_rom[ 5419]='h00001850;  wr_data_rom[ 5419]='h00000000;
    rd_cycle[ 5420] = 1'b0;  wr_cycle[ 5420] = 1'b1;  addr_rom[ 5420]='h00001c40;  wr_data_rom[ 5420]='h000000ef;
    rd_cycle[ 5421] = 1'b0;  wr_cycle[ 5421] = 1'b1;  addr_rom[ 5421]='h00003e28;  wr_data_rom[ 5421]='h00001ad0;
    rd_cycle[ 5422] = 1'b1;  wr_cycle[ 5422] = 1'b0;  addr_rom[ 5422]='h000002dc;  wr_data_rom[ 5422]='h00000000;
    rd_cycle[ 5423] = 1'b0;  wr_cycle[ 5423] = 1'b1;  addr_rom[ 5423]='h00002820;  wr_data_rom[ 5423]='h0000310f;
    rd_cycle[ 5424] = 1'b1;  wr_cycle[ 5424] = 1'b0;  addr_rom[ 5424]='h00002388;  wr_data_rom[ 5424]='h00000000;
    rd_cycle[ 5425] = 1'b1;  wr_cycle[ 5425] = 1'b0;  addr_rom[ 5425]='h00002298;  wr_data_rom[ 5425]='h00000000;
    rd_cycle[ 5426] = 1'b0;  wr_cycle[ 5426] = 1'b1;  addr_rom[ 5426]='h00003fa4;  wr_data_rom[ 5426]='h00003138;
    rd_cycle[ 5427] = 1'b1;  wr_cycle[ 5427] = 1'b0;  addr_rom[ 5427]='h00003dc4;  wr_data_rom[ 5427]='h00000000;
    rd_cycle[ 5428] = 1'b0;  wr_cycle[ 5428] = 1'b1;  addr_rom[ 5428]='h000006d8;  wr_data_rom[ 5428]='h00001f1f;
    rd_cycle[ 5429] = 1'b0;  wr_cycle[ 5429] = 1'b1;  addr_rom[ 5429]='h000033d4;  wr_data_rom[ 5429]='h00003cc5;
    rd_cycle[ 5430] = 1'b1;  wr_cycle[ 5430] = 1'b0;  addr_rom[ 5430]='h000002cc;  wr_data_rom[ 5430]='h00000000;
    rd_cycle[ 5431] = 1'b1;  wr_cycle[ 5431] = 1'b0;  addr_rom[ 5431]='h00001490;  wr_data_rom[ 5431]='h00000000;
    rd_cycle[ 5432] = 1'b0;  wr_cycle[ 5432] = 1'b1;  addr_rom[ 5432]='h00003f40;  wr_data_rom[ 5432]='h00000e48;
    rd_cycle[ 5433] = 1'b1;  wr_cycle[ 5433] = 1'b0;  addr_rom[ 5433]='h0000113c;  wr_data_rom[ 5433]='h00000000;
    rd_cycle[ 5434] = 1'b1;  wr_cycle[ 5434] = 1'b0;  addr_rom[ 5434]='h00002ab0;  wr_data_rom[ 5434]='h00000000;
    rd_cycle[ 5435] = 1'b1;  wr_cycle[ 5435] = 1'b0;  addr_rom[ 5435]='h0000137c;  wr_data_rom[ 5435]='h00000000;
    rd_cycle[ 5436] = 1'b1;  wr_cycle[ 5436] = 1'b0;  addr_rom[ 5436]='h00001070;  wr_data_rom[ 5436]='h00000000;
    rd_cycle[ 5437] = 1'b1;  wr_cycle[ 5437] = 1'b0;  addr_rom[ 5437]='h00000b34;  wr_data_rom[ 5437]='h00000000;
    rd_cycle[ 5438] = 1'b1;  wr_cycle[ 5438] = 1'b0;  addr_rom[ 5438]='h000035c0;  wr_data_rom[ 5438]='h00000000;
    rd_cycle[ 5439] = 1'b0;  wr_cycle[ 5439] = 1'b1;  addr_rom[ 5439]='h00003168;  wr_data_rom[ 5439]='h00000657;
    rd_cycle[ 5440] = 1'b0;  wr_cycle[ 5440] = 1'b1;  addr_rom[ 5440]='h0000292c;  wr_data_rom[ 5440]='h00001191;
    rd_cycle[ 5441] = 1'b0;  wr_cycle[ 5441] = 1'b1;  addr_rom[ 5441]='h00002b1c;  wr_data_rom[ 5441]='h0000249e;
    rd_cycle[ 5442] = 1'b1;  wr_cycle[ 5442] = 1'b0;  addr_rom[ 5442]='h00000510;  wr_data_rom[ 5442]='h00000000;
    rd_cycle[ 5443] = 1'b0;  wr_cycle[ 5443] = 1'b1;  addr_rom[ 5443]='h00000dac;  wr_data_rom[ 5443]='h00003b9f;
    rd_cycle[ 5444] = 1'b1;  wr_cycle[ 5444] = 1'b0;  addr_rom[ 5444]='h00003ff8;  wr_data_rom[ 5444]='h00000000;
    rd_cycle[ 5445] = 1'b1;  wr_cycle[ 5445] = 1'b0;  addr_rom[ 5445]='h00002298;  wr_data_rom[ 5445]='h00000000;
    rd_cycle[ 5446] = 1'b0;  wr_cycle[ 5446] = 1'b1;  addr_rom[ 5446]='h00002f24;  wr_data_rom[ 5446]='h0000016e;
    rd_cycle[ 5447] = 1'b1;  wr_cycle[ 5447] = 1'b0;  addr_rom[ 5447]='h00000c1c;  wr_data_rom[ 5447]='h00000000;
    rd_cycle[ 5448] = 1'b1;  wr_cycle[ 5448] = 1'b0;  addr_rom[ 5448]='h0000273c;  wr_data_rom[ 5448]='h00000000;
    rd_cycle[ 5449] = 1'b0;  wr_cycle[ 5449] = 1'b1;  addr_rom[ 5449]='h00001d30;  wr_data_rom[ 5449]='h0000128f;
    rd_cycle[ 5450] = 1'b1;  wr_cycle[ 5450] = 1'b0;  addr_rom[ 5450]='h00001918;  wr_data_rom[ 5450]='h00000000;
    rd_cycle[ 5451] = 1'b0;  wr_cycle[ 5451] = 1'b1;  addr_rom[ 5451]='h00000310;  wr_data_rom[ 5451]='h00002a9d;
    rd_cycle[ 5452] = 1'b0;  wr_cycle[ 5452] = 1'b1;  addr_rom[ 5452]='h00003dc4;  wr_data_rom[ 5452]='h00002941;
    rd_cycle[ 5453] = 1'b1;  wr_cycle[ 5453] = 1'b0;  addr_rom[ 5453]='h00003f88;  wr_data_rom[ 5453]='h00000000;
    rd_cycle[ 5454] = 1'b0;  wr_cycle[ 5454] = 1'b1;  addr_rom[ 5454]='h00000528;  wr_data_rom[ 5454]='h00001dbc;
    rd_cycle[ 5455] = 1'b1;  wr_cycle[ 5455] = 1'b0;  addr_rom[ 5455]='h000006f4;  wr_data_rom[ 5455]='h00000000;
    rd_cycle[ 5456] = 1'b0;  wr_cycle[ 5456] = 1'b1;  addr_rom[ 5456]='h00003880;  wr_data_rom[ 5456]='h00000ecc;
    rd_cycle[ 5457] = 1'b1;  wr_cycle[ 5457] = 1'b0;  addr_rom[ 5457]='h00000f3c;  wr_data_rom[ 5457]='h00000000;
    rd_cycle[ 5458] = 1'b0;  wr_cycle[ 5458] = 1'b1;  addr_rom[ 5458]='h00001308;  wr_data_rom[ 5458]='h0000131b;
    rd_cycle[ 5459] = 1'b0;  wr_cycle[ 5459] = 1'b1;  addr_rom[ 5459]='h000000d0;  wr_data_rom[ 5459]='h00000eb4;
    rd_cycle[ 5460] = 1'b1;  wr_cycle[ 5460] = 1'b0;  addr_rom[ 5460]='h000012d0;  wr_data_rom[ 5460]='h00000000;
    rd_cycle[ 5461] = 1'b0;  wr_cycle[ 5461] = 1'b1;  addr_rom[ 5461]='h00001278;  wr_data_rom[ 5461]='h00002901;
    rd_cycle[ 5462] = 1'b0;  wr_cycle[ 5462] = 1'b1;  addr_rom[ 5462]='h0000108c;  wr_data_rom[ 5462]='h00002a54;
    rd_cycle[ 5463] = 1'b1;  wr_cycle[ 5463] = 1'b0;  addr_rom[ 5463]='h00001f80;  wr_data_rom[ 5463]='h00000000;
    rd_cycle[ 5464] = 1'b0;  wr_cycle[ 5464] = 1'b1;  addr_rom[ 5464]='h00001078;  wr_data_rom[ 5464]='h00003b28;
    rd_cycle[ 5465] = 1'b0;  wr_cycle[ 5465] = 1'b1;  addr_rom[ 5465]='h00003f8c;  wr_data_rom[ 5465]='h00000246;
    rd_cycle[ 5466] = 1'b1;  wr_cycle[ 5466] = 1'b0;  addr_rom[ 5466]='h00003950;  wr_data_rom[ 5466]='h00000000;
    rd_cycle[ 5467] = 1'b1;  wr_cycle[ 5467] = 1'b0;  addr_rom[ 5467]='h000004d8;  wr_data_rom[ 5467]='h00000000;
    rd_cycle[ 5468] = 1'b0;  wr_cycle[ 5468] = 1'b1;  addr_rom[ 5468]='h00001ce4;  wr_data_rom[ 5468]='h00003bdd;
    rd_cycle[ 5469] = 1'b0;  wr_cycle[ 5469] = 1'b1;  addr_rom[ 5469]='h00000510;  wr_data_rom[ 5469]='h000020fe;
    rd_cycle[ 5470] = 1'b0;  wr_cycle[ 5470] = 1'b1;  addr_rom[ 5470]='h000013fc;  wr_data_rom[ 5470]='h00003b90;
    rd_cycle[ 5471] = 1'b1;  wr_cycle[ 5471] = 1'b0;  addr_rom[ 5471]='h00002c4c;  wr_data_rom[ 5471]='h00000000;
    rd_cycle[ 5472] = 1'b0;  wr_cycle[ 5472] = 1'b1;  addr_rom[ 5472]='h00000b74;  wr_data_rom[ 5472]='h00003601;
    rd_cycle[ 5473] = 1'b0;  wr_cycle[ 5473] = 1'b1;  addr_rom[ 5473]='h0000364c;  wr_data_rom[ 5473]='h000003b1;
    rd_cycle[ 5474] = 1'b1;  wr_cycle[ 5474] = 1'b0;  addr_rom[ 5474]='h000017c8;  wr_data_rom[ 5474]='h00000000;
    rd_cycle[ 5475] = 1'b0;  wr_cycle[ 5475] = 1'b1;  addr_rom[ 5475]='h0000053c;  wr_data_rom[ 5475]='h00000450;
    rd_cycle[ 5476] = 1'b0;  wr_cycle[ 5476] = 1'b1;  addr_rom[ 5476]='h00001544;  wr_data_rom[ 5476]='h0000131e;
    rd_cycle[ 5477] = 1'b0;  wr_cycle[ 5477] = 1'b1;  addr_rom[ 5477]='h000008bc;  wr_data_rom[ 5477]='h00003f46;
    rd_cycle[ 5478] = 1'b0;  wr_cycle[ 5478] = 1'b1;  addr_rom[ 5478]='h00003098;  wr_data_rom[ 5478]='h00000542;
    rd_cycle[ 5479] = 1'b1;  wr_cycle[ 5479] = 1'b0;  addr_rom[ 5479]='h00001b84;  wr_data_rom[ 5479]='h00000000;
    rd_cycle[ 5480] = 1'b1;  wr_cycle[ 5480] = 1'b0;  addr_rom[ 5480]='h000002c8;  wr_data_rom[ 5480]='h00000000;
    rd_cycle[ 5481] = 1'b1;  wr_cycle[ 5481] = 1'b0;  addr_rom[ 5481]='h00002cf8;  wr_data_rom[ 5481]='h00000000;
    rd_cycle[ 5482] = 1'b0;  wr_cycle[ 5482] = 1'b1;  addr_rom[ 5482]='h0000093c;  wr_data_rom[ 5482]='h000033fb;
    rd_cycle[ 5483] = 1'b1;  wr_cycle[ 5483] = 1'b0;  addr_rom[ 5483]='h00001860;  wr_data_rom[ 5483]='h00000000;
    rd_cycle[ 5484] = 1'b0;  wr_cycle[ 5484] = 1'b1;  addr_rom[ 5484]='h00000bdc;  wr_data_rom[ 5484]='h00000c9b;
    rd_cycle[ 5485] = 1'b1;  wr_cycle[ 5485] = 1'b0;  addr_rom[ 5485]='h000000c4;  wr_data_rom[ 5485]='h00000000;
    rd_cycle[ 5486] = 1'b1;  wr_cycle[ 5486] = 1'b0;  addr_rom[ 5486]='h00000d50;  wr_data_rom[ 5486]='h00000000;
    rd_cycle[ 5487] = 1'b1;  wr_cycle[ 5487] = 1'b0;  addr_rom[ 5487]='h00002ea4;  wr_data_rom[ 5487]='h00000000;
    rd_cycle[ 5488] = 1'b1;  wr_cycle[ 5488] = 1'b0;  addr_rom[ 5488]='h00003388;  wr_data_rom[ 5488]='h00000000;
    rd_cycle[ 5489] = 1'b1;  wr_cycle[ 5489] = 1'b0;  addr_rom[ 5489]='h0000145c;  wr_data_rom[ 5489]='h00000000;
    rd_cycle[ 5490] = 1'b0;  wr_cycle[ 5490] = 1'b1;  addr_rom[ 5490]='h00000a9c;  wr_data_rom[ 5490]='h00001902;
    rd_cycle[ 5491] = 1'b0;  wr_cycle[ 5491] = 1'b1;  addr_rom[ 5491]='h00001790;  wr_data_rom[ 5491]='h00000178;
    rd_cycle[ 5492] = 1'b0;  wr_cycle[ 5492] = 1'b1;  addr_rom[ 5492]='h000025c4;  wr_data_rom[ 5492]='h00001d9f;
    rd_cycle[ 5493] = 1'b0;  wr_cycle[ 5493] = 1'b1;  addr_rom[ 5493]='h000018cc;  wr_data_rom[ 5493]='h000028e9;
    rd_cycle[ 5494] = 1'b1;  wr_cycle[ 5494] = 1'b0;  addr_rom[ 5494]='h00000728;  wr_data_rom[ 5494]='h00000000;
    rd_cycle[ 5495] = 1'b1;  wr_cycle[ 5495] = 1'b0;  addr_rom[ 5495]='h00001ac4;  wr_data_rom[ 5495]='h00000000;
    rd_cycle[ 5496] = 1'b0;  wr_cycle[ 5496] = 1'b1;  addr_rom[ 5496]='h00000180;  wr_data_rom[ 5496]='h00002042;
    rd_cycle[ 5497] = 1'b1;  wr_cycle[ 5497] = 1'b0;  addr_rom[ 5497]='h00000b5c;  wr_data_rom[ 5497]='h00000000;
    rd_cycle[ 5498] = 1'b1;  wr_cycle[ 5498] = 1'b0;  addr_rom[ 5498]='h00002c90;  wr_data_rom[ 5498]='h00000000;
    rd_cycle[ 5499] = 1'b0;  wr_cycle[ 5499] = 1'b1;  addr_rom[ 5499]='h000038a0;  wr_data_rom[ 5499]='h000018ac;
    rd_cycle[ 5500] = 1'b1;  wr_cycle[ 5500] = 1'b0;  addr_rom[ 5500]='h000025e0;  wr_data_rom[ 5500]='h00000000;
    rd_cycle[ 5501] = 1'b0;  wr_cycle[ 5501] = 1'b1;  addr_rom[ 5501]='h00003020;  wr_data_rom[ 5501]='h00000f3a;
    rd_cycle[ 5502] = 1'b1;  wr_cycle[ 5502] = 1'b0;  addr_rom[ 5502]='h00002bf8;  wr_data_rom[ 5502]='h00000000;
    rd_cycle[ 5503] = 1'b1;  wr_cycle[ 5503] = 1'b0;  addr_rom[ 5503]='h00002920;  wr_data_rom[ 5503]='h00000000;
    rd_cycle[ 5504] = 1'b0;  wr_cycle[ 5504] = 1'b1;  addr_rom[ 5504]='h00003720;  wr_data_rom[ 5504]='h0000187f;
    rd_cycle[ 5505] = 1'b1;  wr_cycle[ 5505] = 1'b0;  addr_rom[ 5505]='h00002610;  wr_data_rom[ 5505]='h00000000;
    rd_cycle[ 5506] = 1'b0;  wr_cycle[ 5506] = 1'b1;  addr_rom[ 5506]='h00003c30;  wr_data_rom[ 5506]='h000005f4;
    rd_cycle[ 5507] = 1'b1;  wr_cycle[ 5507] = 1'b0;  addr_rom[ 5507]='h00001f1c;  wr_data_rom[ 5507]='h00000000;
    rd_cycle[ 5508] = 1'b1;  wr_cycle[ 5508] = 1'b0;  addr_rom[ 5508]='h00003f00;  wr_data_rom[ 5508]='h00000000;
    rd_cycle[ 5509] = 1'b1;  wr_cycle[ 5509] = 1'b0;  addr_rom[ 5509]='h00003b74;  wr_data_rom[ 5509]='h00000000;
    rd_cycle[ 5510] = 1'b0;  wr_cycle[ 5510] = 1'b1;  addr_rom[ 5510]='h000002f8;  wr_data_rom[ 5510]='h00002263;
    rd_cycle[ 5511] = 1'b0;  wr_cycle[ 5511] = 1'b1;  addr_rom[ 5511]='h00000730;  wr_data_rom[ 5511]='h00000a54;
    rd_cycle[ 5512] = 1'b1;  wr_cycle[ 5512] = 1'b0;  addr_rom[ 5512]='h00002f18;  wr_data_rom[ 5512]='h00000000;
    rd_cycle[ 5513] = 1'b1;  wr_cycle[ 5513] = 1'b0;  addr_rom[ 5513]='h00000ca4;  wr_data_rom[ 5513]='h00000000;
    rd_cycle[ 5514] = 1'b0;  wr_cycle[ 5514] = 1'b1;  addr_rom[ 5514]='h00000380;  wr_data_rom[ 5514]='h00001340;
    rd_cycle[ 5515] = 1'b1;  wr_cycle[ 5515] = 1'b0;  addr_rom[ 5515]='h000026a4;  wr_data_rom[ 5515]='h00000000;
    rd_cycle[ 5516] = 1'b1;  wr_cycle[ 5516] = 1'b0;  addr_rom[ 5516]='h00001854;  wr_data_rom[ 5516]='h00000000;
    rd_cycle[ 5517] = 1'b0;  wr_cycle[ 5517] = 1'b1;  addr_rom[ 5517]='h00001ca8;  wr_data_rom[ 5517]='h0000128f;
    rd_cycle[ 5518] = 1'b0;  wr_cycle[ 5518] = 1'b1;  addr_rom[ 5518]='h000025d4;  wr_data_rom[ 5518]='h000038e8;
    rd_cycle[ 5519] = 1'b0;  wr_cycle[ 5519] = 1'b1;  addr_rom[ 5519]='h00001170;  wr_data_rom[ 5519]='h00003e50;
    rd_cycle[ 5520] = 1'b1;  wr_cycle[ 5520] = 1'b0;  addr_rom[ 5520]='h000024e0;  wr_data_rom[ 5520]='h00000000;
    rd_cycle[ 5521] = 1'b0;  wr_cycle[ 5521] = 1'b1;  addr_rom[ 5521]='h00000cac;  wr_data_rom[ 5521]='h00001b91;
    rd_cycle[ 5522] = 1'b0;  wr_cycle[ 5522] = 1'b1;  addr_rom[ 5522]='h000025f8;  wr_data_rom[ 5522]='h0000333a;
    rd_cycle[ 5523] = 1'b0;  wr_cycle[ 5523] = 1'b1;  addr_rom[ 5523]='h0000385c;  wr_data_rom[ 5523]='h000033f6;
    rd_cycle[ 5524] = 1'b1;  wr_cycle[ 5524] = 1'b0;  addr_rom[ 5524]='h00001c24;  wr_data_rom[ 5524]='h00000000;
    rd_cycle[ 5525] = 1'b0;  wr_cycle[ 5525] = 1'b1;  addr_rom[ 5525]='h00003f90;  wr_data_rom[ 5525]='h00002076;
    rd_cycle[ 5526] = 1'b1;  wr_cycle[ 5526] = 1'b0;  addr_rom[ 5526]='h000034ec;  wr_data_rom[ 5526]='h00000000;
    rd_cycle[ 5527] = 1'b0;  wr_cycle[ 5527] = 1'b1;  addr_rom[ 5527]='h00001d18;  wr_data_rom[ 5527]='h00000fd2;
    rd_cycle[ 5528] = 1'b0;  wr_cycle[ 5528] = 1'b1;  addr_rom[ 5528]='h00003934;  wr_data_rom[ 5528]='h00002c65;
    rd_cycle[ 5529] = 1'b1;  wr_cycle[ 5529] = 1'b0;  addr_rom[ 5529]='h000017c4;  wr_data_rom[ 5529]='h00000000;
    rd_cycle[ 5530] = 1'b0;  wr_cycle[ 5530] = 1'b1;  addr_rom[ 5530]='h00002068;  wr_data_rom[ 5530]='h00000209;
    rd_cycle[ 5531] = 1'b1;  wr_cycle[ 5531] = 1'b0;  addr_rom[ 5531]='h00001528;  wr_data_rom[ 5531]='h00000000;
    rd_cycle[ 5532] = 1'b1;  wr_cycle[ 5532] = 1'b0;  addr_rom[ 5532]='h00001a50;  wr_data_rom[ 5532]='h00000000;
    rd_cycle[ 5533] = 1'b1;  wr_cycle[ 5533] = 1'b0;  addr_rom[ 5533]='h00002efc;  wr_data_rom[ 5533]='h00000000;
    rd_cycle[ 5534] = 1'b1;  wr_cycle[ 5534] = 1'b0;  addr_rom[ 5534]='h00003ad4;  wr_data_rom[ 5534]='h00000000;
    rd_cycle[ 5535] = 1'b0;  wr_cycle[ 5535] = 1'b1;  addr_rom[ 5535]='h00001238;  wr_data_rom[ 5535]='h00000f58;
    rd_cycle[ 5536] = 1'b0;  wr_cycle[ 5536] = 1'b1;  addr_rom[ 5536]='h00003834;  wr_data_rom[ 5536]='h000001d6;
    rd_cycle[ 5537] = 1'b1;  wr_cycle[ 5537] = 1'b0;  addr_rom[ 5537]='h000020ec;  wr_data_rom[ 5537]='h00000000;
    rd_cycle[ 5538] = 1'b1;  wr_cycle[ 5538] = 1'b0;  addr_rom[ 5538]='h00003728;  wr_data_rom[ 5538]='h00000000;
    rd_cycle[ 5539] = 1'b0;  wr_cycle[ 5539] = 1'b1;  addr_rom[ 5539]='h00001af0;  wr_data_rom[ 5539]='h00002c11;
    rd_cycle[ 5540] = 1'b1;  wr_cycle[ 5540] = 1'b0;  addr_rom[ 5540]='h00002224;  wr_data_rom[ 5540]='h00000000;
    rd_cycle[ 5541] = 1'b1;  wr_cycle[ 5541] = 1'b0;  addr_rom[ 5541]='h000017a4;  wr_data_rom[ 5541]='h00000000;
    rd_cycle[ 5542] = 1'b1;  wr_cycle[ 5542] = 1'b0;  addr_rom[ 5542]='h00001c00;  wr_data_rom[ 5542]='h00000000;
    rd_cycle[ 5543] = 1'b1;  wr_cycle[ 5543] = 1'b0;  addr_rom[ 5543]='h00002c88;  wr_data_rom[ 5543]='h00000000;
    rd_cycle[ 5544] = 1'b0;  wr_cycle[ 5544] = 1'b1;  addr_rom[ 5544]='h000029fc;  wr_data_rom[ 5544]='h0000324e;
    rd_cycle[ 5545] = 1'b1;  wr_cycle[ 5545] = 1'b0;  addr_rom[ 5545]='h00003f44;  wr_data_rom[ 5545]='h00000000;
    rd_cycle[ 5546] = 1'b0;  wr_cycle[ 5546] = 1'b1;  addr_rom[ 5546]='h000015d8;  wr_data_rom[ 5546]='h00001a96;
    rd_cycle[ 5547] = 1'b0;  wr_cycle[ 5547] = 1'b1;  addr_rom[ 5547]='h0000388c;  wr_data_rom[ 5547]='h00003c6d;
    rd_cycle[ 5548] = 1'b0;  wr_cycle[ 5548] = 1'b1;  addr_rom[ 5548]='h00002b48;  wr_data_rom[ 5548]='h00002b0e;
    rd_cycle[ 5549] = 1'b0;  wr_cycle[ 5549] = 1'b1;  addr_rom[ 5549]='h00003ec0;  wr_data_rom[ 5549]='h00002665;
    rd_cycle[ 5550] = 1'b0;  wr_cycle[ 5550] = 1'b1;  addr_rom[ 5550]='h00001294;  wr_data_rom[ 5550]='h00000d9d;
    rd_cycle[ 5551] = 1'b0;  wr_cycle[ 5551] = 1'b1;  addr_rom[ 5551]='h00002728;  wr_data_rom[ 5551]='h00001947;
    rd_cycle[ 5552] = 1'b1;  wr_cycle[ 5552] = 1'b0;  addr_rom[ 5552]='h00002294;  wr_data_rom[ 5552]='h00000000;
    rd_cycle[ 5553] = 1'b0;  wr_cycle[ 5553] = 1'b1;  addr_rom[ 5553]='h00003638;  wr_data_rom[ 5553]='h000020ae;
    rd_cycle[ 5554] = 1'b0;  wr_cycle[ 5554] = 1'b1;  addr_rom[ 5554]='h000008c0;  wr_data_rom[ 5554]='h00000303;
    rd_cycle[ 5555] = 1'b0;  wr_cycle[ 5555] = 1'b1;  addr_rom[ 5555]='h00003bdc;  wr_data_rom[ 5555]='h000017e4;
    rd_cycle[ 5556] = 1'b0;  wr_cycle[ 5556] = 1'b1;  addr_rom[ 5556]='h00000564;  wr_data_rom[ 5556]='h0000054e;
    rd_cycle[ 5557] = 1'b1;  wr_cycle[ 5557] = 1'b0;  addr_rom[ 5557]='h0000219c;  wr_data_rom[ 5557]='h00000000;
    rd_cycle[ 5558] = 1'b1;  wr_cycle[ 5558] = 1'b0;  addr_rom[ 5558]='h00003e6c;  wr_data_rom[ 5558]='h00000000;
    rd_cycle[ 5559] = 1'b1;  wr_cycle[ 5559] = 1'b0;  addr_rom[ 5559]='h000038a0;  wr_data_rom[ 5559]='h00000000;
    rd_cycle[ 5560] = 1'b0;  wr_cycle[ 5560] = 1'b1;  addr_rom[ 5560]='h000023ec;  wr_data_rom[ 5560]='h00003a0a;
    rd_cycle[ 5561] = 1'b0;  wr_cycle[ 5561] = 1'b1;  addr_rom[ 5561]='h0000055c;  wr_data_rom[ 5561]='h00002458;
    rd_cycle[ 5562] = 1'b0;  wr_cycle[ 5562] = 1'b1;  addr_rom[ 5562]='h00000c28;  wr_data_rom[ 5562]='h00002506;
    rd_cycle[ 5563] = 1'b0;  wr_cycle[ 5563] = 1'b1;  addr_rom[ 5563]='h00003430;  wr_data_rom[ 5563]='h0000302f;
    rd_cycle[ 5564] = 1'b1;  wr_cycle[ 5564] = 1'b0;  addr_rom[ 5564]='h000028a8;  wr_data_rom[ 5564]='h00000000;
    rd_cycle[ 5565] = 1'b1;  wr_cycle[ 5565] = 1'b0;  addr_rom[ 5565]='h00002ef4;  wr_data_rom[ 5565]='h00000000;
    rd_cycle[ 5566] = 1'b0;  wr_cycle[ 5566] = 1'b1;  addr_rom[ 5566]='h000035b4;  wr_data_rom[ 5566]='h00000eb2;
    rd_cycle[ 5567] = 1'b0;  wr_cycle[ 5567] = 1'b1;  addr_rom[ 5567]='h000034ac;  wr_data_rom[ 5567]='h00000115;
    rd_cycle[ 5568] = 1'b0;  wr_cycle[ 5568] = 1'b1;  addr_rom[ 5568]='h00000e28;  wr_data_rom[ 5568]='h00001217;
    rd_cycle[ 5569] = 1'b1;  wr_cycle[ 5569] = 1'b0;  addr_rom[ 5569]='h0000126c;  wr_data_rom[ 5569]='h00000000;
    rd_cycle[ 5570] = 1'b1;  wr_cycle[ 5570] = 1'b0;  addr_rom[ 5570]='h00002b3c;  wr_data_rom[ 5570]='h00000000;
    rd_cycle[ 5571] = 1'b0;  wr_cycle[ 5571] = 1'b1;  addr_rom[ 5571]='h0000363c;  wr_data_rom[ 5571]='h00000a97;
    rd_cycle[ 5572] = 1'b0;  wr_cycle[ 5572] = 1'b1;  addr_rom[ 5572]='h00002844;  wr_data_rom[ 5572]='h000024cf;
    rd_cycle[ 5573] = 1'b0;  wr_cycle[ 5573] = 1'b1;  addr_rom[ 5573]='h0000233c;  wr_data_rom[ 5573]='h00003681;
    rd_cycle[ 5574] = 1'b0;  wr_cycle[ 5574] = 1'b1;  addr_rom[ 5574]='h00001d84;  wr_data_rom[ 5574]='h00003467;
    rd_cycle[ 5575] = 1'b0;  wr_cycle[ 5575] = 1'b1;  addr_rom[ 5575]='h00000170;  wr_data_rom[ 5575]='h0000261c;
    rd_cycle[ 5576] = 1'b1;  wr_cycle[ 5576] = 1'b0;  addr_rom[ 5576]='h0000207c;  wr_data_rom[ 5576]='h00000000;
    rd_cycle[ 5577] = 1'b0;  wr_cycle[ 5577] = 1'b1;  addr_rom[ 5577]='h00002810;  wr_data_rom[ 5577]='h000034d3;
    rd_cycle[ 5578] = 1'b0;  wr_cycle[ 5578] = 1'b1;  addr_rom[ 5578]='h00002720;  wr_data_rom[ 5578]='h00001713;
    rd_cycle[ 5579] = 1'b0;  wr_cycle[ 5579] = 1'b1;  addr_rom[ 5579]='h00000b24;  wr_data_rom[ 5579]='h00003815;
    rd_cycle[ 5580] = 1'b0;  wr_cycle[ 5580] = 1'b1;  addr_rom[ 5580]='h00003ce4;  wr_data_rom[ 5580]='h00000b8e;
    rd_cycle[ 5581] = 1'b1;  wr_cycle[ 5581] = 1'b0;  addr_rom[ 5581]='h000031bc;  wr_data_rom[ 5581]='h00000000;
    rd_cycle[ 5582] = 1'b0;  wr_cycle[ 5582] = 1'b1;  addr_rom[ 5582]='h00001698;  wr_data_rom[ 5582]='h00003815;
    rd_cycle[ 5583] = 1'b1;  wr_cycle[ 5583] = 1'b0;  addr_rom[ 5583]='h00002ac8;  wr_data_rom[ 5583]='h00000000;
    rd_cycle[ 5584] = 1'b0;  wr_cycle[ 5584] = 1'b1;  addr_rom[ 5584]='h00001ed4;  wr_data_rom[ 5584]='h00001b44;
    rd_cycle[ 5585] = 1'b0;  wr_cycle[ 5585] = 1'b1;  addr_rom[ 5585]='h00001f58;  wr_data_rom[ 5585]='h0000330d;
    rd_cycle[ 5586] = 1'b0;  wr_cycle[ 5586] = 1'b1;  addr_rom[ 5586]='h000018fc;  wr_data_rom[ 5586]='h00003010;
    rd_cycle[ 5587] = 1'b1;  wr_cycle[ 5587] = 1'b0;  addr_rom[ 5587]='h000000e8;  wr_data_rom[ 5587]='h00000000;
    rd_cycle[ 5588] = 1'b0;  wr_cycle[ 5588] = 1'b1;  addr_rom[ 5588]='h000033c4;  wr_data_rom[ 5588]='h00001f57;
    rd_cycle[ 5589] = 1'b1;  wr_cycle[ 5589] = 1'b0;  addr_rom[ 5589]='h00003e94;  wr_data_rom[ 5589]='h00000000;
    rd_cycle[ 5590] = 1'b0;  wr_cycle[ 5590] = 1'b1;  addr_rom[ 5590]='h00002f04;  wr_data_rom[ 5590]='h00000a00;
    rd_cycle[ 5591] = 1'b1;  wr_cycle[ 5591] = 1'b0;  addr_rom[ 5591]='h00002140;  wr_data_rom[ 5591]='h00000000;
    rd_cycle[ 5592] = 1'b0;  wr_cycle[ 5592] = 1'b1;  addr_rom[ 5592]='h0000210c;  wr_data_rom[ 5592]='h00002daf;
    rd_cycle[ 5593] = 1'b1;  wr_cycle[ 5593] = 1'b0;  addr_rom[ 5593]='h00000a04;  wr_data_rom[ 5593]='h00000000;
    rd_cycle[ 5594] = 1'b0;  wr_cycle[ 5594] = 1'b1;  addr_rom[ 5594]='h0000106c;  wr_data_rom[ 5594]='h00003cd6;
    rd_cycle[ 5595] = 1'b1;  wr_cycle[ 5595] = 1'b0;  addr_rom[ 5595]='h00002f50;  wr_data_rom[ 5595]='h00000000;
    rd_cycle[ 5596] = 1'b1;  wr_cycle[ 5596] = 1'b0;  addr_rom[ 5596]='h00003088;  wr_data_rom[ 5596]='h00000000;
    rd_cycle[ 5597] = 1'b1;  wr_cycle[ 5597] = 1'b0;  addr_rom[ 5597]='h000034b8;  wr_data_rom[ 5597]='h00000000;
    rd_cycle[ 5598] = 1'b0;  wr_cycle[ 5598] = 1'b1;  addr_rom[ 5598]='h00000df8;  wr_data_rom[ 5598]='h0000153b;
    rd_cycle[ 5599] = 1'b1;  wr_cycle[ 5599] = 1'b0;  addr_rom[ 5599]='h00000c9c;  wr_data_rom[ 5599]='h00000000;
    rd_cycle[ 5600] = 1'b1;  wr_cycle[ 5600] = 1'b0;  addr_rom[ 5600]='h000017b4;  wr_data_rom[ 5600]='h00000000;
    rd_cycle[ 5601] = 1'b0;  wr_cycle[ 5601] = 1'b1;  addr_rom[ 5601]='h00003cf8;  wr_data_rom[ 5601]='h00001ca9;
    rd_cycle[ 5602] = 1'b0;  wr_cycle[ 5602] = 1'b1;  addr_rom[ 5602]='h00000298;  wr_data_rom[ 5602]='h00003b4e;
    rd_cycle[ 5603] = 1'b0;  wr_cycle[ 5603] = 1'b1;  addr_rom[ 5603]='h000019a4;  wr_data_rom[ 5603]='h00003c73;
    rd_cycle[ 5604] = 1'b0;  wr_cycle[ 5604] = 1'b1;  addr_rom[ 5604]='h00001324;  wr_data_rom[ 5604]='h00000c17;
    rd_cycle[ 5605] = 1'b0;  wr_cycle[ 5605] = 1'b1;  addr_rom[ 5605]='h00002e94;  wr_data_rom[ 5605]='h0000059b;
    rd_cycle[ 5606] = 1'b0;  wr_cycle[ 5606] = 1'b1;  addr_rom[ 5606]='h000020f8;  wr_data_rom[ 5606]='h00003c28;
    rd_cycle[ 5607] = 1'b0;  wr_cycle[ 5607] = 1'b1;  addr_rom[ 5607]='h000016ac;  wr_data_rom[ 5607]='h000005db;
    rd_cycle[ 5608] = 1'b0;  wr_cycle[ 5608] = 1'b1;  addr_rom[ 5608]='h00000ed8;  wr_data_rom[ 5608]='h00001d6d;
    rd_cycle[ 5609] = 1'b0;  wr_cycle[ 5609] = 1'b1;  addr_rom[ 5609]='h00001454;  wr_data_rom[ 5609]='h00002484;
    rd_cycle[ 5610] = 1'b0;  wr_cycle[ 5610] = 1'b1;  addr_rom[ 5610]='h0000202c;  wr_data_rom[ 5610]='h00003b22;
    rd_cycle[ 5611] = 1'b0;  wr_cycle[ 5611] = 1'b1;  addr_rom[ 5611]='h000038dc;  wr_data_rom[ 5611]='h00001bd6;
    rd_cycle[ 5612] = 1'b1;  wr_cycle[ 5612] = 1'b0;  addr_rom[ 5612]='h000020fc;  wr_data_rom[ 5612]='h00000000;
    rd_cycle[ 5613] = 1'b0;  wr_cycle[ 5613] = 1'b1;  addr_rom[ 5613]='h00002200;  wr_data_rom[ 5613]='h000000b2;
    rd_cycle[ 5614] = 1'b0;  wr_cycle[ 5614] = 1'b1;  addr_rom[ 5614]='h000010a8;  wr_data_rom[ 5614]='h000014c8;
    rd_cycle[ 5615] = 1'b0;  wr_cycle[ 5615] = 1'b1;  addr_rom[ 5615]='h0000251c;  wr_data_rom[ 5615]='h00002737;
    rd_cycle[ 5616] = 1'b1;  wr_cycle[ 5616] = 1'b0;  addr_rom[ 5616]='h00000620;  wr_data_rom[ 5616]='h00000000;
    rd_cycle[ 5617] = 1'b1;  wr_cycle[ 5617] = 1'b0;  addr_rom[ 5617]='h00002368;  wr_data_rom[ 5617]='h00000000;
    rd_cycle[ 5618] = 1'b0;  wr_cycle[ 5618] = 1'b1;  addr_rom[ 5618]='h000020f4;  wr_data_rom[ 5618]='h00000964;
    rd_cycle[ 5619] = 1'b1;  wr_cycle[ 5619] = 1'b0;  addr_rom[ 5619]='h00000b04;  wr_data_rom[ 5619]='h00000000;
    rd_cycle[ 5620] = 1'b0;  wr_cycle[ 5620] = 1'b1;  addr_rom[ 5620]='h00001710;  wr_data_rom[ 5620]='h000012f2;
    rd_cycle[ 5621] = 1'b0;  wr_cycle[ 5621] = 1'b1;  addr_rom[ 5621]='h00003328;  wr_data_rom[ 5621]='h00002411;
    rd_cycle[ 5622] = 1'b1;  wr_cycle[ 5622] = 1'b0;  addr_rom[ 5622]='h000024dc;  wr_data_rom[ 5622]='h00000000;
    rd_cycle[ 5623] = 1'b0;  wr_cycle[ 5623] = 1'b1;  addr_rom[ 5623]='h00001dd4;  wr_data_rom[ 5623]='h0000258c;
    rd_cycle[ 5624] = 1'b0;  wr_cycle[ 5624] = 1'b1;  addr_rom[ 5624]='h00003b90;  wr_data_rom[ 5624]='h00002a33;
    rd_cycle[ 5625] = 1'b1;  wr_cycle[ 5625] = 1'b0;  addr_rom[ 5625]='h00002b80;  wr_data_rom[ 5625]='h00000000;
    rd_cycle[ 5626] = 1'b1;  wr_cycle[ 5626] = 1'b0;  addr_rom[ 5626]='h00002ce4;  wr_data_rom[ 5626]='h00000000;
    rd_cycle[ 5627] = 1'b1;  wr_cycle[ 5627] = 1'b0;  addr_rom[ 5627]='h000028ec;  wr_data_rom[ 5627]='h00000000;
    rd_cycle[ 5628] = 1'b0;  wr_cycle[ 5628] = 1'b1;  addr_rom[ 5628]='h00002430;  wr_data_rom[ 5628]='h00001268;
    rd_cycle[ 5629] = 1'b0;  wr_cycle[ 5629] = 1'b1;  addr_rom[ 5629]='h00002074;  wr_data_rom[ 5629]='h000036e5;
    rd_cycle[ 5630] = 1'b0;  wr_cycle[ 5630] = 1'b1;  addr_rom[ 5630]='h00001cf4;  wr_data_rom[ 5630]='h00003859;
    rd_cycle[ 5631] = 1'b1;  wr_cycle[ 5631] = 1'b0;  addr_rom[ 5631]='h00000b50;  wr_data_rom[ 5631]='h00000000;
    rd_cycle[ 5632] = 1'b0;  wr_cycle[ 5632] = 1'b1;  addr_rom[ 5632]='h00003090;  wr_data_rom[ 5632]='h00003b57;
    rd_cycle[ 5633] = 1'b0;  wr_cycle[ 5633] = 1'b1;  addr_rom[ 5633]='h00002d10;  wr_data_rom[ 5633]='h00003477;
    rd_cycle[ 5634] = 1'b0;  wr_cycle[ 5634] = 1'b1;  addr_rom[ 5634]='h00002a10;  wr_data_rom[ 5634]='h00001f45;
    rd_cycle[ 5635] = 1'b1;  wr_cycle[ 5635] = 1'b0;  addr_rom[ 5635]='h00000bd4;  wr_data_rom[ 5635]='h00000000;
    rd_cycle[ 5636] = 1'b0;  wr_cycle[ 5636] = 1'b1;  addr_rom[ 5636]='h00001e3c;  wr_data_rom[ 5636]='h00001ccb;
    rd_cycle[ 5637] = 1'b0;  wr_cycle[ 5637] = 1'b1;  addr_rom[ 5637]='h000011a0;  wr_data_rom[ 5637]='h00002ab6;
    rd_cycle[ 5638] = 1'b0;  wr_cycle[ 5638] = 1'b1;  addr_rom[ 5638]='h000011f8;  wr_data_rom[ 5638]='h0000105f;
    rd_cycle[ 5639] = 1'b0;  wr_cycle[ 5639] = 1'b1;  addr_rom[ 5639]='h00000868;  wr_data_rom[ 5639]='h0000073a;
    rd_cycle[ 5640] = 1'b1;  wr_cycle[ 5640] = 1'b0;  addr_rom[ 5640]='h00002e10;  wr_data_rom[ 5640]='h00000000;
    rd_cycle[ 5641] = 1'b0;  wr_cycle[ 5641] = 1'b1;  addr_rom[ 5641]='h00002874;  wr_data_rom[ 5641]='h000039a5;
    rd_cycle[ 5642] = 1'b0;  wr_cycle[ 5642] = 1'b1;  addr_rom[ 5642]='h0000172c;  wr_data_rom[ 5642]='h00003e91;
    rd_cycle[ 5643] = 1'b1;  wr_cycle[ 5643] = 1'b0;  addr_rom[ 5643]='h000010b0;  wr_data_rom[ 5643]='h00000000;
    rd_cycle[ 5644] = 1'b1;  wr_cycle[ 5644] = 1'b0;  addr_rom[ 5644]='h00000710;  wr_data_rom[ 5644]='h00000000;
    rd_cycle[ 5645] = 1'b1;  wr_cycle[ 5645] = 1'b0;  addr_rom[ 5645]='h00002bd8;  wr_data_rom[ 5645]='h00000000;
    rd_cycle[ 5646] = 1'b1;  wr_cycle[ 5646] = 1'b0;  addr_rom[ 5646]='h0000331c;  wr_data_rom[ 5646]='h00000000;
    rd_cycle[ 5647] = 1'b0;  wr_cycle[ 5647] = 1'b1;  addr_rom[ 5647]='h00003dfc;  wr_data_rom[ 5647]='h00003c1b;
    rd_cycle[ 5648] = 1'b0;  wr_cycle[ 5648] = 1'b1;  addr_rom[ 5648]='h00001370;  wr_data_rom[ 5648]='h00001efa;
    rd_cycle[ 5649] = 1'b0;  wr_cycle[ 5649] = 1'b1;  addr_rom[ 5649]='h00000158;  wr_data_rom[ 5649]='h00003061;
    rd_cycle[ 5650] = 1'b0;  wr_cycle[ 5650] = 1'b1;  addr_rom[ 5650]='h00003398;  wr_data_rom[ 5650]='h00000220;
    rd_cycle[ 5651] = 1'b0;  wr_cycle[ 5651] = 1'b1;  addr_rom[ 5651]='h0000256c;  wr_data_rom[ 5651]='h00003ca8;
    rd_cycle[ 5652] = 1'b0;  wr_cycle[ 5652] = 1'b1;  addr_rom[ 5652]='h000014a4;  wr_data_rom[ 5652]='h00002f9e;
    rd_cycle[ 5653] = 1'b0;  wr_cycle[ 5653] = 1'b1;  addr_rom[ 5653]='h00000a20;  wr_data_rom[ 5653]='h000013b1;
    rd_cycle[ 5654] = 1'b0;  wr_cycle[ 5654] = 1'b1;  addr_rom[ 5654]='h00002c94;  wr_data_rom[ 5654]='h000030dc;
    rd_cycle[ 5655] = 1'b1;  wr_cycle[ 5655] = 1'b0;  addr_rom[ 5655]='h00001bec;  wr_data_rom[ 5655]='h00000000;
    rd_cycle[ 5656] = 1'b0;  wr_cycle[ 5656] = 1'b1;  addr_rom[ 5656]='h00000a20;  wr_data_rom[ 5656]='h000033ea;
    rd_cycle[ 5657] = 1'b1;  wr_cycle[ 5657] = 1'b0;  addr_rom[ 5657]='h00002b9c;  wr_data_rom[ 5657]='h00000000;
    rd_cycle[ 5658] = 1'b1;  wr_cycle[ 5658] = 1'b0;  addr_rom[ 5658]='h00003554;  wr_data_rom[ 5658]='h00000000;
    rd_cycle[ 5659] = 1'b1;  wr_cycle[ 5659] = 1'b0;  addr_rom[ 5659]='h00003b24;  wr_data_rom[ 5659]='h00000000;
    rd_cycle[ 5660] = 1'b1;  wr_cycle[ 5660] = 1'b0;  addr_rom[ 5660]='h00003f84;  wr_data_rom[ 5660]='h00000000;
    rd_cycle[ 5661] = 1'b1;  wr_cycle[ 5661] = 1'b0;  addr_rom[ 5661]='h00002664;  wr_data_rom[ 5661]='h00000000;
    rd_cycle[ 5662] = 1'b0;  wr_cycle[ 5662] = 1'b1;  addr_rom[ 5662]='h000015d4;  wr_data_rom[ 5662]='h00001aab;
    rd_cycle[ 5663] = 1'b0;  wr_cycle[ 5663] = 1'b1;  addr_rom[ 5663]='h00002f14;  wr_data_rom[ 5663]='h00000ef0;
    rd_cycle[ 5664] = 1'b1;  wr_cycle[ 5664] = 1'b0;  addr_rom[ 5664]='h00000884;  wr_data_rom[ 5664]='h00000000;
    rd_cycle[ 5665] = 1'b0;  wr_cycle[ 5665] = 1'b1;  addr_rom[ 5665]='h0000263c;  wr_data_rom[ 5665]='h00003ef1;
    rd_cycle[ 5666] = 1'b1;  wr_cycle[ 5666] = 1'b0;  addr_rom[ 5666]='h000030a0;  wr_data_rom[ 5666]='h00000000;
    rd_cycle[ 5667] = 1'b1;  wr_cycle[ 5667] = 1'b0;  addr_rom[ 5667]='h0000079c;  wr_data_rom[ 5667]='h00000000;
    rd_cycle[ 5668] = 1'b0;  wr_cycle[ 5668] = 1'b1;  addr_rom[ 5668]='h000013e0;  wr_data_rom[ 5668]='h00002683;
    rd_cycle[ 5669] = 1'b1;  wr_cycle[ 5669] = 1'b0;  addr_rom[ 5669]='h00001fa8;  wr_data_rom[ 5669]='h00000000;
    rd_cycle[ 5670] = 1'b0;  wr_cycle[ 5670] = 1'b1;  addr_rom[ 5670]='h000003e4;  wr_data_rom[ 5670]='h00002f70;
    rd_cycle[ 5671] = 1'b1;  wr_cycle[ 5671] = 1'b0;  addr_rom[ 5671]='h00003f68;  wr_data_rom[ 5671]='h00000000;
    rd_cycle[ 5672] = 1'b0;  wr_cycle[ 5672] = 1'b1;  addr_rom[ 5672]='h000015a4;  wr_data_rom[ 5672]='h00000a78;
    rd_cycle[ 5673] = 1'b1;  wr_cycle[ 5673] = 1'b0;  addr_rom[ 5673]='h00001dd8;  wr_data_rom[ 5673]='h00000000;
    rd_cycle[ 5674] = 1'b1;  wr_cycle[ 5674] = 1'b0;  addr_rom[ 5674]='h00000df0;  wr_data_rom[ 5674]='h00000000;
    rd_cycle[ 5675] = 1'b0;  wr_cycle[ 5675] = 1'b1;  addr_rom[ 5675]='h000035b8;  wr_data_rom[ 5675]='h000014c0;
    rd_cycle[ 5676] = 1'b1;  wr_cycle[ 5676] = 1'b0;  addr_rom[ 5676]='h000005e8;  wr_data_rom[ 5676]='h00000000;
    rd_cycle[ 5677] = 1'b0;  wr_cycle[ 5677] = 1'b1;  addr_rom[ 5677]='h000002dc;  wr_data_rom[ 5677]='h0000343a;
    rd_cycle[ 5678] = 1'b1;  wr_cycle[ 5678] = 1'b0;  addr_rom[ 5678]='h00003e6c;  wr_data_rom[ 5678]='h00000000;
    rd_cycle[ 5679] = 1'b0;  wr_cycle[ 5679] = 1'b1;  addr_rom[ 5679]='h00000a88;  wr_data_rom[ 5679]='h00000865;
    rd_cycle[ 5680] = 1'b1;  wr_cycle[ 5680] = 1'b0;  addr_rom[ 5680]='h00002040;  wr_data_rom[ 5680]='h00000000;
    rd_cycle[ 5681] = 1'b0;  wr_cycle[ 5681] = 1'b1;  addr_rom[ 5681]='h00001278;  wr_data_rom[ 5681]='h00000bf6;
    rd_cycle[ 5682] = 1'b0;  wr_cycle[ 5682] = 1'b1;  addr_rom[ 5682]='h00003ed8;  wr_data_rom[ 5682]='h00001319;
    rd_cycle[ 5683] = 1'b0;  wr_cycle[ 5683] = 1'b1;  addr_rom[ 5683]='h000025a8;  wr_data_rom[ 5683]='h00001328;
    rd_cycle[ 5684] = 1'b0;  wr_cycle[ 5684] = 1'b1;  addr_rom[ 5684]='h0000042c;  wr_data_rom[ 5684]='h00003810;
    rd_cycle[ 5685] = 1'b1;  wr_cycle[ 5685] = 1'b0;  addr_rom[ 5685]='h0000180c;  wr_data_rom[ 5685]='h00000000;
    rd_cycle[ 5686] = 1'b0;  wr_cycle[ 5686] = 1'b1;  addr_rom[ 5686]='h00000b9c;  wr_data_rom[ 5686]='h00000e68;
    rd_cycle[ 5687] = 1'b0;  wr_cycle[ 5687] = 1'b1;  addr_rom[ 5687]='h000029ac;  wr_data_rom[ 5687]='h00000e77;
    rd_cycle[ 5688] = 1'b0;  wr_cycle[ 5688] = 1'b1;  addr_rom[ 5688]='h00002118;  wr_data_rom[ 5688]='h00000a15;
    rd_cycle[ 5689] = 1'b0;  wr_cycle[ 5689] = 1'b1;  addr_rom[ 5689]='h000038fc;  wr_data_rom[ 5689]='h000015ee;
    rd_cycle[ 5690] = 1'b0;  wr_cycle[ 5690] = 1'b1;  addr_rom[ 5690]='h00001d9c;  wr_data_rom[ 5690]='h000013a2;
    rd_cycle[ 5691] = 1'b0;  wr_cycle[ 5691] = 1'b1;  addr_rom[ 5691]='h000032ac;  wr_data_rom[ 5691]='h000025ca;
    rd_cycle[ 5692] = 1'b1;  wr_cycle[ 5692] = 1'b0;  addr_rom[ 5692]='h00001b48;  wr_data_rom[ 5692]='h00000000;
    rd_cycle[ 5693] = 1'b0;  wr_cycle[ 5693] = 1'b1;  addr_rom[ 5693]='h00001274;  wr_data_rom[ 5693]='h00002c8d;
    rd_cycle[ 5694] = 1'b0;  wr_cycle[ 5694] = 1'b1;  addr_rom[ 5694]='h0000121c;  wr_data_rom[ 5694]='h00003aed;
    rd_cycle[ 5695] = 1'b0;  wr_cycle[ 5695] = 1'b1;  addr_rom[ 5695]='h00002260;  wr_data_rom[ 5695]='h00000eb6;
    rd_cycle[ 5696] = 1'b1;  wr_cycle[ 5696] = 1'b0;  addr_rom[ 5696]='h00003128;  wr_data_rom[ 5696]='h00000000;
    rd_cycle[ 5697] = 1'b0;  wr_cycle[ 5697] = 1'b1;  addr_rom[ 5697]='h000019ac;  wr_data_rom[ 5697]='h000017d8;
    rd_cycle[ 5698] = 1'b0;  wr_cycle[ 5698] = 1'b1;  addr_rom[ 5698]='h0000328c;  wr_data_rom[ 5698]='h00000370;
    rd_cycle[ 5699] = 1'b0;  wr_cycle[ 5699] = 1'b1;  addr_rom[ 5699]='h00003cbc;  wr_data_rom[ 5699]='h000029b3;
    rd_cycle[ 5700] = 1'b0;  wr_cycle[ 5700] = 1'b1;  addr_rom[ 5700]='h00000798;  wr_data_rom[ 5700]='h00003766;
    rd_cycle[ 5701] = 1'b1;  wr_cycle[ 5701] = 1'b0;  addr_rom[ 5701]='h0000218c;  wr_data_rom[ 5701]='h00000000;
    rd_cycle[ 5702] = 1'b1;  wr_cycle[ 5702] = 1'b0;  addr_rom[ 5702]='h00001b7c;  wr_data_rom[ 5702]='h00000000;
    rd_cycle[ 5703] = 1'b0;  wr_cycle[ 5703] = 1'b1;  addr_rom[ 5703]='h000007ac;  wr_data_rom[ 5703]='h00001b64;
    rd_cycle[ 5704] = 1'b1;  wr_cycle[ 5704] = 1'b0;  addr_rom[ 5704]='h00000948;  wr_data_rom[ 5704]='h00000000;
    rd_cycle[ 5705] = 1'b0;  wr_cycle[ 5705] = 1'b1;  addr_rom[ 5705]='h00001ae4;  wr_data_rom[ 5705]='h00002fb1;
    rd_cycle[ 5706] = 1'b1;  wr_cycle[ 5706] = 1'b0;  addr_rom[ 5706]='h00003e38;  wr_data_rom[ 5706]='h00000000;
    rd_cycle[ 5707] = 1'b0;  wr_cycle[ 5707] = 1'b1;  addr_rom[ 5707]='h00002e44;  wr_data_rom[ 5707]='h00002046;
    rd_cycle[ 5708] = 1'b1;  wr_cycle[ 5708] = 1'b0;  addr_rom[ 5708]='h00002f64;  wr_data_rom[ 5708]='h00000000;
    rd_cycle[ 5709] = 1'b0;  wr_cycle[ 5709] = 1'b1;  addr_rom[ 5709]='h000000a4;  wr_data_rom[ 5709]='h00002c7e;
    rd_cycle[ 5710] = 1'b1;  wr_cycle[ 5710] = 1'b0;  addr_rom[ 5710]='h00001b70;  wr_data_rom[ 5710]='h00000000;
    rd_cycle[ 5711] = 1'b1;  wr_cycle[ 5711] = 1'b0;  addr_rom[ 5711]='h000026ec;  wr_data_rom[ 5711]='h00000000;
    rd_cycle[ 5712] = 1'b1;  wr_cycle[ 5712] = 1'b0;  addr_rom[ 5712]='h000036a8;  wr_data_rom[ 5712]='h00000000;
    rd_cycle[ 5713] = 1'b0;  wr_cycle[ 5713] = 1'b1;  addr_rom[ 5713]='h000008c0;  wr_data_rom[ 5713]='h00001f2f;
    rd_cycle[ 5714] = 1'b0;  wr_cycle[ 5714] = 1'b1;  addr_rom[ 5714]='h0000014c;  wr_data_rom[ 5714]='h0000322a;
    rd_cycle[ 5715] = 1'b1;  wr_cycle[ 5715] = 1'b0;  addr_rom[ 5715]='h0000062c;  wr_data_rom[ 5715]='h00000000;
    rd_cycle[ 5716] = 1'b1;  wr_cycle[ 5716] = 1'b0;  addr_rom[ 5716]='h00002440;  wr_data_rom[ 5716]='h00000000;
    rd_cycle[ 5717] = 1'b0;  wr_cycle[ 5717] = 1'b1;  addr_rom[ 5717]='h000028e0;  wr_data_rom[ 5717]='h00001216;
    rd_cycle[ 5718] = 1'b1;  wr_cycle[ 5718] = 1'b0;  addr_rom[ 5718]='h000026e4;  wr_data_rom[ 5718]='h00000000;
    rd_cycle[ 5719] = 1'b0;  wr_cycle[ 5719] = 1'b1;  addr_rom[ 5719]='h0000183c;  wr_data_rom[ 5719]='h000022ec;
    rd_cycle[ 5720] = 1'b0;  wr_cycle[ 5720] = 1'b1;  addr_rom[ 5720]='h00003cb8;  wr_data_rom[ 5720]='h00002797;
    rd_cycle[ 5721] = 1'b1;  wr_cycle[ 5721] = 1'b0;  addr_rom[ 5721]='h000023cc;  wr_data_rom[ 5721]='h00000000;
    rd_cycle[ 5722] = 1'b1;  wr_cycle[ 5722] = 1'b0;  addr_rom[ 5722]='h00000ac4;  wr_data_rom[ 5722]='h00000000;
    rd_cycle[ 5723] = 1'b1;  wr_cycle[ 5723] = 1'b0;  addr_rom[ 5723]='h00003178;  wr_data_rom[ 5723]='h00000000;
    rd_cycle[ 5724] = 1'b0;  wr_cycle[ 5724] = 1'b1;  addr_rom[ 5724]='h00002b38;  wr_data_rom[ 5724]='h00001285;
    rd_cycle[ 5725] = 1'b0;  wr_cycle[ 5725] = 1'b1;  addr_rom[ 5725]='h00001ef8;  wr_data_rom[ 5725]='h0000136e;
    rd_cycle[ 5726] = 1'b0;  wr_cycle[ 5726] = 1'b1;  addr_rom[ 5726]='h00002114;  wr_data_rom[ 5726]='h0000366f;
    rd_cycle[ 5727] = 1'b0;  wr_cycle[ 5727] = 1'b1;  addr_rom[ 5727]='h00003360;  wr_data_rom[ 5727]='h000017f1;
    rd_cycle[ 5728] = 1'b1;  wr_cycle[ 5728] = 1'b0;  addr_rom[ 5728]='h00001f44;  wr_data_rom[ 5728]='h00000000;
    rd_cycle[ 5729] = 1'b1;  wr_cycle[ 5729] = 1'b0;  addr_rom[ 5729]='h00002d18;  wr_data_rom[ 5729]='h00000000;
    rd_cycle[ 5730] = 1'b0;  wr_cycle[ 5730] = 1'b1;  addr_rom[ 5730]='h00000824;  wr_data_rom[ 5730]='h0000190e;
    rd_cycle[ 5731] = 1'b0;  wr_cycle[ 5731] = 1'b1;  addr_rom[ 5731]='h00003368;  wr_data_rom[ 5731]='h00003e16;
    rd_cycle[ 5732] = 1'b1;  wr_cycle[ 5732] = 1'b0;  addr_rom[ 5732]='h00002088;  wr_data_rom[ 5732]='h00000000;
    rd_cycle[ 5733] = 1'b0;  wr_cycle[ 5733] = 1'b1;  addr_rom[ 5733]='h00003488;  wr_data_rom[ 5733]='h00001623;
    rd_cycle[ 5734] = 1'b1;  wr_cycle[ 5734] = 1'b0;  addr_rom[ 5734]='h00001728;  wr_data_rom[ 5734]='h00000000;
    rd_cycle[ 5735] = 1'b1;  wr_cycle[ 5735] = 1'b0;  addr_rom[ 5735]='h000025f0;  wr_data_rom[ 5735]='h00000000;
    rd_cycle[ 5736] = 1'b1;  wr_cycle[ 5736] = 1'b0;  addr_rom[ 5736]='h000008d0;  wr_data_rom[ 5736]='h00000000;
    rd_cycle[ 5737] = 1'b0;  wr_cycle[ 5737] = 1'b1;  addr_rom[ 5737]='h00002da8;  wr_data_rom[ 5737]='h00001732;
    rd_cycle[ 5738] = 1'b0;  wr_cycle[ 5738] = 1'b1;  addr_rom[ 5738]='h00002404;  wr_data_rom[ 5738]='h00002f94;
    rd_cycle[ 5739] = 1'b0;  wr_cycle[ 5739] = 1'b1;  addr_rom[ 5739]='h00002ab0;  wr_data_rom[ 5739]='h00001800;
    rd_cycle[ 5740] = 1'b0;  wr_cycle[ 5740] = 1'b1;  addr_rom[ 5740]='h00003690;  wr_data_rom[ 5740]='h000029bc;
    rd_cycle[ 5741] = 1'b0;  wr_cycle[ 5741] = 1'b1;  addr_rom[ 5741]='h00001c18;  wr_data_rom[ 5741]='h00002ea1;
    rd_cycle[ 5742] = 1'b1;  wr_cycle[ 5742] = 1'b0;  addr_rom[ 5742]='h00003850;  wr_data_rom[ 5742]='h00000000;
    rd_cycle[ 5743] = 1'b1;  wr_cycle[ 5743] = 1'b0;  addr_rom[ 5743]='h00003640;  wr_data_rom[ 5743]='h00000000;
    rd_cycle[ 5744] = 1'b0;  wr_cycle[ 5744] = 1'b1;  addr_rom[ 5744]='h00002f48;  wr_data_rom[ 5744]='h00003546;
    rd_cycle[ 5745] = 1'b1;  wr_cycle[ 5745] = 1'b0;  addr_rom[ 5745]='h00002134;  wr_data_rom[ 5745]='h00000000;
    rd_cycle[ 5746] = 1'b1;  wr_cycle[ 5746] = 1'b0;  addr_rom[ 5746]='h00000b5c;  wr_data_rom[ 5746]='h00000000;
    rd_cycle[ 5747] = 1'b0;  wr_cycle[ 5747] = 1'b1;  addr_rom[ 5747]='h000002ec;  wr_data_rom[ 5747]='h00003e39;
    rd_cycle[ 5748] = 1'b1;  wr_cycle[ 5748] = 1'b0;  addr_rom[ 5748]='h00003fb8;  wr_data_rom[ 5748]='h00000000;
    rd_cycle[ 5749] = 1'b1;  wr_cycle[ 5749] = 1'b0;  addr_rom[ 5749]='h00000d3c;  wr_data_rom[ 5749]='h00000000;
    rd_cycle[ 5750] = 1'b0;  wr_cycle[ 5750] = 1'b1;  addr_rom[ 5750]='h00000c58;  wr_data_rom[ 5750]='h0000199e;
    rd_cycle[ 5751] = 1'b0;  wr_cycle[ 5751] = 1'b1;  addr_rom[ 5751]='h000014cc;  wr_data_rom[ 5751]='h00003cb5;
    rd_cycle[ 5752] = 1'b1;  wr_cycle[ 5752] = 1'b0;  addr_rom[ 5752]='h00003ca4;  wr_data_rom[ 5752]='h00000000;
    rd_cycle[ 5753] = 1'b0;  wr_cycle[ 5753] = 1'b1;  addr_rom[ 5753]='h000039b8;  wr_data_rom[ 5753]='h000022d7;
    rd_cycle[ 5754] = 1'b0;  wr_cycle[ 5754] = 1'b1;  addr_rom[ 5754]='h00000ec0;  wr_data_rom[ 5754]='h00001000;
    rd_cycle[ 5755] = 1'b1;  wr_cycle[ 5755] = 1'b0;  addr_rom[ 5755]='h00003228;  wr_data_rom[ 5755]='h00000000;
    rd_cycle[ 5756] = 1'b0;  wr_cycle[ 5756] = 1'b1;  addr_rom[ 5756]='h00003840;  wr_data_rom[ 5756]='h000025cf;
    rd_cycle[ 5757] = 1'b0;  wr_cycle[ 5757] = 1'b1;  addr_rom[ 5757]='h000022bc;  wr_data_rom[ 5757]='h00000db3;
    rd_cycle[ 5758] = 1'b0;  wr_cycle[ 5758] = 1'b1;  addr_rom[ 5758]='h00002524;  wr_data_rom[ 5758]='h00003b20;
    rd_cycle[ 5759] = 1'b1;  wr_cycle[ 5759] = 1'b0;  addr_rom[ 5759]='h00001888;  wr_data_rom[ 5759]='h00000000;
    rd_cycle[ 5760] = 1'b1;  wr_cycle[ 5760] = 1'b0;  addr_rom[ 5760]='h000034dc;  wr_data_rom[ 5760]='h00000000;
    rd_cycle[ 5761] = 1'b0;  wr_cycle[ 5761] = 1'b1;  addr_rom[ 5761]='h000019ec;  wr_data_rom[ 5761]='h00001c06;
    rd_cycle[ 5762] = 1'b1;  wr_cycle[ 5762] = 1'b0;  addr_rom[ 5762]='h00002f4c;  wr_data_rom[ 5762]='h00000000;
    rd_cycle[ 5763] = 1'b1;  wr_cycle[ 5763] = 1'b0;  addr_rom[ 5763]='h00000f78;  wr_data_rom[ 5763]='h00000000;
    rd_cycle[ 5764] = 1'b0;  wr_cycle[ 5764] = 1'b1;  addr_rom[ 5764]='h00000d64;  wr_data_rom[ 5764]='h0000197c;
    rd_cycle[ 5765] = 1'b1;  wr_cycle[ 5765] = 1'b0;  addr_rom[ 5765]='h00000918;  wr_data_rom[ 5765]='h00000000;
    rd_cycle[ 5766] = 1'b0;  wr_cycle[ 5766] = 1'b1;  addr_rom[ 5766]='h00002e30;  wr_data_rom[ 5766]='h0000098d;
    rd_cycle[ 5767] = 1'b1;  wr_cycle[ 5767] = 1'b0;  addr_rom[ 5767]='h00002550;  wr_data_rom[ 5767]='h00000000;
    rd_cycle[ 5768] = 1'b0;  wr_cycle[ 5768] = 1'b1;  addr_rom[ 5768]='h0000359c;  wr_data_rom[ 5768]='h00003fb4;
    rd_cycle[ 5769] = 1'b1;  wr_cycle[ 5769] = 1'b0;  addr_rom[ 5769]='h000026b8;  wr_data_rom[ 5769]='h00000000;
    rd_cycle[ 5770] = 1'b1;  wr_cycle[ 5770] = 1'b0;  addr_rom[ 5770]='h000021e0;  wr_data_rom[ 5770]='h00000000;
    rd_cycle[ 5771] = 1'b1;  wr_cycle[ 5771] = 1'b0;  addr_rom[ 5771]='h00001690;  wr_data_rom[ 5771]='h00000000;
    rd_cycle[ 5772] = 1'b1;  wr_cycle[ 5772] = 1'b0;  addr_rom[ 5772]='h0000010c;  wr_data_rom[ 5772]='h00000000;
    rd_cycle[ 5773] = 1'b0;  wr_cycle[ 5773] = 1'b1;  addr_rom[ 5773]='h000031b8;  wr_data_rom[ 5773]='h000036a8;
    rd_cycle[ 5774] = 1'b1;  wr_cycle[ 5774] = 1'b0;  addr_rom[ 5774]='h00002518;  wr_data_rom[ 5774]='h00000000;
    rd_cycle[ 5775] = 1'b1;  wr_cycle[ 5775] = 1'b0;  addr_rom[ 5775]='h00003198;  wr_data_rom[ 5775]='h00000000;
    rd_cycle[ 5776] = 1'b0;  wr_cycle[ 5776] = 1'b1;  addr_rom[ 5776]='h0000003c;  wr_data_rom[ 5776]='h000005da;
    rd_cycle[ 5777] = 1'b1;  wr_cycle[ 5777] = 1'b0;  addr_rom[ 5777]='h000019ec;  wr_data_rom[ 5777]='h00000000;
    rd_cycle[ 5778] = 1'b1;  wr_cycle[ 5778] = 1'b0;  addr_rom[ 5778]='h0000004c;  wr_data_rom[ 5778]='h00000000;
    rd_cycle[ 5779] = 1'b1;  wr_cycle[ 5779] = 1'b0;  addr_rom[ 5779]='h000035a8;  wr_data_rom[ 5779]='h00000000;
    rd_cycle[ 5780] = 1'b0;  wr_cycle[ 5780] = 1'b1;  addr_rom[ 5780]='h00002c60;  wr_data_rom[ 5780]='h000032ca;
    rd_cycle[ 5781] = 1'b1;  wr_cycle[ 5781] = 1'b0;  addr_rom[ 5781]='h00002194;  wr_data_rom[ 5781]='h00000000;
    rd_cycle[ 5782] = 1'b1;  wr_cycle[ 5782] = 1'b0;  addr_rom[ 5782]='h00003df0;  wr_data_rom[ 5782]='h00000000;
    rd_cycle[ 5783] = 1'b0;  wr_cycle[ 5783] = 1'b1;  addr_rom[ 5783]='h00001288;  wr_data_rom[ 5783]='h00001035;
    rd_cycle[ 5784] = 1'b1;  wr_cycle[ 5784] = 1'b0;  addr_rom[ 5784]='h00000020;  wr_data_rom[ 5784]='h00000000;
    rd_cycle[ 5785] = 1'b1;  wr_cycle[ 5785] = 1'b0;  addr_rom[ 5785]='h00003840;  wr_data_rom[ 5785]='h00000000;
    rd_cycle[ 5786] = 1'b1;  wr_cycle[ 5786] = 1'b0;  addr_rom[ 5786]='h00000e74;  wr_data_rom[ 5786]='h00000000;
    rd_cycle[ 5787] = 1'b1;  wr_cycle[ 5787] = 1'b0;  addr_rom[ 5787]='h0000217c;  wr_data_rom[ 5787]='h00000000;
    rd_cycle[ 5788] = 1'b0;  wr_cycle[ 5788] = 1'b1;  addr_rom[ 5788]='h00000de0;  wr_data_rom[ 5788]='h00000315;
    rd_cycle[ 5789] = 1'b0;  wr_cycle[ 5789] = 1'b1;  addr_rom[ 5789]='h000016c0;  wr_data_rom[ 5789]='h00000ab6;
    rd_cycle[ 5790] = 1'b0;  wr_cycle[ 5790] = 1'b1;  addr_rom[ 5790]='h00003204;  wr_data_rom[ 5790]='h00001dd8;
    rd_cycle[ 5791] = 1'b0;  wr_cycle[ 5791] = 1'b1;  addr_rom[ 5791]='h0000285c;  wr_data_rom[ 5791]='h00000685;
    rd_cycle[ 5792] = 1'b0;  wr_cycle[ 5792] = 1'b1;  addr_rom[ 5792]='h0000221c;  wr_data_rom[ 5792]='h00000e4c;
    rd_cycle[ 5793] = 1'b0;  wr_cycle[ 5793] = 1'b1;  addr_rom[ 5793]='h00002a0c;  wr_data_rom[ 5793]='h00003bb0;
    rd_cycle[ 5794] = 1'b0;  wr_cycle[ 5794] = 1'b1;  addr_rom[ 5794]='h0000081c;  wr_data_rom[ 5794]='h00003ec7;
    rd_cycle[ 5795] = 1'b0;  wr_cycle[ 5795] = 1'b1;  addr_rom[ 5795]='h000025f8;  wr_data_rom[ 5795]='h00001762;
    rd_cycle[ 5796] = 1'b0;  wr_cycle[ 5796] = 1'b1;  addr_rom[ 5796]='h00001354;  wr_data_rom[ 5796]='h00000d37;
    rd_cycle[ 5797] = 1'b1;  wr_cycle[ 5797] = 1'b0;  addr_rom[ 5797]='h000032d4;  wr_data_rom[ 5797]='h00000000;
    rd_cycle[ 5798] = 1'b0;  wr_cycle[ 5798] = 1'b1;  addr_rom[ 5798]='h00000528;  wr_data_rom[ 5798]='h00002687;
    rd_cycle[ 5799] = 1'b0;  wr_cycle[ 5799] = 1'b1;  addr_rom[ 5799]='h000032e4;  wr_data_rom[ 5799]='h000035ed;
    rd_cycle[ 5800] = 1'b0;  wr_cycle[ 5800] = 1'b1;  addr_rom[ 5800]='h00003dc0;  wr_data_rom[ 5800]='h00001db0;
    rd_cycle[ 5801] = 1'b0;  wr_cycle[ 5801] = 1'b1;  addr_rom[ 5801]='h0000055c;  wr_data_rom[ 5801]='h00000dac;
    rd_cycle[ 5802] = 1'b0;  wr_cycle[ 5802] = 1'b1;  addr_rom[ 5802]='h0000141c;  wr_data_rom[ 5802]='h0000025f;
    rd_cycle[ 5803] = 1'b1;  wr_cycle[ 5803] = 1'b0;  addr_rom[ 5803]='h00000824;  wr_data_rom[ 5803]='h00000000;
    rd_cycle[ 5804] = 1'b0;  wr_cycle[ 5804] = 1'b1;  addr_rom[ 5804]='h000000b4;  wr_data_rom[ 5804]='h00001ade;
    rd_cycle[ 5805] = 1'b0;  wr_cycle[ 5805] = 1'b1;  addr_rom[ 5805]='h00001968;  wr_data_rom[ 5805]='h0000238c;
    rd_cycle[ 5806] = 1'b0;  wr_cycle[ 5806] = 1'b1;  addr_rom[ 5806]='h00000ddc;  wr_data_rom[ 5806]='h00001803;
    rd_cycle[ 5807] = 1'b0;  wr_cycle[ 5807] = 1'b1;  addr_rom[ 5807]='h000019f0;  wr_data_rom[ 5807]='h00003149;
    rd_cycle[ 5808] = 1'b1;  wr_cycle[ 5808] = 1'b0;  addr_rom[ 5808]='h000029e8;  wr_data_rom[ 5808]='h00000000;
    rd_cycle[ 5809] = 1'b1;  wr_cycle[ 5809] = 1'b0;  addr_rom[ 5809]='h00001178;  wr_data_rom[ 5809]='h00000000;
    rd_cycle[ 5810] = 1'b0;  wr_cycle[ 5810] = 1'b1;  addr_rom[ 5810]='h00001298;  wr_data_rom[ 5810]='h00003311;
    rd_cycle[ 5811] = 1'b1;  wr_cycle[ 5811] = 1'b0;  addr_rom[ 5811]='h00003e14;  wr_data_rom[ 5811]='h00000000;
    rd_cycle[ 5812] = 1'b1;  wr_cycle[ 5812] = 1'b0;  addr_rom[ 5812]='h00002e30;  wr_data_rom[ 5812]='h00000000;
    rd_cycle[ 5813] = 1'b0;  wr_cycle[ 5813] = 1'b1;  addr_rom[ 5813]='h000025ec;  wr_data_rom[ 5813]='h00003a9d;
    rd_cycle[ 5814] = 1'b0;  wr_cycle[ 5814] = 1'b1;  addr_rom[ 5814]='h0000007c;  wr_data_rom[ 5814]='h0000134e;
    rd_cycle[ 5815] = 1'b0;  wr_cycle[ 5815] = 1'b1;  addr_rom[ 5815]='h0000203c;  wr_data_rom[ 5815]='h00000f98;
    rd_cycle[ 5816] = 1'b0;  wr_cycle[ 5816] = 1'b1;  addr_rom[ 5816]='h00003d58;  wr_data_rom[ 5816]='h00002f12;
    rd_cycle[ 5817] = 1'b0;  wr_cycle[ 5817] = 1'b1;  addr_rom[ 5817]='h00002764;  wr_data_rom[ 5817]='h00003231;
    rd_cycle[ 5818] = 1'b1;  wr_cycle[ 5818] = 1'b0;  addr_rom[ 5818]='h000030d0;  wr_data_rom[ 5818]='h00000000;
    rd_cycle[ 5819] = 1'b1;  wr_cycle[ 5819] = 1'b0;  addr_rom[ 5819]='h00002898;  wr_data_rom[ 5819]='h00000000;
    rd_cycle[ 5820] = 1'b0;  wr_cycle[ 5820] = 1'b1;  addr_rom[ 5820]='h00002430;  wr_data_rom[ 5820]='h000004dd;
    rd_cycle[ 5821] = 1'b0;  wr_cycle[ 5821] = 1'b1;  addr_rom[ 5821]='h00003c44;  wr_data_rom[ 5821]='h00000d4a;
    rd_cycle[ 5822] = 1'b1;  wr_cycle[ 5822] = 1'b0;  addr_rom[ 5822]='h000035ac;  wr_data_rom[ 5822]='h00000000;
    rd_cycle[ 5823] = 1'b0;  wr_cycle[ 5823] = 1'b1;  addr_rom[ 5823]='h00003a38;  wr_data_rom[ 5823]='h000004e2;
    rd_cycle[ 5824] = 1'b0;  wr_cycle[ 5824] = 1'b1;  addr_rom[ 5824]='h0000133c;  wr_data_rom[ 5824]='h000020be;
    rd_cycle[ 5825] = 1'b0;  wr_cycle[ 5825] = 1'b1;  addr_rom[ 5825]='h00003f94;  wr_data_rom[ 5825]='h00002348;
    rd_cycle[ 5826] = 1'b1;  wr_cycle[ 5826] = 1'b0;  addr_rom[ 5826]='h000037e4;  wr_data_rom[ 5826]='h00000000;
    rd_cycle[ 5827] = 1'b1;  wr_cycle[ 5827] = 1'b0;  addr_rom[ 5827]='h000016f0;  wr_data_rom[ 5827]='h00000000;
    rd_cycle[ 5828] = 1'b0;  wr_cycle[ 5828] = 1'b1;  addr_rom[ 5828]='h00003c40;  wr_data_rom[ 5828]='h00001113;
    rd_cycle[ 5829] = 1'b1;  wr_cycle[ 5829] = 1'b0;  addr_rom[ 5829]='h00002bd8;  wr_data_rom[ 5829]='h00000000;
    rd_cycle[ 5830] = 1'b1;  wr_cycle[ 5830] = 1'b0;  addr_rom[ 5830]='h00002c88;  wr_data_rom[ 5830]='h00000000;
    rd_cycle[ 5831] = 1'b1;  wr_cycle[ 5831] = 1'b0;  addr_rom[ 5831]='h00000c08;  wr_data_rom[ 5831]='h00000000;
    rd_cycle[ 5832] = 1'b0;  wr_cycle[ 5832] = 1'b1;  addr_rom[ 5832]='h000001d8;  wr_data_rom[ 5832]='h00003862;
    rd_cycle[ 5833] = 1'b1;  wr_cycle[ 5833] = 1'b0;  addr_rom[ 5833]='h00000f64;  wr_data_rom[ 5833]='h00000000;
    rd_cycle[ 5834] = 1'b0;  wr_cycle[ 5834] = 1'b1;  addr_rom[ 5834]='h00000820;  wr_data_rom[ 5834]='h0000016a;
    rd_cycle[ 5835] = 1'b1;  wr_cycle[ 5835] = 1'b0;  addr_rom[ 5835]='h00001728;  wr_data_rom[ 5835]='h00000000;
    rd_cycle[ 5836] = 1'b1;  wr_cycle[ 5836] = 1'b0;  addr_rom[ 5836]='h00000ba0;  wr_data_rom[ 5836]='h00000000;
    rd_cycle[ 5837] = 1'b0;  wr_cycle[ 5837] = 1'b1;  addr_rom[ 5837]='h00000b3c;  wr_data_rom[ 5837]='h0000291f;
    rd_cycle[ 5838] = 1'b1;  wr_cycle[ 5838] = 1'b0;  addr_rom[ 5838]='h00003b04;  wr_data_rom[ 5838]='h00000000;
    rd_cycle[ 5839] = 1'b1;  wr_cycle[ 5839] = 1'b0;  addr_rom[ 5839]='h0000281c;  wr_data_rom[ 5839]='h00000000;
    rd_cycle[ 5840] = 1'b1;  wr_cycle[ 5840] = 1'b0;  addr_rom[ 5840]='h0000023c;  wr_data_rom[ 5840]='h00000000;
    rd_cycle[ 5841] = 1'b1;  wr_cycle[ 5841] = 1'b0;  addr_rom[ 5841]='h00003280;  wr_data_rom[ 5841]='h00000000;
    rd_cycle[ 5842] = 1'b0;  wr_cycle[ 5842] = 1'b1;  addr_rom[ 5842]='h00000068;  wr_data_rom[ 5842]='h000021b9;
    rd_cycle[ 5843] = 1'b1;  wr_cycle[ 5843] = 1'b0;  addr_rom[ 5843]='h000021b8;  wr_data_rom[ 5843]='h00000000;
    rd_cycle[ 5844] = 1'b1;  wr_cycle[ 5844] = 1'b0;  addr_rom[ 5844]='h00002054;  wr_data_rom[ 5844]='h00000000;
    rd_cycle[ 5845] = 1'b0;  wr_cycle[ 5845] = 1'b1;  addr_rom[ 5845]='h00000760;  wr_data_rom[ 5845]='h00001c44;
    rd_cycle[ 5846] = 1'b1;  wr_cycle[ 5846] = 1'b0;  addr_rom[ 5846]='h00003bf4;  wr_data_rom[ 5846]='h00000000;
    rd_cycle[ 5847] = 1'b0;  wr_cycle[ 5847] = 1'b1;  addr_rom[ 5847]='h0000299c;  wr_data_rom[ 5847]='h00002cb0;
    rd_cycle[ 5848] = 1'b1;  wr_cycle[ 5848] = 1'b0;  addr_rom[ 5848]='h00001ab8;  wr_data_rom[ 5848]='h00000000;
    rd_cycle[ 5849] = 1'b0;  wr_cycle[ 5849] = 1'b1;  addr_rom[ 5849]='h000030a0;  wr_data_rom[ 5849]='h00003205;
    rd_cycle[ 5850] = 1'b1;  wr_cycle[ 5850] = 1'b0;  addr_rom[ 5850]='h00001390;  wr_data_rom[ 5850]='h00000000;
    rd_cycle[ 5851] = 1'b0;  wr_cycle[ 5851] = 1'b1;  addr_rom[ 5851]='h000016f4;  wr_data_rom[ 5851]='h0000244e;
    rd_cycle[ 5852] = 1'b1;  wr_cycle[ 5852] = 1'b0;  addr_rom[ 5852]='h0000062c;  wr_data_rom[ 5852]='h00000000;
    rd_cycle[ 5853] = 1'b0;  wr_cycle[ 5853] = 1'b1;  addr_rom[ 5853]='h000024f4;  wr_data_rom[ 5853]='h000039cd;
    rd_cycle[ 5854] = 1'b0;  wr_cycle[ 5854] = 1'b1;  addr_rom[ 5854]='h00001dd8;  wr_data_rom[ 5854]='h00001a43;
    rd_cycle[ 5855] = 1'b0;  wr_cycle[ 5855] = 1'b1;  addr_rom[ 5855]='h00003d98;  wr_data_rom[ 5855]='h000036c1;
    rd_cycle[ 5856] = 1'b0;  wr_cycle[ 5856] = 1'b1;  addr_rom[ 5856]='h00001300;  wr_data_rom[ 5856]='h00002196;
    rd_cycle[ 5857] = 1'b0;  wr_cycle[ 5857] = 1'b1;  addr_rom[ 5857]='h00001b70;  wr_data_rom[ 5857]='h000000ad;
    rd_cycle[ 5858] = 1'b1;  wr_cycle[ 5858] = 1'b0;  addr_rom[ 5858]='h00001d74;  wr_data_rom[ 5858]='h00000000;
    rd_cycle[ 5859] = 1'b1;  wr_cycle[ 5859] = 1'b0;  addr_rom[ 5859]='h00003910;  wr_data_rom[ 5859]='h00000000;
    rd_cycle[ 5860] = 1'b0;  wr_cycle[ 5860] = 1'b1;  addr_rom[ 5860]='h00003d14;  wr_data_rom[ 5860]='h00000ddb;
    rd_cycle[ 5861] = 1'b1;  wr_cycle[ 5861] = 1'b0;  addr_rom[ 5861]='h000023e0;  wr_data_rom[ 5861]='h00000000;
    rd_cycle[ 5862] = 1'b1;  wr_cycle[ 5862] = 1'b0;  addr_rom[ 5862]='h00002e5c;  wr_data_rom[ 5862]='h00000000;
    rd_cycle[ 5863] = 1'b0;  wr_cycle[ 5863] = 1'b1;  addr_rom[ 5863]='h00003108;  wr_data_rom[ 5863]='h00003754;
    rd_cycle[ 5864] = 1'b0;  wr_cycle[ 5864] = 1'b1;  addr_rom[ 5864]='h0000041c;  wr_data_rom[ 5864]='h00003cbe;
    rd_cycle[ 5865] = 1'b0;  wr_cycle[ 5865] = 1'b1;  addr_rom[ 5865]='h00002ef0;  wr_data_rom[ 5865]='h00001a13;
    rd_cycle[ 5866] = 1'b1;  wr_cycle[ 5866] = 1'b0;  addr_rom[ 5866]='h000025d0;  wr_data_rom[ 5866]='h00000000;
    rd_cycle[ 5867] = 1'b1;  wr_cycle[ 5867] = 1'b0;  addr_rom[ 5867]='h00001c84;  wr_data_rom[ 5867]='h00000000;
    rd_cycle[ 5868] = 1'b1;  wr_cycle[ 5868] = 1'b0;  addr_rom[ 5868]='h00000cf0;  wr_data_rom[ 5868]='h00000000;
    rd_cycle[ 5869] = 1'b0;  wr_cycle[ 5869] = 1'b1;  addr_rom[ 5869]='h00001748;  wr_data_rom[ 5869]='h00002657;
    rd_cycle[ 5870] = 1'b0;  wr_cycle[ 5870] = 1'b1;  addr_rom[ 5870]='h000033b4;  wr_data_rom[ 5870]='h00003231;
    rd_cycle[ 5871] = 1'b0;  wr_cycle[ 5871] = 1'b1;  addr_rom[ 5871]='h00000a64;  wr_data_rom[ 5871]='h00001dcb;
    rd_cycle[ 5872] = 1'b1;  wr_cycle[ 5872] = 1'b0;  addr_rom[ 5872]='h0000213c;  wr_data_rom[ 5872]='h00000000;
    rd_cycle[ 5873] = 1'b1;  wr_cycle[ 5873] = 1'b0;  addr_rom[ 5873]='h00003e14;  wr_data_rom[ 5873]='h00000000;
    rd_cycle[ 5874] = 1'b1;  wr_cycle[ 5874] = 1'b0;  addr_rom[ 5874]='h000030c0;  wr_data_rom[ 5874]='h00000000;
    rd_cycle[ 5875] = 1'b1;  wr_cycle[ 5875] = 1'b0;  addr_rom[ 5875]='h00001628;  wr_data_rom[ 5875]='h00000000;
    rd_cycle[ 5876] = 1'b1;  wr_cycle[ 5876] = 1'b0;  addr_rom[ 5876]='h000006e0;  wr_data_rom[ 5876]='h00000000;
    rd_cycle[ 5877] = 1'b0;  wr_cycle[ 5877] = 1'b1;  addr_rom[ 5877]='h00000304;  wr_data_rom[ 5877]='h00000a18;
    rd_cycle[ 5878] = 1'b1;  wr_cycle[ 5878] = 1'b0;  addr_rom[ 5878]='h00002a60;  wr_data_rom[ 5878]='h00000000;
    rd_cycle[ 5879] = 1'b1;  wr_cycle[ 5879] = 1'b0;  addr_rom[ 5879]='h00001d08;  wr_data_rom[ 5879]='h00000000;
    rd_cycle[ 5880] = 1'b1;  wr_cycle[ 5880] = 1'b0;  addr_rom[ 5880]='h000026cc;  wr_data_rom[ 5880]='h00000000;
    rd_cycle[ 5881] = 1'b0;  wr_cycle[ 5881] = 1'b1;  addr_rom[ 5881]='h00002808;  wr_data_rom[ 5881]='h000012fd;
    rd_cycle[ 5882] = 1'b1;  wr_cycle[ 5882] = 1'b0;  addr_rom[ 5882]='h00000730;  wr_data_rom[ 5882]='h00000000;
    rd_cycle[ 5883] = 1'b1;  wr_cycle[ 5883] = 1'b0;  addr_rom[ 5883]='h000013b4;  wr_data_rom[ 5883]='h00000000;
    rd_cycle[ 5884] = 1'b1;  wr_cycle[ 5884] = 1'b0;  addr_rom[ 5884]='h000039a8;  wr_data_rom[ 5884]='h00000000;
    rd_cycle[ 5885] = 1'b1;  wr_cycle[ 5885] = 1'b0;  addr_rom[ 5885]='h000026f4;  wr_data_rom[ 5885]='h00000000;
    rd_cycle[ 5886] = 1'b1;  wr_cycle[ 5886] = 1'b0;  addr_rom[ 5886]='h0000310c;  wr_data_rom[ 5886]='h00000000;
    rd_cycle[ 5887] = 1'b1;  wr_cycle[ 5887] = 1'b0;  addr_rom[ 5887]='h00003804;  wr_data_rom[ 5887]='h00000000;
    rd_cycle[ 5888] = 1'b1;  wr_cycle[ 5888] = 1'b0;  addr_rom[ 5888]='h00000f38;  wr_data_rom[ 5888]='h00000000;
    rd_cycle[ 5889] = 1'b0;  wr_cycle[ 5889] = 1'b1;  addr_rom[ 5889]='h00000644;  wr_data_rom[ 5889]='h00003fa8;
    rd_cycle[ 5890] = 1'b0;  wr_cycle[ 5890] = 1'b1;  addr_rom[ 5890]='h00002aa4;  wr_data_rom[ 5890]='h00003a86;
    rd_cycle[ 5891] = 1'b1;  wr_cycle[ 5891] = 1'b0;  addr_rom[ 5891]='h00001670;  wr_data_rom[ 5891]='h00000000;
    rd_cycle[ 5892] = 1'b1;  wr_cycle[ 5892] = 1'b0;  addr_rom[ 5892]='h00001038;  wr_data_rom[ 5892]='h00000000;
    rd_cycle[ 5893] = 1'b0;  wr_cycle[ 5893] = 1'b1;  addr_rom[ 5893]='h000029f8;  wr_data_rom[ 5893]='h000030fa;
    rd_cycle[ 5894] = 1'b1;  wr_cycle[ 5894] = 1'b0;  addr_rom[ 5894]='h00001004;  wr_data_rom[ 5894]='h00000000;
    rd_cycle[ 5895] = 1'b1;  wr_cycle[ 5895] = 1'b0;  addr_rom[ 5895]='h0000077c;  wr_data_rom[ 5895]='h00000000;
    rd_cycle[ 5896] = 1'b0;  wr_cycle[ 5896] = 1'b1;  addr_rom[ 5896]='h00003fcc;  wr_data_rom[ 5896]='h0000163a;
    rd_cycle[ 5897] = 1'b1;  wr_cycle[ 5897] = 1'b0;  addr_rom[ 5897]='h000018d8;  wr_data_rom[ 5897]='h00000000;
    rd_cycle[ 5898] = 1'b0;  wr_cycle[ 5898] = 1'b1;  addr_rom[ 5898]='h000020e4;  wr_data_rom[ 5898]='h0000305f;
    rd_cycle[ 5899] = 1'b1;  wr_cycle[ 5899] = 1'b0;  addr_rom[ 5899]='h00003658;  wr_data_rom[ 5899]='h00000000;
    rd_cycle[ 5900] = 1'b1;  wr_cycle[ 5900] = 1'b0;  addr_rom[ 5900]='h000024cc;  wr_data_rom[ 5900]='h00000000;
    rd_cycle[ 5901] = 1'b1;  wr_cycle[ 5901] = 1'b0;  addr_rom[ 5901]='h00001c80;  wr_data_rom[ 5901]='h00000000;
    rd_cycle[ 5902] = 1'b0;  wr_cycle[ 5902] = 1'b1;  addr_rom[ 5902]='h00002768;  wr_data_rom[ 5902]='h00003667;
    rd_cycle[ 5903] = 1'b0;  wr_cycle[ 5903] = 1'b1;  addr_rom[ 5903]='h00003598;  wr_data_rom[ 5903]='h00000179;
    rd_cycle[ 5904] = 1'b0;  wr_cycle[ 5904] = 1'b1;  addr_rom[ 5904]='h00002f54;  wr_data_rom[ 5904]='h00003531;
    rd_cycle[ 5905] = 1'b0;  wr_cycle[ 5905] = 1'b1;  addr_rom[ 5905]='h00001834;  wr_data_rom[ 5905]='h000004b5;
    rd_cycle[ 5906] = 1'b0;  wr_cycle[ 5906] = 1'b1;  addr_rom[ 5906]='h00000288;  wr_data_rom[ 5906]='h00000c7b;
    rd_cycle[ 5907] = 1'b0;  wr_cycle[ 5907] = 1'b1;  addr_rom[ 5907]='h00001a48;  wr_data_rom[ 5907]='h000014d9;
    rd_cycle[ 5908] = 1'b1;  wr_cycle[ 5908] = 1'b0;  addr_rom[ 5908]='h00003fc0;  wr_data_rom[ 5908]='h00000000;
    rd_cycle[ 5909] = 1'b0;  wr_cycle[ 5909] = 1'b1;  addr_rom[ 5909]='h00003968;  wr_data_rom[ 5909]='h00003a7f;
    rd_cycle[ 5910] = 1'b0;  wr_cycle[ 5910] = 1'b1;  addr_rom[ 5910]='h000005c0;  wr_data_rom[ 5910]='h0000365c;
    rd_cycle[ 5911] = 1'b1;  wr_cycle[ 5911] = 1'b0;  addr_rom[ 5911]='h0000370c;  wr_data_rom[ 5911]='h00000000;
    rd_cycle[ 5912] = 1'b0;  wr_cycle[ 5912] = 1'b1;  addr_rom[ 5912]='h000032c4;  wr_data_rom[ 5912]='h00000940;
    rd_cycle[ 5913] = 1'b0;  wr_cycle[ 5913] = 1'b1;  addr_rom[ 5913]='h000002c8;  wr_data_rom[ 5913]='h00000d78;
    rd_cycle[ 5914] = 1'b1;  wr_cycle[ 5914] = 1'b0;  addr_rom[ 5914]='h00003f74;  wr_data_rom[ 5914]='h00000000;
    rd_cycle[ 5915] = 1'b1;  wr_cycle[ 5915] = 1'b0;  addr_rom[ 5915]='h00002f18;  wr_data_rom[ 5915]='h00000000;
    rd_cycle[ 5916] = 1'b0;  wr_cycle[ 5916] = 1'b1;  addr_rom[ 5916]='h00000408;  wr_data_rom[ 5916]='h00000ce5;
    rd_cycle[ 5917] = 1'b0;  wr_cycle[ 5917] = 1'b1;  addr_rom[ 5917]='h0000145c;  wr_data_rom[ 5917]='h000022ee;
    rd_cycle[ 5918] = 1'b0;  wr_cycle[ 5918] = 1'b1;  addr_rom[ 5918]='h00000200;  wr_data_rom[ 5918]='h00003288;
    rd_cycle[ 5919] = 1'b0;  wr_cycle[ 5919] = 1'b1;  addr_rom[ 5919]='h00002a38;  wr_data_rom[ 5919]='h00000a6c;
    rd_cycle[ 5920] = 1'b1;  wr_cycle[ 5920] = 1'b0;  addr_rom[ 5920]='h00002224;  wr_data_rom[ 5920]='h00000000;
    rd_cycle[ 5921] = 1'b1;  wr_cycle[ 5921] = 1'b0;  addr_rom[ 5921]='h00000254;  wr_data_rom[ 5921]='h00000000;
    rd_cycle[ 5922] = 1'b0;  wr_cycle[ 5922] = 1'b1;  addr_rom[ 5922]='h000039ec;  wr_data_rom[ 5922]='h00002857;
    rd_cycle[ 5923] = 1'b0;  wr_cycle[ 5923] = 1'b1;  addr_rom[ 5923]='h00003d80;  wr_data_rom[ 5923]='h000017e2;
    rd_cycle[ 5924] = 1'b1;  wr_cycle[ 5924] = 1'b0;  addr_rom[ 5924]='h00001b98;  wr_data_rom[ 5924]='h00000000;
    rd_cycle[ 5925] = 1'b1;  wr_cycle[ 5925] = 1'b0;  addr_rom[ 5925]='h00001d70;  wr_data_rom[ 5925]='h00000000;
    rd_cycle[ 5926] = 1'b0;  wr_cycle[ 5926] = 1'b1;  addr_rom[ 5926]='h000021e8;  wr_data_rom[ 5926]='h000000a7;
    rd_cycle[ 5927] = 1'b1;  wr_cycle[ 5927] = 1'b0;  addr_rom[ 5927]='h00003920;  wr_data_rom[ 5927]='h00000000;
    rd_cycle[ 5928] = 1'b1;  wr_cycle[ 5928] = 1'b0;  addr_rom[ 5928]='h00001914;  wr_data_rom[ 5928]='h00000000;
    rd_cycle[ 5929] = 1'b1;  wr_cycle[ 5929] = 1'b0;  addr_rom[ 5929]='h00001ad4;  wr_data_rom[ 5929]='h00000000;
    rd_cycle[ 5930] = 1'b1;  wr_cycle[ 5930] = 1'b0;  addr_rom[ 5930]='h00003fbc;  wr_data_rom[ 5930]='h00000000;
    rd_cycle[ 5931] = 1'b1;  wr_cycle[ 5931] = 1'b0;  addr_rom[ 5931]='h0000215c;  wr_data_rom[ 5931]='h00000000;
    rd_cycle[ 5932] = 1'b1;  wr_cycle[ 5932] = 1'b0;  addr_rom[ 5932]='h00003028;  wr_data_rom[ 5932]='h00000000;
    rd_cycle[ 5933] = 1'b1;  wr_cycle[ 5933] = 1'b0;  addr_rom[ 5933]='h00002b80;  wr_data_rom[ 5933]='h00000000;
    rd_cycle[ 5934] = 1'b0;  wr_cycle[ 5934] = 1'b1;  addr_rom[ 5934]='h0000034c;  wr_data_rom[ 5934]='h00002cb4;
    rd_cycle[ 5935] = 1'b1;  wr_cycle[ 5935] = 1'b0;  addr_rom[ 5935]='h00000ad8;  wr_data_rom[ 5935]='h00000000;
    rd_cycle[ 5936] = 1'b1;  wr_cycle[ 5936] = 1'b0;  addr_rom[ 5936]='h00003de4;  wr_data_rom[ 5936]='h00000000;
    rd_cycle[ 5937] = 1'b1;  wr_cycle[ 5937] = 1'b0;  addr_rom[ 5937]='h00002d40;  wr_data_rom[ 5937]='h00000000;
    rd_cycle[ 5938] = 1'b1;  wr_cycle[ 5938] = 1'b0;  addr_rom[ 5938]='h00003594;  wr_data_rom[ 5938]='h00000000;
    rd_cycle[ 5939] = 1'b1;  wr_cycle[ 5939] = 1'b0;  addr_rom[ 5939]='h0000300c;  wr_data_rom[ 5939]='h00000000;
    rd_cycle[ 5940] = 1'b0;  wr_cycle[ 5940] = 1'b1;  addr_rom[ 5940]='h00002b78;  wr_data_rom[ 5940]='h00002f2c;
    rd_cycle[ 5941] = 1'b0;  wr_cycle[ 5941] = 1'b1;  addr_rom[ 5941]='h00001668;  wr_data_rom[ 5941]='h0000012a;
    rd_cycle[ 5942] = 1'b1;  wr_cycle[ 5942] = 1'b0;  addr_rom[ 5942]='h00003b48;  wr_data_rom[ 5942]='h00000000;
    rd_cycle[ 5943] = 1'b1;  wr_cycle[ 5943] = 1'b0;  addr_rom[ 5943]='h00003e44;  wr_data_rom[ 5943]='h00000000;
    rd_cycle[ 5944] = 1'b0;  wr_cycle[ 5944] = 1'b1;  addr_rom[ 5944]='h0000231c;  wr_data_rom[ 5944]='h00000af7;
    rd_cycle[ 5945] = 1'b1;  wr_cycle[ 5945] = 1'b0;  addr_rom[ 5945]='h000034a0;  wr_data_rom[ 5945]='h00000000;
    rd_cycle[ 5946] = 1'b1;  wr_cycle[ 5946] = 1'b0;  addr_rom[ 5946]='h00003090;  wr_data_rom[ 5946]='h00000000;
    rd_cycle[ 5947] = 1'b0;  wr_cycle[ 5947] = 1'b1;  addr_rom[ 5947]='h00003834;  wr_data_rom[ 5947]='h000029ae;
    rd_cycle[ 5948] = 1'b1;  wr_cycle[ 5948] = 1'b0;  addr_rom[ 5948]='h000008a0;  wr_data_rom[ 5948]='h00000000;
    rd_cycle[ 5949] = 1'b0;  wr_cycle[ 5949] = 1'b1;  addr_rom[ 5949]='h00003a7c;  wr_data_rom[ 5949]='h00002811;
    rd_cycle[ 5950] = 1'b0;  wr_cycle[ 5950] = 1'b1;  addr_rom[ 5950]='h000035fc;  wr_data_rom[ 5950]='h00002f34;
    rd_cycle[ 5951] = 1'b0;  wr_cycle[ 5951] = 1'b1;  addr_rom[ 5951]='h000038e0;  wr_data_rom[ 5951]='h00000ad9;
    rd_cycle[ 5952] = 1'b1;  wr_cycle[ 5952] = 1'b0;  addr_rom[ 5952]='h00003ef8;  wr_data_rom[ 5952]='h00000000;
    rd_cycle[ 5953] = 1'b1;  wr_cycle[ 5953] = 1'b0;  addr_rom[ 5953]='h0000232c;  wr_data_rom[ 5953]='h00000000;
    rd_cycle[ 5954] = 1'b0;  wr_cycle[ 5954] = 1'b1;  addr_rom[ 5954]='h0000134c;  wr_data_rom[ 5954]='h0000077a;
    rd_cycle[ 5955] = 1'b0;  wr_cycle[ 5955] = 1'b1;  addr_rom[ 5955]='h00003e84;  wr_data_rom[ 5955]='h00003c7e;
    rd_cycle[ 5956] = 1'b0;  wr_cycle[ 5956] = 1'b1;  addr_rom[ 5956]='h000031e4;  wr_data_rom[ 5956]='h000021d1;
    rd_cycle[ 5957] = 1'b1;  wr_cycle[ 5957] = 1'b0;  addr_rom[ 5957]='h00002df0;  wr_data_rom[ 5957]='h00000000;
    rd_cycle[ 5958] = 1'b1;  wr_cycle[ 5958] = 1'b0;  addr_rom[ 5958]='h00001284;  wr_data_rom[ 5958]='h00000000;
    rd_cycle[ 5959] = 1'b1;  wr_cycle[ 5959] = 1'b0;  addr_rom[ 5959]='h00000c50;  wr_data_rom[ 5959]='h00000000;
    rd_cycle[ 5960] = 1'b1;  wr_cycle[ 5960] = 1'b0;  addr_rom[ 5960]='h00003160;  wr_data_rom[ 5960]='h00000000;
    rd_cycle[ 5961] = 1'b0;  wr_cycle[ 5961] = 1'b1;  addr_rom[ 5961]='h000005b0;  wr_data_rom[ 5961]='h00000481;
    rd_cycle[ 5962] = 1'b0;  wr_cycle[ 5962] = 1'b1;  addr_rom[ 5962]='h000005e8;  wr_data_rom[ 5962]='h000009f1;
    rd_cycle[ 5963] = 1'b0;  wr_cycle[ 5963] = 1'b1;  addr_rom[ 5963]='h00001c40;  wr_data_rom[ 5963]='h000030dd;
    rd_cycle[ 5964] = 1'b0;  wr_cycle[ 5964] = 1'b1;  addr_rom[ 5964]='h00001444;  wr_data_rom[ 5964]='h000000ca;
    rd_cycle[ 5965] = 1'b1;  wr_cycle[ 5965] = 1'b0;  addr_rom[ 5965]='h00003370;  wr_data_rom[ 5965]='h00000000;
    rd_cycle[ 5966] = 1'b0;  wr_cycle[ 5966] = 1'b1;  addr_rom[ 5966]='h0000188c;  wr_data_rom[ 5966]='h00002f16;
    rd_cycle[ 5967] = 1'b0;  wr_cycle[ 5967] = 1'b1;  addr_rom[ 5967]='h00000870;  wr_data_rom[ 5967]='h000033ae;
    rd_cycle[ 5968] = 1'b0;  wr_cycle[ 5968] = 1'b1;  addr_rom[ 5968]='h000023ac;  wr_data_rom[ 5968]='h00003b4f;
    rd_cycle[ 5969] = 1'b0;  wr_cycle[ 5969] = 1'b1;  addr_rom[ 5969]='h00002a5c;  wr_data_rom[ 5969]='h00001621;
    rd_cycle[ 5970] = 1'b1;  wr_cycle[ 5970] = 1'b0;  addr_rom[ 5970]='h0000193c;  wr_data_rom[ 5970]='h00000000;
    rd_cycle[ 5971] = 1'b1;  wr_cycle[ 5971] = 1'b0;  addr_rom[ 5971]='h00000814;  wr_data_rom[ 5971]='h00000000;
    rd_cycle[ 5972] = 1'b1;  wr_cycle[ 5972] = 1'b0;  addr_rom[ 5972]='h00002074;  wr_data_rom[ 5972]='h00000000;
    rd_cycle[ 5973] = 1'b1;  wr_cycle[ 5973] = 1'b0;  addr_rom[ 5973]='h000034b8;  wr_data_rom[ 5973]='h00000000;
    rd_cycle[ 5974] = 1'b0;  wr_cycle[ 5974] = 1'b1;  addr_rom[ 5974]='h00000868;  wr_data_rom[ 5974]='h0000244f;
    rd_cycle[ 5975] = 1'b0;  wr_cycle[ 5975] = 1'b1;  addr_rom[ 5975]='h00002e00;  wr_data_rom[ 5975]='h00000064;
    rd_cycle[ 5976] = 1'b1;  wr_cycle[ 5976] = 1'b0;  addr_rom[ 5976]='h00003be4;  wr_data_rom[ 5976]='h00000000;
    rd_cycle[ 5977] = 1'b0;  wr_cycle[ 5977] = 1'b1;  addr_rom[ 5977]='h0000188c;  wr_data_rom[ 5977]='h000029d1;
    rd_cycle[ 5978] = 1'b1;  wr_cycle[ 5978] = 1'b0;  addr_rom[ 5978]='h00001068;  wr_data_rom[ 5978]='h00000000;
    rd_cycle[ 5979] = 1'b0;  wr_cycle[ 5979] = 1'b1;  addr_rom[ 5979]='h00002b24;  wr_data_rom[ 5979]='h00001646;
    rd_cycle[ 5980] = 1'b1;  wr_cycle[ 5980] = 1'b0;  addr_rom[ 5980]='h00001bcc;  wr_data_rom[ 5980]='h00000000;
    rd_cycle[ 5981] = 1'b1;  wr_cycle[ 5981] = 1'b0;  addr_rom[ 5981]='h00001bb0;  wr_data_rom[ 5981]='h00000000;
    rd_cycle[ 5982] = 1'b1;  wr_cycle[ 5982] = 1'b0;  addr_rom[ 5982]='h00002d58;  wr_data_rom[ 5982]='h00000000;
    rd_cycle[ 5983] = 1'b1;  wr_cycle[ 5983] = 1'b0;  addr_rom[ 5983]='h00000e08;  wr_data_rom[ 5983]='h00000000;
    rd_cycle[ 5984] = 1'b0;  wr_cycle[ 5984] = 1'b1;  addr_rom[ 5984]='h000004b0;  wr_data_rom[ 5984]='h00001a83;
    rd_cycle[ 5985] = 1'b1;  wr_cycle[ 5985] = 1'b0;  addr_rom[ 5985]='h00000bbc;  wr_data_rom[ 5985]='h00000000;
    rd_cycle[ 5986] = 1'b0;  wr_cycle[ 5986] = 1'b1;  addr_rom[ 5986]='h00000aa8;  wr_data_rom[ 5986]='h00003d5e;
    rd_cycle[ 5987] = 1'b1;  wr_cycle[ 5987] = 1'b0;  addr_rom[ 5987]='h00001b28;  wr_data_rom[ 5987]='h00000000;
    rd_cycle[ 5988] = 1'b1;  wr_cycle[ 5988] = 1'b0;  addr_rom[ 5988]='h000019c0;  wr_data_rom[ 5988]='h00000000;
    rd_cycle[ 5989] = 1'b1;  wr_cycle[ 5989] = 1'b0;  addr_rom[ 5989]='h000028f4;  wr_data_rom[ 5989]='h00000000;
    rd_cycle[ 5990] = 1'b0;  wr_cycle[ 5990] = 1'b1;  addr_rom[ 5990]='h00001218;  wr_data_rom[ 5990]='h000014eb;
    rd_cycle[ 5991] = 1'b1;  wr_cycle[ 5991] = 1'b0;  addr_rom[ 5991]='h00003040;  wr_data_rom[ 5991]='h00000000;
    rd_cycle[ 5992] = 1'b1;  wr_cycle[ 5992] = 1'b0;  addr_rom[ 5992]='h00003ca0;  wr_data_rom[ 5992]='h00000000;
    rd_cycle[ 5993] = 1'b1;  wr_cycle[ 5993] = 1'b0;  addr_rom[ 5993]='h00000cf4;  wr_data_rom[ 5993]='h00000000;
    rd_cycle[ 5994] = 1'b0;  wr_cycle[ 5994] = 1'b1;  addr_rom[ 5994]='h00003470;  wr_data_rom[ 5994]='h00003bbc;
    rd_cycle[ 5995] = 1'b1;  wr_cycle[ 5995] = 1'b0;  addr_rom[ 5995]='h000006f4;  wr_data_rom[ 5995]='h00000000;
    rd_cycle[ 5996] = 1'b0;  wr_cycle[ 5996] = 1'b1;  addr_rom[ 5996]='h000038f4;  wr_data_rom[ 5996]='h0000267c;
    rd_cycle[ 5997] = 1'b1;  wr_cycle[ 5997] = 1'b0;  addr_rom[ 5997]='h00000218;  wr_data_rom[ 5997]='h00000000;
    rd_cycle[ 5998] = 1'b0;  wr_cycle[ 5998] = 1'b1;  addr_rom[ 5998]='h000035f4;  wr_data_rom[ 5998]='h00000101;
    rd_cycle[ 5999] = 1'b1;  wr_cycle[ 5999] = 1'b0;  addr_rom[ 5999]='h000004b0;  wr_data_rom[ 5999]='h00000000;
    rd_cycle[ 6000] = 1'b1;  wr_cycle[ 6000] = 1'b0;  addr_rom[ 6000]='h00001a48;  wr_data_rom[ 6000]='h00000000;
    rd_cycle[ 6001] = 1'b0;  wr_cycle[ 6001] = 1'b1;  addr_rom[ 6001]='h00001cdc;  wr_data_rom[ 6001]='h000000b4;
    rd_cycle[ 6002] = 1'b1;  wr_cycle[ 6002] = 1'b0;  addr_rom[ 6002]='h0000368c;  wr_data_rom[ 6002]='h00000000;
    rd_cycle[ 6003] = 1'b0;  wr_cycle[ 6003] = 1'b1;  addr_rom[ 6003]='h00003f48;  wr_data_rom[ 6003]='h000022fa;
    rd_cycle[ 6004] = 1'b0;  wr_cycle[ 6004] = 1'b1;  addr_rom[ 6004]='h00001da4;  wr_data_rom[ 6004]='h00002fc6;
    rd_cycle[ 6005] = 1'b0;  wr_cycle[ 6005] = 1'b1;  addr_rom[ 6005]='h00001810;  wr_data_rom[ 6005]='h000006c5;
    rd_cycle[ 6006] = 1'b0;  wr_cycle[ 6006] = 1'b1;  addr_rom[ 6006]='h000000b4;  wr_data_rom[ 6006]='h000015c7;
    rd_cycle[ 6007] = 1'b0;  wr_cycle[ 6007] = 1'b1;  addr_rom[ 6007]='h000024b4;  wr_data_rom[ 6007]='h000004aa;
    rd_cycle[ 6008] = 1'b0;  wr_cycle[ 6008] = 1'b1;  addr_rom[ 6008]='h0000223c;  wr_data_rom[ 6008]='h000019de;
    rd_cycle[ 6009] = 1'b0;  wr_cycle[ 6009] = 1'b1;  addr_rom[ 6009]='h00002ca0;  wr_data_rom[ 6009]='h00003dfc;
    rd_cycle[ 6010] = 1'b0;  wr_cycle[ 6010] = 1'b1;  addr_rom[ 6010]='h00000aa0;  wr_data_rom[ 6010]='h00002d62;
    rd_cycle[ 6011] = 1'b1;  wr_cycle[ 6011] = 1'b0;  addr_rom[ 6011]='h000023e8;  wr_data_rom[ 6011]='h00000000;
    rd_cycle[ 6012] = 1'b1;  wr_cycle[ 6012] = 1'b0;  addr_rom[ 6012]='h00001be0;  wr_data_rom[ 6012]='h00000000;
    rd_cycle[ 6013] = 1'b0;  wr_cycle[ 6013] = 1'b1;  addr_rom[ 6013]='h000024b0;  wr_data_rom[ 6013]='h00000c53;
    rd_cycle[ 6014] = 1'b0;  wr_cycle[ 6014] = 1'b1;  addr_rom[ 6014]='h00003898;  wr_data_rom[ 6014]='h000010eb;
    rd_cycle[ 6015] = 1'b1;  wr_cycle[ 6015] = 1'b0;  addr_rom[ 6015]='h00000fa4;  wr_data_rom[ 6015]='h00000000;
    rd_cycle[ 6016] = 1'b0;  wr_cycle[ 6016] = 1'b1;  addr_rom[ 6016]='h00003b64;  wr_data_rom[ 6016]='h00000e98;
    rd_cycle[ 6017] = 1'b1;  wr_cycle[ 6017] = 1'b0;  addr_rom[ 6017]='h00003f70;  wr_data_rom[ 6017]='h00000000;
    rd_cycle[ 6018] = 1'b1;  wr_cycle[ 6018] = 1'b0;  addr_rom[ 6018]='h00003bd8;  wr_data_rom[ 6018]='h00000000;
    rd_cycle[ 6019] = 1'b1;  wr_cycle[ 6019] = 1'b0;  addr_rom[ 6019]='h00003000;  wr_data_rom[ 6019]='h00000000;
    rd_cycle[ 6020] = 1'b1;  wr_cycle[ 6020] = 1'b0;  addr_rom[ 6020]='h00002688;  wr_data_rom[ 6020]='h00000000;
    rd_cycle[ 6021] = 1'b0;  wr_cycle[ 6021] = 1'b1;  addr_rom[ 6021]='h00003968;  wr_data_rom[ 6021]='h0000066d;
    rd_cycle[ 6022] = 1'b1;  wr_cycle[ 6022] = 1'b0;  addr_rom[ 6022]='h000005a0;  wr_data_rom[ 6022]='h00000000;
    rd_cycle[ 6023] = 1'b0;  wr_cycle[ 6023] = 1'b1;  addr_rom[ 6023]='h00001b7c;  wr_data_rom[ 6023]='h0000061e;
    rd_cycle[ 6024] = 1'b1;  wr_cycle[ 6024] = 1'b0;  addr_rom[ 6024]='h000023e0;  wr_data_rom[ 6024]='h00000000;
    rd_cycle[ 6025] = 1'b1;  wr_cycle[ 6025] = 1'b0;  addr_rom[ 6025]='h00002d04;  wr_data_rom[ 6025]='h00000000;
    rd_cycle[ 6026] = 1'b1;  wr_cycle[ 6026] = 1'b0;  addr_rom[ 6026]='h00000d58;  wr_data_rom[ 6026]='h00000000;
    rd_cycle[ 6027] = 1'b1;  wr_cycle[ 6027] = 1'b0;  addr_rom[ 6027]='h00001f0c;  wr_data_rom[ 6027]='h00000000;
    rd_cycle[ 6028] = 1'b0;  wr_cycle[ 6028] = 1'b1;  addr_rom[ 6028]='h000036a8;  wr_data_rom[ 6028]='h00003510;
    rd_cycle[ 6029] = 1'b1;  wr_cycle[ 6029] = 1'b0;  addr_rom[ 6029]='h00003564;  wr_data_rom[ 6029]='h00000000;
    rd_cycle[ 6030] = 1'b0;  wr_cycle[ 6030] = 1'b1;  addr_rom[ 6030]='h00002740;  wr_data_rom[ 6030]='h00003a70;
    rd_cycle[ 6031] = 1'b1;  wr_cycle[ 6031] = 1'b0;  addr_rom[ 6031]='h00000818;  wr_data_rom[ 6031]='h00000000;
    rd_cycle[ 6032] = 1'b1;  wr_cycle[ 6032] = 1'b0;  addr_rom[ 6032]='h00002ab0;  wr_data_rom[ 6032]='h00000000;
    rd_cycle[ 6033] = 1'b1;  wr_cycle[ 6033] = 1'b0;  addr_rom[ 6033]='h00002d4c;  wr_data_rom[ 6033]='h00000000;
    rd_cycle[ 6034] = 1'b1;  wr_cycle[ 6034] = 1'b0;  addr_rom[ 6034]='h0000010c;  wr_data_rom[ 6034]='h00000000;
    rd_cycle[ 6035] = 1'b1;  wr_cycle[ 6035] = 1'b0;  addr_rom[ 6035]='h0000174c;  wr_data_rom[ 6035]='h00000000;
    rd_cycle[ 6036] = 1'b0;  wr_cycle[ 6036] = 1'b1;  addr_rom[ 6036]='h000033fc;  wr_data_rom[ 6036]='h00000b32;
    rd_cycle[ 6037] = 1'b0;  wr_cycle[ 6037] = 1'b1;  addr_rom[ 6037]='h000028c4;  wr_data_rom[ 6037]='h00000abc;
    rd_cycle[ 6038] = 1'b0;  wr_cycle[ 6038] = 1'b1;  addr_rom[ 6038]='h000026d4;  wr_data_rom[ 6038]='h00001381;
    rd_cycle[ 6039] = 1'b0;  wr_cycle[ 6039] = 1'b1;  addr_rom[ 6039]='h00002a78;  wr_data_rom[ 6039]='h000008e0;
    rd_cycle[ 6040] = 1'b0;  wr_cycle[ 6040] = 1'b1;  addr_rom[ 6040]='h00000278;  wr_data_rom[ 6040]='h000000b4;
    rd_cycle[ 6041] = 1'b1;  wr_cycle[ 6041] = 1'b0;  addr_rom[ 6041]='h00002a10;  wr_data_rom[ 6041]='h00000000;
    rd_cycle[ 6042] = 1'b0;  wr_cycle[ 6042] = 1'b1;  addr_rom[ 6042]='h00000790;  wr_data_rom[ 6042]='h00000316;
    rd_cycle[ 6043] = 1'b1;  wr_cycle[ 6043] = 1'b0;  addr_rom[ 6043]='h000027d4;  wr_data_rom[ 6043]='h00000000;
    rd_cycle[ 6044] = 1'b0;  wr_cycle[ 6044] = 1'b1;  addr_rom[ 6044]='h000004e0;  wr_data_rom[ 6044]='h00003eaf;
    rd_cycle[ 6045] = 1'b0;  wr_cycle[ 6045] = 1'b1;  addr_rom[ 6045]='h000017f8;  wr_data_rom[ 6045]='h00003f15;
    rd_cycle[ 6046] = 1'b0;  wr_cycle[ 6046] = 1'b1;  addr_rom[ 6046]='h00001dec;  wr_data_rom[ 6046]='h000023a4;
    rd_cycle[ 6047] = 1'b1;  wr_cycle[ 6047] = 1'b0;  addr_rom[ 6047]='h00003680;  wr_data_rom[ 6047]='h00000000;
    rd_cycle[ 6048] = 1'b1;  wr_cycle[ 6048] = 1'b0;  addr_rom[ 6048]='h00002a88;  wr_data_rom[ 6048]='h00000000;
    rd_cycle[ 6049] = 1'b0;  wr_cycle[ 6049] = 1'b1;  addr_rom[ 6049]='h000003f4;  wr_data_rom[ 6049]='h00002a7e;
    rd_cycle[ 6050] = 1'b1;  wr_cycle[ 6050] = 1'b0;  addr_rom[ 6050]='h00002d70;  wr_data_rom[ 6050]='h00000000;
    rd_cycle[ 6051] = 1'b0;  wr_cycle[ 6051] = 1'b1;  addr_rom[ 6051]='h000004d0;  wr_data_rom[ 6051]='h00002c64;
    rd_cycle[ 6052] = 1'b0;  wr_cycle[ 6052] = 1'b1;  addr_rom[ 6052]='h000039fc;  wr_data_rom[ 6052]='h0000226b;
    rd_cycle[ 6053] = 1'b0;  wr_cycle[ 6053] = 1'b1;  addr_rom[ 6053]='h00001da0;  wr_data_rom[ 6053]='h00000aca;
    rd_cycle[ 6054] = 1'b1;  wr_cycle[ 6054] = 1'b0;  addr_rom[ 6054]='h00002aec;  wr_data_rom[ 6054]='h00000000;
    rd_cycle[ 6055] = 1'b1;  wr_cycle[ 6055] = 1'b0;  addr_rom[ 6055]='h00003b24;  wr_data_rom[ 6055]='h00000000;
    rd_cycle[ 6056] = 1'b0;  wr_cycle[ 6056] = 1'b1;  addr_rom[ 6056]='h00002060;  wr_data_rom[ 6056]='h00000679;
    rd_cycle[ 6057] = 1'b0;  wr_cycle[ 6057] = 1'b1;  addr_rom[ 6057]='h00003640;  wr_data_rom[ 6057]='h0000002b;
    rd_cycle[ 6058] = 1'b1;  wr_cycle[ 6058] = 1'b0;  addr_rom[ 6058]='h00001630;  wr_data_rom[ 6058]='h00000000;
    rd_cycle[ 6059] = 1'b1;  wr_cycle[ 6059] = 1'b0;  addr_rom[ 6059]='h00003b24;  wr_data_rom[ 6059]='h00000000;
    rd_cycle[ 6060] = 1'b0;  wr_cycle[ 6060] = 1'b1;  addr_rom[ 6060]='h00003e38;  wr_data_rom[ 6060]='h00003f29;
    rd_cycle[ 6061] = 1'b1;  wr_cycle[ 6061] = 1'b0;  addr_rom[ 6061]='h00000d14;  wr_data_rom[ 6061]='h00000000;
    rd_cycle[ 6062] = 1'b1;  wr_cycle[ 6062] = 1'b0;  addr_rom[ 6062]='h00003c20;  wr_data_rom[ 6062]='h00000000;
    rd_cycle[ 6063] = 1'b0;  wr_cycle[ 6063] = 1'b1;  addr_rom[ 6063]='h000013bc;  wr_data_rom[ 6063]='h00002b7c;
    rd_cycle[ 6064] = 1'b0;  wr_cycle[ 6064] = 1'b1;  addr_rom[ 6064]='h00002654;  wr_data_rom[ 6064]='h00002056;
    rd_cycle[ 6065] = 1'b0;  wr_cycle[ 6065] = 1'b1;  addr_rom[ 6065]='h000001a0;  wr_data_rom[ 6065]='h0000172b;
    rd_cycle[ 6066] = 1'b0;  wr_cycle[ 6066] = 1'b1;  addr_rom[ 6066]='h00002bbc;  wr_data_rom[ 6066]='h00001e45;
    rd_cycle[ 6067] = 1'b1;  wr_cycle[ 6067] = 1'b0;  addr_rom[ 6067]='h000004ec;  wr_data_rom[ 6067]='h00000000;
    rd_cycle[ 6068] = 1'b0;  wr_cycle[ 6068] = 1'b1;  addr_rom[ 6068]='h00000d4c;  wr_data_rom[ 6068]='h00000df9;
    rd_cycle[ 6069] = 1'b0;  wr_cycle[ 6069] = 1'b1;  addr_rom[ 6069]='h00002bf8;  wr_data_rom[ 6069]='h00001a3f;
    rd_cycle[ 6070] = 1'b1;  wr_cycle[ 6070] = 1'b0;  addr_rom[ 6070]='h00001b70;  wr_data_rom[ 6070]='h00000000;
    rd_cycle[ 6071] = 1'b0;  wr_cycle[ 6071] = 1'b1;  addr_rom[ 6071]='h00000fec;  wr_data_rom[ 6071]='h0000350e;
    rd_cycle[ 6072] = 1'b0;  wr_cycle[ 6072] = 1'b1;  addr_rom[ 6072]='h00001900;  wr_data_rom[ 6072]='h00002d38;
    rd_cycle[ 6073] = 1'b1;  wr_cycle[ 6073] = 1'b0;  addr_rom[ 6073]='h00003f28;  wr_data_rom[ 6073]='h00000000;
    rd_cycle[ 6074] = 1'b1;  wr_cycle[ 6074] = 1'b0;  addr_rom[ 6074]='h000037d4;  wr_data_rom[ 6074]='h00000000;
    rd_cycle[ 6075] = 1'b0;  wr_cycle[ 6075] = 1'b1;  addr_rom[ 6075]='h00001824;  wr_data_rom[ 6075]='h00000bad;
    rd_cycle[ 6076] = 1'b0;  wr_cycle[ 6076] = 1'b1;  addr_rom[ 6076]='h00003a5c;  wr_data_rom[ 6076]='h00000948;
    rd_cycle[ 6077] = 1'b0;  wr_cycle[ 6077] = 1'b1;  addr_rom[ 6077]='h000023b4;  wr_data_rom[ 6077]='h000020a5;
    rd_cycle[ 6078] = 1'b1;  wr_cycle[ 6078] = 1'b0;  addr_rom[ 6078]='h00000c3c;  wr_data_rom[ 6078]='h00000000;
    rd_cycle[ 6079] = 1'b0;  wr_cycle[ 6079] = 1'b1;  addr_rom[ 6079]='h00000500;  wr_data_rom[ 6079]='h0000197d;
    rd_cycle[ 6080] = 1'b0;  wr_cycle[ 6080] = 1'b1;  addr_rom[ 6080]='h00001720;  wr_data_rom[ 6080]='h00003141;
    rd_cycle[ 6081] = 1'b1;  wr_cycle[ 6081] = 1'b0;  addr_rom[ 6081]='h00002dec;  wr_data_rom[ 6081]='h00000000;
    rd_cycle[ 6082] = 1'b0;  wr_cycle[ 6082] = 1'b1;  addr_rom[ 6082]='h000028c8;  wr_data_rom[ 6082]='h00003f47;
    rd_cycle[ 6083] = 1'b1;  wr_cycle[ 6083] = 1'b0;  addr_rom[ 6083]='h00000908;  wr_data_rom[ 6083]='h00000000;
    rd_cycle[ 6084] = 1'b0;  wr_cycle[ 6084] = 1'b1;  addr_rom[ 6084]='h00002c94;  wr_data_rom[ 6084]='h000027ba;
    rd_cycle[ 6085] = 1'b1;  wr_cycle[ 6085] = 1'b0;  addr_rom[ 6085]='h00002b04;  wr_data_rom[ 6085]='h00000000;
    rd_cycle[ 6086] = 1'b0;  wr_cycle[ 6086] = 1'b1;  addr_rom[ 6086]='h00003eec;  wr_data_rom[ 6086]='h00003a7a;
    rd_cycle[ 6087] = 1'b0;  wr_cycle[ 6087] = 1'b1;  addr_rom[ 6087]='h00000cbc;  wr_data_rom[ 6087]='h000001c3;
    rd_cycle[ 6088] = 1'b0;  wr_cycle[ 6088] = 1'b1;  addr_rom[ 6088]='h00002dc8;  wr_data_rom[ 6088]='h000029d9;
    rd_cycle[ 6089] = 1'b1;  wr_cycle[ 6089] = 1'b0;  addr_rom[ 6089]='h0000058c;  wr_data_rom[ 6089]='h00000000;
    rd_cycle[ 6090] = 1'b1;  wr_cycle[ 6090] = 1'b0;  addr_rom[ 6090]='h00000c50;  wr_data_rom[ 6090]='h00000000;
    rd_cycle[ 6091] = 1'b0;  wr_cycle[ 6091] = 1'b1;  addr_rom[ 6091]='h00000394;  wr_data_rom[ 6091]='h00002dda;
    rd_cycle[ 6092] = 1'b0;  wr_cycle[ 6092] = 1'b1;  addr_rom[ 6092]='h00002b88;  wr_data_rom[ 6092]='h0000243f;
    rd_cycle[ 6093] = 1'b0;  wr_cycle[ 6093] = 1'b1;  addr_rom[ 6093]='h000009a8;  wr_data_rom[ 6093]='h00002fe4;
    rd_cycle[ 6094] = 1'b0;  wr_cycle[ 6094] = 1'b1;  addr_rom[ 6094]='h00003bd8;  wr_data_rom[ 6094]='h00001d40;
    rd_cycle[ 6095] = 1'b1;  wr_cycle[ 6095] = 1'b0;  addr_rom[ 6095]='h00002654;  wr_data_rom[ 6095]='h00000000;
    rd_cycle[ 6096] = 1'b1;  wr_cycle[ 6096] = 1'b0;  addr_rom[ 6096]='h00001614;  wr_data_rom[ 6096]='h00000000;
    rd_cycle[ 6097] = 1'b0;  wr_cycle[ 6097] = 1'b1;  addr_rom[ 6097]='h00002ab8;  wr_data_rom[ 6097]='h00003068;
    rd_cycle[ 6098] = 1'b1;  wr_cycle[ 6098] = 1'b0;  addr_rom[ 6098]='h00002ca0;  wr_data_rom[ 6098]='h00000000;
    rd_cycle[ 6099] = 1'b1;  wr_cycle[ 6099] = 1'b0;  addr_rom[ 6099]='h00001344;  wr_data_rom[ 6099]='h00000000;
    rd_cycle[ 6100] = 1'b0;  wr_cycle[ 6100] = 1'b1;  addr_rom[ 6100]='h00002710;  wr_data_rom[ 6100]='h00001c6f;
    rd_cycle[ 6101] = 1'b0;  wr_cycle[ 6101] = 1'b1;  addr_rom[ 6101]='h00001c9c;  wr_data_rom[ 6101]='h000003f6;
    rd_cycle[ 6102] = 1'b0;  wr_cycle[ 6102] = 1'b1;  addr_rom[ 6102]='h000025d4;  wr_data_rom[ 6102]='h000034af;
    rd_cycle[ 6103] = 1'b1;  wr_cycle[ 6103] = 1'b0;  addr_rom[ 6103]='h00000f5c;  wr_data_rom[ 6103]='h00000000;
    rd_cycle[ 6104] = 1'b1;  wr_cycle[ 6104] = 1'b0;  addr_rom[ 6104]='h00001768;  wr_data_rom[ 6104]='h00000000;
    rd_cycle[ 6105] = 1'b1;  wr_cycle[ 6105] = 1'b0;  addr_rom[ 6105]='h00000514;  wr_data_rom[ 6105]='h00000000;
    rd_cycle[ 6106] = 1'b1;  wr_cycle[ 6106] = 1'b0;  addr_rom[ 6106]='h00000580;  wr_data_rom[ 6106]='h00000000;
    rd_cycle[ 6107] = 1'b0;  wr_cycle[ 6107] = 1'b1;  addr_rom[ 6107]='h00001420;  wr_data_rom[ 6107]='h00001a43;
    rd_cycle[ 6108] = 1'b1;  wr_cycle[ 6108] = 1'b0;  addr_rom[ 6108]='h00000e68;  wr_data_rom[ 6108]='h00000000;
    rd_cycle[ 6109] = 1'b1;  wr_cycle[ 6109] = 1'b0;  addr_rom[ 6109]='h000009b0;  wr_data_rom[ 6109]='h00000000;
    rd_cycle[ 6110] = 1'b0;  wr_cycle[ 6110] = 1'b1;  addr_rom[ 6110]='h000016a8;  wr_data_rom[ 6110]='h0000384b;
    rd_cycle[ 6111] = 1'b1;  wr_cycle[ 6111] = 1'b0;  addr_rom[ 6111]='h00001acc;  wr_data_rom[ 6111]='h00000000;
    rd_cycle[ 6112] = 1'b1;  wr_cycle[ 6112] = 1'b0;  addr_rom[ 6112]='h00002a60;  wr_data_rom[ 6112]='h00000000;
    rd_cycle[ 6113] = 1'b0;  wr_cycle[ 6113] = 1'b1;  addr_rom[ 6113]='h00002690;  wr_data_rom[ 6113]='h000015a5;
    rd_cycle[ 6114] = 1'b1;  wr_cycle[ 6114] = 1'b0;  addr_rom[ 6114]='h000020c4;  wr_data_rom[ 6114]='h00000000;
    rd_cycle[ 6115] = 1'b0;  wr_cycle[ 6115] = 1'b1;  addr_rom[ 6115]='h00001c20;  wr_data_rom[ 6115]='h00000ab0;
    rd_cycle[ 6116] = 1'b0;  wr_cycle[ 6116] = 1'b1;  addr_rom[ 6116]='h00003ed0;  wr_data_rom[ 6116]='h0000022c;
    rd_cycle[ 6117] = 1'b1;  wr_cycle[ 6117] = 1'b0;  addr_rom[ 6117]='h00002e4c;  wr_data_rom[ 6117]='h00000000;
    rd_cycle[ 6118] = 1'b1;  wr_cycle[ 6118] = 1'b0;  addr_rom[ 6118]='h000010b8;  wr_data_rom[ 6118]='h00000000;
    rd_cycle[ 6119] = 1'b0;  wr_cycle[ 6119] = 1'b1;  addr_rom[ 6119]='h00003fb0;  wr_data_rom[ 6119]='h0000263f;
    rd_cycle[ 6120] = 1'b0;  wr_cycle[ 6120] = 1'b1;  addr_rom[ 6120]='h00000eb8;  wr_data_rom[ 6120]='h00001a61;
    rd_cycle[ 6121] = 1'b1;  wr_cycle[ 6121] = 1'b0;  addr_rom[ 6121]='h0000023c;  wr_data_rom[ 6121]='h00000000;
    rd_cycle[ 6122] = 1'b0;  wr_cycle[ 6122] = 1'b1;  addr_rom[ 6122]='h00003144;  wr_data_rom[ 6122]='h000019b8;
    rd_cycle[ 6123] = 1'b1;  wr_cycle[ 6123] = 1'b0;  addr_rom[ 6123]='h000000dc;  wr_data_rom[ 6123]='h00000000;
    rd_cycle[ 6124] = 1'b0;  wr_cycle[ 6124] = 1'b1;  addr_rom[ 6124]='h00001f44;  wr_data_rom[ 6124]='h00001734;
    rd_cycle[ 6125] = 1'b1;  wr_cycle[ 6125] = 1'b0;  addr_rom[ 6125]='h00003f2c;  wr_data_rom[ 6125]='h00000000;
    rd_cycle[ 6126] = 1'b1;  wr_cycle[ 6126] = 1'b0;  addr_rom[ 6126]='h00003924;  wr_data_rom[ 6126]='h00000000;
    rd_cycle[ 6127] = 1'b1;  wr_cycle[ 6127] = 1'b0;  addr_rom[ 6127]='h00002614;  wr_data_rom[ 6127]='h00000000;
    rd_cycle[ 6128] = 1'b0;  wr_cycle[ 6128] = 1'b1;  addr_rom[ 6128]='h0000345c;  wr_data_rom[ 6128]='h00001530;
    rd_cycle[ 6129] = 1'b0;  wr_cycle[ 6129] = 1'b1;  addr_rom[ 6129]='h00003954;  wr_data_rom[ 6129]='h00000913;
    rd_cycle[ 6130] = 1'b0;  wr_cycle[ 6130] = 1'b1;  addr_rom[ 6130]='h00001c84;  wr_data_rom[ 6130]='h00003bb6;
    rd_cycle[ 6131] = 1'b0;  wr_cycle[ 6131] = 1'b1;  addr_rom[ 6131]='h00003490;  wr_data_rom[ 6131]='h0000134b;
    rd_cycle[ 6132] = 1'b0;  wr_cycle[ 6132] = 1'b1;  addr_rom[ 6132]='h00002014;  wr_data_rom[ 6132]='h00002178;
    rd_cycle[ 6133] = 1'b0;  wr_cycle[ 6133] = 1'b1;  addr_rom[ 6133]='h0000318c;  wr_data_rom[ 6133]='h00001895;
    rd_cycle[ 6134] = 1'b1;  wr_cycle[ 6134] = 1'b0;  addr_rom[ 6134]='h00003ff4;  wr_data_rom[ 6134]='h00000000;
    rd_cycle[ 6135] = 1'b0;  wr_cycle[ 6135] = 1'b1;  addr_rom[ 6135]='h00000b44;  wr_data_rom[ 6135]='h00002f48;
    rd_cycle[ 6136] = 1'b0;  wr_cycle[ 6136] = 1'b1;  addr_rom[ 6136]='h00001d7c;  wr_data_rom[ 6136]='h00000a3c;
    rd_cycle[ 6137] = 1'b0;  wr_cycle[ 6137] = 1'b1;  addr_rom[ 6137]='h00003f90;  wr_data_rom[ 6137]='h0000165c;
    rd_cycle[ 6138] = 1'b0;  wr_cycle[ 6138] = 1'b1;  addr_rom[ 6138]='h000012d8;  wr_data_rom[ 6138]='h00000fd9;
    rd_cycle[ 6139] = 1'b1;  wr_cycle[ 6139] = 1'b0;  addr_rom[ 6139]='h00003c48;  wr_data_rom[ 6139]='h00000000;
    rd_cycle[ 6140] = 1'b0;  wr_cycle[ 6140] = 1'b1;  addr_rom[ 6140]='h00002864;  wr_data_rom[ 6140]='h00003333;
    rd_cycle[ 6141] = 1'b1;  wr_cycle[ 6141] = 1'b0;  addr_rom[ 6141]='h000039c0;  wr_data_rom[ 6141]='h00000000;
    rd_cycle[ 6142] = 1'b0;  wr_cycle[ 6142] = 1'b1;  addr_rom[ 6142]='h00000180;  wr_data_rom[ 6142]='h000019d9;
    rd_cycle[ 6143] = 1'b0;  wr_cycle[ 6143] = 1'b1;  addr_rom[ 6143]='h00001774;  wr_data_rom[ 6143]='h00000bca;
    rd_cycle[ 6144] = 1'b1;  wr_cycle[ 6144] = 1'b0;  addr_rom[ 6144]='h0000142c;  wr_data_rom[ 6144]='h00000000;
    rd_cycle[ 6145] = 1'b1;  wr_cycle[ 6145] = 1'b0;  addr_rom[ 6145]='h0000140c;  wr_data_rom[ 6145]='h00000000;
    rd_cycle[ 6146] = 1'b0;  wr_cycle[ 6146] = 1'b1;  addr_rom[ 6146]='h000020c0;  wr_data_rom[ 6146]='h00000874;
    rd_cycle[ 6147] = 1'b0;  wr_cycle[ 6147] = 1'b1;  addr_rom[ 6147]='h00000770;  wr_data_rom[ 6147]='h0000287a;
    rd_cycle[ 6148] = 1'b1;  wr_cycle[ 6148] = 1'b0;  addr_rom[ 6148]='h000001d8;  wr_data_rom[ 6148]='h00000000;
    rd_cycle[ 6149] = 1'b1;  wr_cycle[ 6149] = 1'b0;  addr_rom[ 6149]='h00000b2c;  wr_data_rom[ 6149]='h00000000;
    rd_cycle[ 6150] = 1'b1;  wr_cycle[ 6150] = 1'b0;  addr_rom[ 6150]='h00000778;  wr_data_rom[ 6150]='h00000000;
    rd_cycle[ 6151] = 1'b0;  wr_cycle[ 6151] = 1'b1;  addr_rom[ 6151]='h00001438;  wr_data_rom[ 6151]='h0000255c;
    rd_cycle[ 6152] = 1'b1;  wr_cycle[ 6152] = 1'b0;  addr_rom[ 6152]='h000032a8;  wr_data_rom[ 6152]='h00000000;
    rd_cycle[ 6153] = 1'b0;  wr_cycle[ 6153] = 1'b1;  addr_rom[ 6153]='h00000f84;  wr_data_rom[ 6153]='h00002627;
    rd_cycle[ 6154] = 1'b1;  wr_cycle[ 6154] = 1'b0;  addr_rom[ 6154]='h00002c7c;  wr_data_rom[ 6154]='h00000000;
    rd_cycle[ 6155] = 1'b0;  wr_cycle[ 6155] = 1'b1;  addr_rom[ 6155]='h00003f20;  wr_data_rom[ 6155]='h00003348;
    rd_cycle[ 6156] = 1'b0;  wr_cycle[ 6156] = 1'b1;  addr_rom[ 6156]='h000035c8;  wr_data_rom[ 6156]='h000030b4;
    rd_cycle[ 6157] = 1'b0;  wr_cycle[ 6157] = 1'b1;  addr_rom[ 6157]='h0000169c;  wr_data_rom[ 6157]='h000029db;
    rd_cycle[ 6158] = 1'b1;  wr_cycle[ 6158] = 1'b0;  addr_rom[ 6158]='h000011d8;  wr_data_rom[ 6158]='h00000000;
    rd_cycle[ 6159] = 1'b0;  wr_cycle[ 6159] = 1'b1;  addr_rom[ 6159]='h00000b70;  wr_data_rom[ 6159]='h000026a1;
    rd_cycle[ 6160] = 1'b0;  wr_cycle[ 6160] = 1'b1;  addr_rom[ 6160]='h00000fc0;  wr_data_rom[ 6160]='h00003c8c;
    rd_cycle[ 6161] = 1'b0;  wr_cycle[ 6161] = 1'b1;  addr_rom[ 6161]='h00001f2c;  wr_data_rom[ 6161]='h00001263;
    rd_cycle[ 6162] = 1'b1;  wr_cycle[ 6162] = 1'b0;  addr_rom[ 6162]='h000012c0;  wr_data_rom[ 6162]='h00000000;
    rd_cycle[ 6163] = 1'b0;  wr_cycle[ 6163] = 1'b1;  addr_rom[ 6163]='h00001690;  wr_data_rom[ 6163]='h00001fab;
    rd_cycle[ 6164] = 1'b0;  wr_cycle[ 6164] = 1'b1;  addr_rom[ 6164]='h00003994;  wr_data_rom[ 6164]='h00003b38;
    rd_cycle[ 6165] = 1'b0;  wr_cycle[ 6165] = 1'b1;  addr_rom[ 6165]='h00002280;  wr_data_rom[ 6165]='h00003624;
    rd_cycle[ 6166] = 1'b1;  wr_cycle[ 6166] = 1'b0;  addr_rom[ 6166]='h000027d0;  wr_data_rom[ 6166]='h00000000;
    rd_cycle[ 6167] = 1'b1;  wr_cycle[ 6167] = 1'b0;  addr_rom[ 6167]='h00001124;  wr_data_rom[ 6167]='h00000000;
    rd_cycle[ 6168] = 1'b0;  wr_cycle[ 6168] = 1'b1;  addr_rom[ 6168]='h00000278;  wr_data_rom[ 6168]='h00000700;
    rd_cycle[ 6169] = 1'b0;  wr_cycle[ 6169] = 1'b1;  addr_rom[ 6169]='h00002c30;  wr_data_rom[ 6169]='h00000bb7;
    rd_cycle[ 6170] = 1'b1;  wr_cycle[ 6170] = 1'b0;  addr_rom[ 6170]='h00003dd8;  wr_data_rom[ 6170]='h00000000;
    rd_cycle[ 6171] = 1'b1;  wr_cycle[ 6171] = 1'b0;  addr_rom[ 6171]='h000006b0;  wr_data_rom[ 6171]='h00000000;
    rd_cycle[ 6172] = 1'b0;  wr_cycle[ 6172] = 1'b1;  addr_rom[ 6172]='h0000101c;  wr_data_rom[ 6172]='h000031ea;
    rd_cycle[ 6173] = 1'b1;  wr_cycle[ 6173] = 1'b0;  addr_rom[ 6173]='h00001df8;  wr_data_rom[ 6173]='h00000000;
    rd_cycle[ 6174] = 1'b1;  wr_cycle[ 6174] = 1'b0;  addr_rom[ 6174]='h00003194;  wr_data_rom[ 6174]='h00000000;
    rd_cycle[ 6175] = 1'b0;  wr_cycle[ 6175] = 1'b1;  addr_rom[ 6175]='h00002b78;  wr_data_rom[ 6175]='h00001c72;
    rd_cycle[ 6176] = 1'b0;  wr_cycle[ 6176] = 1'b1;  addr_rom[ 6176]='h000002e4;  wr_data_rom[ 6176]='h00000053;
    rd_cycle[ 6177] = 1'b1;  wr_cycle[ 6177] = 1'b0;  addr_rom[ 6177]='h000011c4;  wr_data_rom[ 6177]='h00000000;
    rd_cycle[ 6178] = 1'b0;  wr_cycle[ 6178] = 1'b1;  addr_rom[ 6178]='h00003c20;  wr_data_rom[ 6178]='h000000fa;
    rd_cycle[ 6179] = 1'b1;  wr_cycle[ 6179] = 1'b0;  addr_rom[ 6179]='h00003220;  wr_data_rom[ 6179]='h00000000;
    rd_cycle[ 6180] = 1'b1;  wr_cycle[ 6180] = 1'b0;  addr_rom[ 6180]='h00000620;  wr_data_rom[ 6180]='h00000000;
    rd_cycle[ 6181] = 1'b1;  wr_cycle[ 6181] = 1'b0;  addr_rom[ 6181]='h000031d4;  wr_data_rom[ 6181]='h00000000;
    rd_cycle[ 6182] = 1'b1;  wr_cycle[ 6182] = 1'b0;  addr_rom[ 6182]='h0000003c;  wr_data_rom[ 6182]='h00000000;
    rd_cycle[ 6183] = 1'b0;  wr_cycle[ 6183] = 1'b1;  addr_rom[ 6183]='h00003408;  wr_data_rom[ 6183]='h000030ce;
    rd_cycle[ 6184] = 1'b1;  wr_cycle[ 6184] = 1'b0;  addr_rom[ 6184]='h00000680;  wr_data_rom[ 6184]='h00000000;
    rd_cycle[ 6185] = 1'b1;  wr_cycle[ 6185] = 1'b0;  addr_rom[ 6185]='h00002bdc;  wr_data_rom[ 6185]='h00000000;
    rd_cycle[ 6186] = 1'b1;  wr_cycle[ 6186] = 1'b0;  addr_rom[ 6186]='h00003658;  wr_data_rom[ 6186]='h00000000;
    rd_cycle[ 6187] = 1'b1;  wr_cycle[ 6187] = 1'b0;  addr_rom[ 6187]='h000005d8;  wr_data_rom[ 6187]='h00000000;
    rd_cycle[ 6188] = 1'b0;  wr_cycle[ 6188] = 1'b1;  addr_rom[ 6188]='h00001da8;  wr_data_rom[ 6188]='h000008af;
    rd_cycle[ 6189] = 1'b0;  wr_cycle[ 6189] = 1'b1;  addr_rom[ 6189]='h000013dc;  wr_data_rom[ 6189]='h00002e78;
    rd_cycle[ 6190] = 1'b0;  wr_cycle[ 6190] = 1'b1;  addr_rom[ 6190]='h00003664;  wr_data_rom[ 6190]='h000030a4;
    rd_cycle[ 6191] = 1'b0;  wr_cycle[ 6191] = 1'b1;  addr_rom[ 6191]='h00000d6c;  wr_data_rom[ 6191]='h00000219;
    rd_cycle[ 6192] = 1'b0;  wr_cycle[ 6192] = 1'b1;  addr_rom[ 6192]='h00000458;  wr_data_rom[ 6192]='h000010b4;
    rd_cycle[ 6193] = 1'b0;  wr_cycle[ 6193] = 1'b1;  addr_rom[ 6193]='h00000238;  wr_data_rom[ 6193]='h00001a29;
    rd_cycle[ 6194] = 1'b0;  wr_cycle[ 6194] = 1'b1;  addr_rom[ 6194]='h00003e70;  wr_data_rom[ 6194]='h0000318d;
    rd_cycle[ 6195] = 1'b0;  wr_cycle[ 6195] = 1'b1;  addr_rom[ 6195]='h0000156c;  wr_data_rom[ 6195]='h0000204c;
    rd_cycle[ 6196] = 1'b1;  wr_cycle[ 6196] = 1'b0;  addr_rom[ 6196]='h000032ac;  wr_data_rom[ 6196]='h00000000;
    rd_cycle[ 6197] = 1'b0;  wr_cycle[ 6197] = 1'b1;  addr_rom[ 6197]='h00000460;  wr_data_rom[ 6197]='h00003dca;
    rd_cycle[ 6198] = 1'b0;  wr_cycle[ 6198] = 1'b1;  addr_rom[ 6198]='h00000880;  wr_data_rom[ 6198]='h00000f9e;
    rd_cycle[ 6199] = 1'b1;  wr_cycle[ 6199] = 1'b0;  addr_rom[ 6199]='h00000514;  wr_data_rom[ 6199]='h00000000;
    rd_cycle[ 6200] = 1'b1;  wr_cycle[ 6200] = 1'b0;  addr_rom[ 6200]='h00002fdc;  wr_data_rom[ 6200]='h00000000;
    rd_cycle[ 6201] = 1'b0;  wr_cycle[ 6201] = 1'b1;  addr_rom[ 6201]='h00002e0c;  wr_data_rom[ 6201]='h00003eec;
    rd_cycle[ 6202] = 1'b1;  wr_cycle[ 6202] = 1'b0;  addr_rom[ 6202]='h0000330c;  wr_data_rom[ 6202]='h00000000;
    rd_cycle[ 6203] = 1'b1;  wr_cycle[ 6203] = 1'b0;  addr_rom[ 6203]='h0000226c;  wr_data_rom[ 6203]='h00000000;
    rd_cycle[ 6204] = 1'b1;  wr_cycle[ 6204] = 1'b0;  addr_rom[ 6204]='h0000011c;  wr_data_rom[ 6204]='h00000000;
    rd_cycle[ 6205] = 1'b1;  wr_cycle[ 6205] = 1'b0;  addr_rom[ 6205]='h00003fcc;  wr_data_rom[ 6205]='h00000000;
    rd_cycle[ 6206] = 1'b0;  wr_cycle[ 6206] = 1'b1;  addr_rom[ 6206]='h00001d44;  wr_data_rom[ 6206]='h00001a5d;
    rd_cycle[ 6207] = 1'b0;  wr_cycle[ 6207] = 1'b1;  addr_rom[ 6207]='h00003964;  wr_data_rom[ 6207]='h000028c0;
    rd_cycle[ 6208] = 1'b0;  wr_cycle[ 6208] = 1'b1;  addr_rom[ 6208]='h00000d70;  wr_data_rom[ 6208]='h000017d0;
    rd_cycle[ 6209] = 1'b0;  wr_cycle[ 6209] = 1'b1;  addr_rom[ 6209]='h00003998;  wr_data_rom[ 6209]='h00001b22;
    rd_cycle[ 6210] = 1'b1;  wr_cycle[ 6210] = 1'b0;  addr_rom[ 6210]='h00000560;  wr_data_rom[ 6210]='h00000000;
    rd_cycle[ 6211] = 1'b1;  wr_cycle[ 6211] = 1'b0;  addr_rom[ 6211]='h00001c50;  wr_data_rom[ 6211]='h00000000;
    rd_cycle[ 6212] = 1'b0;  wr_cycle[ 6212] = 1'b1;  addr_rom[ 6212]='h00000380;  wr_data_rom[ 6212]='h00002fe6;
    rd_cycle[ 6213] = 1'b0;  wr_cycle[ 6213] = 1'b1;  addr_rom[ 6213]='h00001ab0;  wr_data_rom[ 6213]='h00003dbd;
    rd_cycle[ 6214] = 1'b1;  wr_cycle[ 6214] = 1'b0;  addr_rom[ 6214]='h0000271c;  wr_data_rom[ 6214]='h00000000;
    rd_cycle[ 6215] = 1'b1;  wr_cycle[ 6215] = 1'b0;  addr_rom[ 6215]='h00000f0c;  wr_data_rom[ 6215]='h00000000;
    rd_cycle[ 6216] = 1'b0;  wr_cycle[ 6216] = 1'b1;  addr_rom[ 6216]='h0000187c;  wr_data_rom[ 6216]='h00003113;
    rd_cycle[ 6217] = 1'b1;  wr_cycle[ 6217] = 1'b0;  addr_rom[ 6217]='h00001aa8;  wr_data_rom[ 6217]='h00000000;
    rd_cycle[ 6218] = 1'b1;  wr_cycle[ 6218] = 1'b0;  addr_rom[ 6218]='h00000820;  wr_data_rom[ 6218]='h00000000;
    rd_cycle[ 6219] = 1'b1;  wr_cycle[ 6219] = 1'b0;  addr_rom[ 6219]='h00000008;  wr_data_rom[ 6219]='h00000000;
    rd_cycle[ 6220] = 1'b1;  wr_cycle[ 6220] = 1'b0;  addr_rom[ 6220]='h000028cc;  wr_data_rom[ 6220]='h00000000;
    rd_cycle[ 6221] = 1'b1;  wr_cycle[ 6221] = 1'b0;  addr_rom[ 6221]='h00002cc4;  wr_data_rom[ 6221]='h00000000;
    rd_cycle[ 6222] = 1'b0;  wr_cycle[ 6222] = 1'b1;  addr_rom[ 6222]='h000006b0;  wr_data_rom[ 6222]='h00001add;
    rd_cycle[ 6223] = 1'b1;  wr_cycle[ 6223] = 1'b0;  addr_rom[ 6223]='h00000304;  wr_data_rom[ 6223]='h00000000;
    rd_cycle[ 6224] = 1'b1;  wr_cycle[ 6224] = 1'b0;  addr_rom[ 6224]='h000035fc;  wr_data_rom[ 6224]='h00000000;
    rd_cycle[ 6225] = 1'b0;  wr_cycle[ 6225] = 1'b1;  addr_rom[ 6225]='h000026f4;  wr_data_rom[ 6225]='h000037fd;
    rd_cycle[ 6226] = 1'b1;  wr_cycle[ 6226] = 1'b0;  addr_rom[ 6226]='h00003b30;  wr_data_rom[ 6226]='h00000000;
    rd_cycle[ 6227] = 1'b0;  wr_cycle[ 6227] = 1'b1;  addr_rom[ 6227]='h00000250;  wr_data_rom[ 6227]='h00002eb9;
    rd_cycle[ 6228] = 1'b0;  wr_cycle[ 6228] = 1'b1;  addr_rom[ 6228]='h00002c9c;  wr_data_rom[ 6228]='h00001cb5;
    rd_cycle[ 6229] = 1'b0;  wr_cycle[ 6229] = 1'b1;  addr_rom[ 6229]='h0000149c;  wr_data_rom[ 6229]='h00002bbf;
    rd_cycle[ 6230] = 1'b1;  wr_cycle[ 6230] = 1'b0;  addr_rom[ 6230]='h00001ab8;  wr_data_rom[ 6230]='h00000000;
    rd_cycle[ 6231] = 1'b1;  wr_cycle[ 6231] = 1'b0;  addr_rom[ 6231]='h00000db4;  wr_data_rom[ 6231]='h00000000;
    rd_cycle[ 6232] = 1'b0;  wr_cycle[ 6232] = 1'b1;  addr_rom[ 6232]='h0000061c;  wr_data_rom[ 6232]='h00000edf;
    rd_cycle[ 6233] = 1'b0;  wr_cycle[ 6233] = 1'b1;  addr_rom[ 6233]='h00001e44;  wr_data_rom[ 6233]='h0000223e;
    rd_cycle[ 6234] = 1'b1;  wr_cycle[ 6234] = 1'b0;  addr_rom[ 6234]='h000031a8;  wr_data_rom[ 6234]='h00000000;
    rd_cycle[ 6235] = 1'b1;  wr_cycle[ 6235] = 1'b0;  addr_rom[ 6235]='h00002c44;  wr_data_rom[ 6235]='h00000000;
    rd_cycle[ 6236] = 1'b0;  wr_cycle[ 6236] = 1'b1;  addr_rom[ 6236]='h000006d4;  wr_data_rom[ 6236]='h00000510;
    rd_cycle[ 6237] = 1'b0;  wr_cycle[ 6237] = 1'b1;  addr_rom[ 6237]='h00001d70;  wr_data_rom[ 6237]='h00002e77;
    rd_cycle[ 6238] = 1'b1;  wr_cycle[ 6238] = 1'b0;  addr_rom[ 6238]='h00000ac4;  wr_data_rom[ 6238]='h00000000;
    rd_cycle[ 6239] = 1'b0;  wr_cycle[ 6239] = 1'b1;  addr_rom[ 6239]='h00001e28;  wr_data_rom[ 6239]='h0000092d;
    rd_cycle[ 6240] = 1'b0;  wr_cycle[ 6240] = 1'b1;  addr_rom[ 6240]='h00002d88;  wr_data_rom[ 6240]='h00001914;
    rd_cycle[ 6241] = 1'b1;  wr_cycle[ 6241] = 1'b0;  addr_rom[ 6241]='h00001040;  wr_data_rom[ 6241]='h00000000;
    rd_cycle[ 6242] = 1'b1;  wr_cycle[ 6242] = 1'b0;  addr_rom[ 6242]='h00002d9c;  wr_data_rom[ 6242]='h00000000;
    rd_cycle[ 6243] = 1'b1;  wr_cycle[ 6243] = 1'b0;  addr_rom[ 6243]='h00002330;  wr_data_rom[ 6243]='h00000000;
    rd_cycle[ 6244] = 1'b1;  wr_cycle[ 6244] = 1'b0;  addr_rom[ 6244]='h00000fb8;  wr_data_rom[ 6244]='h00000000;
    rd_cycle[ 6245] = 1'b0;  wr_cycle[ 6245] = 1'b1;  addr_rom[ 6245]='h00001f7c;  wr_data_rom[ 6245]='h0000087f;
    rd_cycle[ 6246] = 1'b0;  wr_cycle[ 6246] = 1'b1;  addr_rom[ 6246]='h00001a24;  wr_data_rom[ 6246]='h000007bf;
    rd_cycle[ 6247] = 1'b0;  wr_cycle[ 6247] = 1'b1;  addr_rom[ 6247]='h00003d74;  wr_data_rom[ 6247]='h00001975;
    rd_cycle[ 6248] = 1'b1;  wr_cycle[ 6248] = 1'b0;  addr_rom[ 6248]='h00001010;  wr_data_rom[ 6248]='h00000000;
    rd_cycle[ 6249] = 1'b0;  wr_cycle[ 6249] = 1'b1;  addr_rom[ 6249]='h00002794;  wr_data_rom[ 6249]='h000037d9;
    rd_cycle[ 6250] = 1'b1;  wr_cycle[ 6250] = 1'b0;  addr_rom[ 6250]='h000035f4;  wr_data_rom[ 6250]='h00000000;
    rd_cycle[ 6251] = 1'b0;  wr_cycle[ 6251] = 1'b1;  addr_rom[ 6251]='h00000b18;  wr_data_rom[ 6251]='h00003477;
    rd_cycle[ 6252] = 1'b1;  wr_cycle[ 6252] = 1'b0;  addr_rom[ 6252]='h00003f04;  wr_data_rom[ 6252]='h00000000;
    rd_cycle[ 6253] = 1'b1;  wr_cycle[ 6253] = 1'b0;  addr_rom[ 6253]='h00002c6c;  wr_data_rom[ 6253]='h00000000;
    rd_cycle[ 6254] = 1'b1;  wr_cycle[ 6254] = 1'b0;  addr_rom[ 6254]='h00001f00;  wr_data_rom[ 6254]='h00000000;
    rd_cycle[ 6255] = 1'b0;  wr_cycle[ 6255] = 1'b1;  addr_rom[ 6255]='h000000f0;  wr_data_rom[ 6255]='h0000376b;
    rd_cycle[ 6256] = 1'b1;  wr_cycle[ 6256] = 1'b0;  addr_rom[ 6256]='h000019c8;  wr_data_rom[ 6256]='h00000000;
    rd_cycle[ 6257] = 1'b0;  wr_cycle[ 6257] = 1'b1;  addr_rom[ 6257]='h000025b8;  wr_data_rom[ 6257]='h00003349;
    rd_cycle[ 6258] = 1'b1;  wr_cycle[ 6258] = 1'b0;  addr_rom[ 6258]='h00003638;  wr_data_rom[ 6258]='h00000000;
    rd_cycle[ 6259] = 1'b1;  wr_cycle[ 6259] = 1'b0;  addr_rom[ 6259]='h00002ec4;  wr_data_rom[ 6259]='h00000000;
    rd_cycle[ 6260] = 1'b0;  wr_cycle[ 6260] = 1'b1;  addr_rom[ 6260]='h00003578;  wr_data_rom[ 6260]='h00003732;
    rd_cycle[ 6261] = 1'b1;  wr_cycle[ 6261] = 1'b0;  addr_rom[ 6261]='h00001b3c;  wr_data_rom[ 6261]='h00000000;
    rd_cycle[ 6262] = 1'b1;  wr_cycle[ 6262] = 1'b0;  addr_rom[ 6262]='h000020a0;  wr_data_rom[ 6262]='h00000000;
    rd_cycle[ 6263] = 1'b0;  wr_cycle[ 6263] = 1'b1;  addr_rom[ 6263]='h0000178c;  wr_data_rom[ 6263]='h00002a3b;
    rd_cycle[ 6264] = 1'b0;  wr_cycle[ 6264] = 1'b1;  addr_rom[ 6264]='h00000f3c;  wr_data_rom[ 6264]='h000021e0;
    rd_cycle[ 6265] = 1'b1;  wr_cycle[ 6265] = 1'b0;  addr_rom[ 6265]='h00001198;  wr_data_rom[ 6265]='h00000000;
    rd_cycle[ 6266] = 1'b0;  wr_cycle[ 6266] = 1'b1;  addr_rom[ 6266]='h00000db0;  wr_data_rom[ 6266]='h0000387f;
    rd_cycle[ 6267] = 1'b1;  wr_cycle[ 6267] = 1'b0;  addr_rom[ 6267]='h00000594;  wr_data_rom[ 6267]='h00000000;
    rd_cycle[ 6268] = 1'b0;  wr_cycle[ 6268] = 1'b1;  addr_rom[ 6268]='h000002d0;  wr_data_rom[ 6268]='h00001bde;
    rd_cycle[ 6269] = 1'b1;  wr_cycle[ 6269] = 1'b0;  addr_rom[ 6269]='h00000a64;  wr_data_rom[ 6269]='h00000000;
    rd_cycle[ 6270] = 1'b1;  wr_cycle[ 6270] = 1'b0;  addr_rom[ 6270]='h00000af0;  wr_data_rom[ 6270]='h00000000;
    rd_cycle[ 6271] = 1'b0;  wr_cycle[ 6271] = 1'b1;  addr_rom[ 6271]='h00001c70;  wr_data_rom[ 6271]='h00001f73;
    rd_cycle[ 6272] = 1'b0;  wr_cycle[ 6272] = 1'b1;  addr_rom[ 6272]='h00001c54;  wr_data_rom[ 6272]='h00003f08;
    rd_cycle[ 6273] = 1'b0;  wr_cycle[ 6273] = 1'b1;  addr_rom[ 6273]='h00002b20;  wr_data_rom[ 6273]='h0000131b;
    rd_cycle[ 6274] = 1'b0;  wr_cycle[ 6274] = 1'b1;  addr_rom[ 6274]='h00002160;  wr_data_rom[ 6274]='h0000101e;
    rd_cycle[ 6275] = 1'b1;  wr_cycle[ 6275] = 1'b0;  addr_rom[ 6275]='h000034c8;  wr_data_rom[ 6275]='h00000000;
    rd_cycle[ 6276] = 1'b1;  wr_cycle[ 6276] = 1'b0;  addr_rom[ 6276]='h000034cc;  wr_data_rom[ 6276]='h00000000;
    rd_cycle[ 6277] = 1'b1;  wr_cycle[ 6277] = 1'b0;  addr_rom[ 6277]='h00002e90;  wr_data_rom[ 6277]='h00000000;
    rd_cycle[ 6278] = 1'b1;  wr_cycle[ 6278] = 1'b0;  addr_rom[ 6278]='h00000830;  wr_data_rom[ 6278]='h00000000;
    rd_cycle[ 6279] = 1'b1;  wr_cycle[ 6279] = 1'b0;  addr_rom[ 6279]='h000029f4;  wr_data_rom[ 6279]='h00000000;
    rd_cycle[ 6280] = 1'b1;  wr_cycle[ 6280] = 1'b0;  addr_rom[ 6280]='h0000174c;  wr_data_rom[ 6280]='h00000000;
    rd_cycle[ 6281] = 1'b1;  wr_cycle[ 6281] = 1'b0;  addr_rom[ 6281]='h00003704;  wr_data_rom[ 6281]='h00000000;
    rd_cycle[ 6282] = 1'b0;  wr_cycle[ 6282] = 1'b1;  addr_rom[ 6282]='h00003728;  wr_data_rom[ 6282]='h00003af4;
    rd_cycle[ 6283] = 1'b1;  wr_cycle[ 6283] = 1'b0;  addr_rom[ 6283]='h00000680;  wr_data_rom[ 6283]='h00000000;
    rd_cycle[ 6284] = 1'b1;  wr_cycle[ 6284] = 1'b0;  addr_rom[ 6284]='h00001558;  wr_data_rom[ 6284]='h00000000;
    rd_cycle[ 6285] = 1'b0;  wr_cycle[ 6285] = 1'b1;  addr_rom[ 6285]='h000007d0;  wr_data_rom[ 6285]='h00003528;
    rd_cycle[ 6286] = 1'b1;  wr_cycle[ 6286] = 1'b0;  addr_rom[ 6286]='h000026c8;  wr_data_rom[ 6286]='h00000000;
    rd_cycle[ 6287] = 1'b0;  wr_cycle[ 6287] = 1'b1;  addr_rom[ 6287]='h000024d8;  wr_data_rom[ 6287]='h00003a1e;
    rd_cycle[ 6288] = 1'b0;  wr_cycle[ 6288] = 1'b1;  addr_rom[ 6288]='h000025f8;  wr_data_rom[ 6288]='h000038d5;
    rd_cycle[ 6289] = 1'b0;  wr_cycle[ 6289] = 1'b1;  addr_rom[ 6289]='h00001d30;  wr_data_rom[ 6289]='h00002c16;
    rd_cycle[ 6290] = 1'b1;  wr_cycle[ 6290] = 1'b0;  addr_rom[ 6290]='h00001f30;  wr_data_rom[ 6290]='h00000000;
    rd_cycle[ 6291] = 1'b1;  wr_cycle[ 6291] = 1'b0;  addr_rom[ 6291]='h00000540;  wr_data_rom[ 6291]='h00000000;
    rd_cycle[ 6292] = 1'b1;  wr_cycle[ 6292] = 1'b0;  addr_rom[ 6292]='h00002e48;  wr_data_rom[ 6292]='h00000000;
    rd_cycle[ 6293] = 1'b0;  wr_cycle[ 6293] = 1'b1;  addr_rom[ 6293]='h00003fc0;  wr_data_rom[ 6293]='h00003ed6;
    rd_cycle[ 6294] = 1'b0;  wr_cycle[ 6294] = 1'b1;  addr_rom[ 6294]='h00000564;  wr_data_rom[ 6294]='h0000257e;
    rd_cycle[ 6295] = 1'b1;  wr_cycle[ 6295] = 1'b0;  addr_rom[ 6295]='h00003114;  wr_data_rom[ 6295]='h00000000;
    rd_cycle[ 6296] = 1'b1;  wr_cycle[ 6296] = 1'b0;  addr_rom[ 6296]='h00002be8;  wr_data_rom[ 6296]='h00000000;
    rd_cycle[ 6297] = 1'b0;  wr_cycle[ 6297] = 1'b1;  addr_rom[ 6297]='h00003ad4;  wr_data_rom[ 6297]='h000022f2;
    rd_cycle[ 6298] = 1'b0;  wr_cycle[ 6298] = 1'b1;  addr_rom[ 6298]='h000018f4;  wr_data_rom[ 6298]='h000019fa;
    rd_cycle[ 6299] = 1'b1;  wr_cycle[ 6299] = 1'b0;  addr_rom[ 6299]='h00000340;  wr_data_rom[ 6299]='h00000000;
    rd_cycle[ 6300] = 1'b1;  wr_cycle[ 6300] = 1'b0;  addr_rom[ 6300]='h00000214;  wr_data_rom[ 6300]='h00000000;
    rd_cycle[ 6301] = 1'b1;  wr_cycle[ 6301] = 1'b0;  addr_rom[ 6301]='h0000048c;  wr_data_rom[ 6301]='h00000000;
    rd_cycle[ 6302] = 1'b1;  wr_cycle[ 6302] = 1'b0;  addr_rom[ 6302]='h0000266c;  wr_data_rom[ 6302]='h00000000;
    rd_cycle[ 6303] = 1'b0;  wr_cycle[ 6303] = 1'b1;  addr_rom[ 6303]='h00002568;  wr_data_rom[ 6303]='h00001229;
    rd_cycle[ 6304] = 1'b0;  wr_cycle[ 6304] = 1'b1;  addr_rom[ 6304]='h000011cc;  wr_data_rom[ 6304]='h00002538;
    rd_cycle[ 6305] = 1'b1;  wr_cycle[ 6305] = 1'b0;  addr_rom[ 6305]='h00000474;  wr_data_rom[ 6305]='h00000000;
    rd_cycle[ 6306] = 1'b1;  wr_cycle[ 6306] = 1'b0;  addr_rom[ 6306]='h00002060;  wr_data_rom[ 6306]='h00000000;
    rd_cycle[ 6307] = 1'b1;  wr_cycle[ 6307] = 1'b0;  addr_rom[ 6307]='h00000f30;  wr_data_rom[ 6307]='h00000000;
    rd_cycle[ 6308] = 1'b1;  wr_cycle[ 6308] = 1'b0;  addr_rom[ 6308]='h00002cbc;  wr_data_rom[ 6308]='h00000000;
    rd_cycle[ 6309] = 1'b1;  wr_cycle[ 6309] = 1'b0;  addr_rom[ 6309]='h00003ff8;  wr_data_rom[ 6309]='h00000000;
    rd_cycle[ 6310] = 1'b1;  wr_cycle[ 6310] = 1'b0;  addr_rom[ 6310]='h000000c4;  wr_data_rom[ 6310]='h00000000;
    rd_cycle[ 6311] = 1'b0;  wr_cycle[ 6311] = 1'b1;  addr_rom[ 6311]='h00003d80;  wr_data_rom[ 6311]='h00003c73;
    rd_cycle[ 6312] = 1'b1;  wr_cycle[ 6312] = 1'b0;  addr_rom[ 6312]='h0000112c;  wr_data_rom[ 6312]='h00000000;
    rd_cycle[ 6313] = 1'b0;  wr_cycle[ 6313] = 1'b1;  addr_rom[ 6313]='h00003464;  wr_data_rom[ 6313]='h00003c9f;
    rd_cycle[ 6314] = 1'b1;  wr_cycle[ 6314] = 1'b0;  addr_rom[ 6314]='h00001744;  wr_data_rom[ 6314]='h00000000;
    rd_cycle[ 6315] = 1'b1;  wr_cycle[ 6315] = 1'b0;  addr_rom[ 6315]='h00002bc8;  wr_data_rom[ 6315]='h00000000;
    rd_cycle[ 6316] = 1'b0;  wr_cycle[ 6316] = 1'b1;  addr_rom[ 6316]='h000029dc;  wr_data_rom[ 6316]='h000028cb;
    rd_cycle[ 6317] = 1'b0;  wr_cycle[ 6317] = 1'b1;  addr_rom[ 6317]='h00001528;  wr_data_rom[ 6317]='h00002ed4;
    rd_cycle[ 6318] = 1'b1;  wr_cycle[ 6318] = 1'b0;  addr_rom[ 6318]='h00003170;  wr_data_rom[ 6318]='h00000000;
    rd_cycle[ 6319] = 1'b0;  wr_cycle[ 6319] = 1'b1;  addr_rom[ 6319]='h00002728;  wr_data_rom[ 6319]='h00000081;
    rd_cycle[ 6320] = 1'b1;  wr_cycle[ 6320] = 1'b0;  addr_rom[ 6320]='h0000320c;  wr_data_rom[ 6320]='h00000000;
    rd_cycle[ 6321] = 1'b1;  wr_cycle[ 6321] = 1'b0;  addr_rom[ 6321]='h00003974;  wr_data_rom[ 6321]='h00000000;
    rd_cycle[ 6322] = 1'b1;  wr_cycle[ 6322] = 1'b0;  addr_rom[ 6322]='h0000239c;  wr_data_rom[ 6322]='h00000000;
    rd_cycle[ 6323] = 1'b0;  wr_cycle[ 6323] = 1'b1;  addr_rom[ 6323]='h00001178;  wr_data_rom[ 6323]='h00003e02;
    rd_cycle[ 6324] = 1'b0;  wr_cycle[ 6324] = 1'b1;  addr_rom[ 6324]='h000007a4;  wr_data_rom[ 6324]='h00000567;
    rd_cycle[ 6325] = 1'b0;  wr_cycle[ 6325] = 1'b1;  addr_rom[ 6325]='h00000a74;  wr_data_rom[ 6325]='h0000175c;
    rd_cycle[ 6326] = 1'b1;  wr_cycle[ 6326] = 1'b0;  addr_rom[ 6326]='h000005fc;  wr_data_rom[ 6326]='h00000000;
    rd_cycle[ 6327] = 1'b0;  wr_cycle[ 6327] = 1'b1;  addr_rom[ 6327]='h00002ecc;  wr_data_rom[ 6327]='h00002bde;
    rd_cycle[ 6328] = 1'b0;  wr_cycle[ 6328] = 1'b1;  addr_rom[ 6328]='h00002cd4;  wr_data_rom[ 6328]='h00002197;
    rd_cycle[ 6329] = 1'b1;  wr_cycle[ 6329] = 1'b0;  addr_rom[ 6329]='h00003b64;  wr_data_rom[ 6329]='h00000000;
    rd_cycle[ 6330] = 1'b0;  wr_cycle[ 6330] = 1'b1;  addr_rom[ 6330]='h00001d54;  wr_data_rom[ 6330]='h00003f65;
    rd_cycle[ 6331] = 1'b0;  wr_cycle[ 6331] = 1'b1;  addr_rom[ 6331]='h00003a88;  wr_data_rom[ 6331]='h00003f35;
    rd_cycle[ 6332] = 1'b1;  wr_cycle[ 6332] = 1'b0;  addr_rom[ 6332]='h00002ff0;  wr_data_rom[ 6332]='h00000000;
    rd_cycle[ 6333] = 1'b0;  wr_cycle[ 6333] = 1'b1;  addr_rom[ 6333]='h000038d8;  wr_data_rom[ 6333]='h00002b38;
    rd_cycle[ 6334] = 1'b0;  wr_cycle[ 6334] = 1'b1;  addr_rom[ 6334]='h00003584;  wr_data_rom[ 6334]='h00002100;
    rd_cycle[ 6335] = 1'b1;  wr_cycle[ 6335] = 1'b0;  addr_rom[ 6335]='h00003344;  wr_data_rom[ 6335]='h00000000;
    rd_cycle[ 6336] = 1'b0;  wr_cycle[ 6336] = 1'b1;  addr_rom[ 6336]='h000017a0;  wr_data_rom[ 6336]='h00003f83;
    rd_cycle[ 6337] = 1'b0;  wr_cycle[ 6337] = 1'b1;  addr_rom[ 6337]='h00001044;  wr_data_rom[ 6337]='h00003259;
    rd_cycle[ 6338] = 1'b0;  wr_cycle[ 6338] = 1'b1;  addr_rom[ 6338]='h000038dc;  wr_data_rom[ 6338]='h000022de;
    rd_cycle[ 6339] = 1'b1;  wr_cycle[ 6339] = 1'b0;  addr_rom[ 6339]='h00003b2c;  wr_data_rom[ 6339]='h00000000;
    rd_cycle[ 6340] = 1'b0;  wr_cycle[ 6340] = 1'b1;  addr_rom[ 6340]='h000038f8;  wr_data_rom[ 6340]='h00002428;
    rd_cycle[ 6341] = 1'b1;  wr_cycle[ 6341] = 1'b0;  addr_rom[ 6341]='h00002f78;  wr_data_rom[ 6341]='h00000000;
    rd_cycle[ 6342] = 1'b0;  wr_cycle[ 6342] = 1'b1;  addr_rom[ 6342]='h00002968;  wr_data_rom[ 6342]='h0000036e;
    rd_cycle[ 6343] = 1'b0;  wr_cycle[ 6343] = 1'b1;  addr_rom[ 6343]='h000002c8;  wr_data_rom[ 6343]='h00000865;
    rd_cycle[ 6344] = 1'b0;  wr_cycle[ 6344] = 1'b1;  addr_rom[ 6344]='h00003a54;  wr_data_rom[ 6344]='h00001f93;
    rd_cycle[ 6345] = 1'b1;  wr_cycle[ 6345] = 1'b0;  addr_rom[ 6345]='h00001898;  wr_data_rom[ 6345]='h00000000;
    rd_cycle[ 6346] = 1'b1;  wr_cycle[ 6346] = 1'b0;  addr_rom[ 6346]='h00001ff8;  wr_data_rom[ 6346]='h00000000;
    rd_cycle[ 6347] = 1'b0;  wr_cycle[ 6347] = 1'b1;  addr_rom[ 6347]='h000035dc;  wr_data_rom[ 6347]='h00003d2e;
    rd_cycle[ 6348] = 1'b0;  wr_cycle[ 6348] = 1'b1;  addr_rom[ 6348]='h00002918;  wr_data_rom[ 6348]='h000008b6;
    rd_cycle[ 6349] = 1'b0;  wr_cycle[ 6349] = 1'b1;  addr_rom[ 6349]='h00003098;  wr_data_rom[ 6349]='h00002df6;
    rd_cycle[ 6350] = 1'b0;  wr_cycle[ 6350] = 1'b1;  addr_rom[ 6350]='h00001dc4;  wr_data_rom[ 6350]='h00003382;
    rd_cycle[ 6351] = 1'b1;  wr_cycle[ 6351] = 1'b0;  addr_rom[ 6351]='h00003c54;  wr_data_rom[ 6351]='h00000000;
    rd_cycle[ 6352] = 1'b0;  wr_cycle[ 6352] = 1'b1;  addr_rom[ 6352]='h000013f8;  wr_data_rom[ 6352]='h00002e56;
    rd_cycle[ 6353] = 1'b0;  wr_cycle[ 6353] = 1'b1;  addr_rom[ 6353]='h000008dc;  wr_data_rom[ 6353]='h000024fb;
    rd_cycle[ 6354] = 1'b1;  wr_cycle[ 6354] = 1'b0;  addr_rom[ 6354]='h00002bd0;  wr_data_rom[ 6354]='h00000000;
    rd_cycle[ 6355] = 1'b0;  wr_cycle[ 6355] = 1'b1;  addr_rom[ 6355]='h00003b68;  wr_data_rom[ 6355]='h00000226;
    rd_cycle[ 6356] = 1'b1;  wr_cycle[ 6356] = 1'b0;  addr_rom[ 6356]='h000006a4;  wr_data_rom[ 6356]='h00000000;
    rd_cycle[ 6357] = 1'b1;  wr_cycle[ 6357] = 1'b0;  addr_rom[ 6357]='h0000038c;  wr_data_rom[ 6357]='h00000000;
    rd_cycle[ 6358] = 1'b1;  wr_cycle[ 6358] = 1'b0;  addr_rom[ 6358]='h00003ff4;  wr_data_rom[ 6358]='h00000000;
    rd_cycle[ 6359] = 1'b0;  wr_cycle[ 6359] = 1'b1;  addr_rom[ 6359]='h00002d80;  wr_data_rom[ 6359]='h00003a2e;
    rd_cycle[ 6360] = 1'b0;  wr_cycle[ 6360] = 1'b1;  addr_rom[ 6360]='h00003ffc;  wr_data_rom[ 6360]='h000023f0;
    rd_cycle[ 6361] = 1'b0;  wr_cycle[ 6361] = 1'b1;  addr_rom[ 6361]='h000011a0;  wr_data_rom[ 6361]='h000028a8;
    rd_cycle[ 6362] = 1'b1;  wr_cycle[ 6362] = 1'b0;  addr_rom[ 6362]='h000036cc;  wr_data_rom[ 6362]='h00000000;
    rd_cycle[ 6363] = 1'b1;  wr_cycle[ 6363] = 1'b0;  addr_rom[ 6363]='h00002c2c;  wr_data_rom[ 6363]='h00000000;
    rd_cycle[ 6364] = 1'b0;  wr_cycle[ 6364] = 1'b1;  addr_rom[ 6364]='h00002b70;  wr_data_rom[ 6364]='h00003b32;
    rd_cycle[ 6365] = 1'b0;  wr_cycle[ 6365] = 1'b1;  addr_rom[ 6365]='h000014e0;  wr_data_rom[ 6365]='h00003854;
    rd_cycle[ 6366] = 1'b0;  wr_cycle[ 6366] = 1'b1;  addr_rom[ 6366]='h000025f4;  wr_data_rom[ 6366]='h00000278;
    rd_cycle[ 6367] = 1'b1;  wr_cycle[ 6367] = 1'b0;  addr_rom[ 6367]='h0000134c;  wr_data_rom[ 6367]='h00000000;
    rd_cycle[ 6368] = 1'b0;  wr_cycle[ 6368] = 1'b1;  addr_rom[ 6368]='h00002f78;  wr_data_rom[ 6368]='h000001e0;
    rd_cycle[ 6369] = 1'b0;  wr_cycle[ 6369] = 1'b1;  addr_rom[ 6369]='h000005b4;  wr_data_rom[ 6369]='h00002301;
    rd_cycle[ 6370] = 1'b0;  wr_cycle[ 6370] = 1'b1;  addr_rom[ 6370]='h000003a0;  wr_data_rom[ 6370]='h00002bc1;
    rd_cycle[ 6371] = 1'b1;  wr_cycle[ 6371] = 1'b0;  addr_rom[ 6371]='h00002490;  wr_data_rom[ 6371]='h00000000;
    rd_cycle[ 6372] = 1'b1;  wr_cycle[ 6372] = 1'b0;  addr_rom[ 6372]='h00002b6c;  wr_data_rom[ 6372]='h00000000;
    rd_cycle[ 6373] = 1'b0;  wr_cycle[ 6373] = 1'b1;  addr_rom[ 6373]='h00003a80;  wr_data_rom[ 6373]='h00003877;
    rd_cycle[ 6374] = 1'b1;  wr_cycle[ 6374] = 1'b0;  addr_rom[ 6374]='h000006d8;  wr_data_rom[ 6374]='h00000000;
    rd_cycle[ 6375] = 1'b0;  wr_cycle[ 6375] = 1'b1;  addr_rom[ 6375]='h00001590;  wr_data_rom[ 6375]='h00002ba3;
    rd_cycle[ 6376] = 1'b1;  wr_cycle[ 6376] = 1'b0;  addr_rom[ 6376]='h000005cc;  wr_data_rom[ 6376]='h00000000;
    rd_cycle[ 6377] = 1'b1;  wr_cycle[ 6377] = 1'b0;  addr_rom[ 6377]='h000033c0;  wr_data_rom[ 6377]='h00000000;
    rd_cycle[ 6378] = 1'b1;  wr_cycle[ 6378] = 1'b0;  addr_rom[ 6378]='h000010a4;  wr_data_rom[ 6378]='h00000000;
    rd_cycle[ 6379] = 1'b1;  wr_cycle[ 6379] = 1'b0;  addr_rom[ 6379]='h00002c98;  wr_data_rom[ 6379]='h00000000;
    rd_cycle[ 6380] = 1'b1;  wr_cycle[ 6380] = 1'b0;  addr_rom[ 6380]='h00002954;  wr_data_rom[ 6380]='h00000000;
    rd_cycle[ 6381] = 1'b0;  wr_cycle[ 6381] = 1'b1;  addr_rom[ 6381]='h000009e8;  wr_data_rom[ 6381]='h0000108d;
    rd_cycle[ 6382] = 1'b1;  wr_cycle[ 6382] = 1'b0;  addr_rom[ 6382]='h00000bf0;  wr_data_rom[ 6382]='h00000000;
    rd_cycle[ 6383] = 1'b0;  wr_cycle[ 6383] = 1'b1;  addr_rom[ 6383]='h00001d50;  wr_data_rom[ 6383]='h000001d0;
    rd_cycle[ 6384] = 1'b0;  wr_cycle[ 6384] = 1'b1;  addr_rom[ 6384]='h00000b28;  wr_data_rom[ 6384]='h000022a9;
    rd_cycle[ 6385] = 1'b1;  wr_cycle[ 6385] = 1'b0;  addr_rom[ 6385]='h000018c8;  wr_data_rom[ 6385]='h00000000;
    rd_cycle[ 6386] = 1'b0;  wr_cycle[ 6386] = 1'b1;  addr_rom[ 6386]='h00000e98;  wr_data_rom[ 6386]='h00002f3d;
    rd_cycle[ 6387] = 1'b0;  wr_cycle[ 6387] = 1'b1;  addr_rom[ 6387]='h0000052c;  wr_data_rom[ 6387]='h00000bab;
    rd_cycle[ 6388] = 1'b1;  wr_cycle[ 6388] = 1'b0;  addr_rom[ 6388]='h00002620;  wr_data_rom[ 6388]='h00000000;
    rd_cycle[ 6389] = 1'b0;  wr_cycle[ 6389] = 1'b1;  addr_rom[ 6389]='h00002df0;  wr_data_rom[ 6389]='h00002ed8;
    rd_cycle[ 6390] = 1'b0;  wr_cycle[ 6390] = 1'b1;  addr_rom[ 6390]='h000018a8;  wr_data_rom[ 6390]='h0000394a;
    rd_cycle[ 6391] = 1'b1;  wr_cycle[ 6391] = 1'b0;  addr_rom[ 6391]='h00000334;  wr_data_rom[ 6391]='h00000000;
    rd_cycle[ 6392] = 1'b0;  wr_cycle[ 6392] = 1'b1;  addr_rom[ 6392]='h00000fec;  wr_data_rom[ 6392]='h000038a0;
    rd_cycle[ 6393] = 1'b0;  wr_cycle[ 6393] = 1'b1;  addr_rom[ 6393]='h00000884;  wr_data_rom[ 6393]='h00001398;
    rd_cycle[ 6394] = 1'b1;  wr_cycle[ 6394] = 1'b0;  addr_rom[ 6394]='h0000357c;  wr_data_rom[ 6394]='h00000000;
    rd_cycle[ 6395] = 1'b0;  wr_cycle[ 6395] = 1'b1;  addr_rom[ 6395]='h00001a50;  wr_data_rom[ 6395]='h0000097c;
    rd_cycle[ 6396] = 1'b1;  wr_cycle[ 6396] = 1'b0;  addr_rom[ 6396]='h00003364;  wr_data_rom[ 6396]='h00000000;
    rd_cycle[ 6397] = 1'b0;  wr_cycle[ 6397] = 1'b1;  addr_rom[ 6397]='h000011d8;  wr_data_rom[ 6397]='h00002afc;
    rd_cycle[ 6398] = 1'b0;  wr_cycle[ 6398] = 1'b1;  addr_rom[ 6398]='h00001560;  wr_data_rom[ 6398]='h00003eaf;
    rd_cycle[ 6399] = 1'b0;  wr_cycle[ 6399] = 1'b1;  addr_rom[ 6399]='h00001f20;  wr_data_rom[ 6399]='h0000149e;
    rd_cycle[ 6400] = 1'b0;  wr_cycle[ 6400] = 1'b1;  addr_rom[ 6400]='h00002f08;  wr_data_rom[ 6400]='h00001a3c;
    rd_cycle[ 6401] = 1'b1;  wr_cycle[ 6401] = 1'b0;  addr_rom[ 6401]='h00000014;  wr_data_rom[ 6401]='h00000000;
    rd_cycle[ 6402] = 1'b1;  wr_cycle[ 6402] = 1'b0;  addr_rom[ 6402]='h000004a4;  wr_data_rom[ 6402]='h00000000;
    rd_cycle[ 6403] = 1'b1;  wr_cycle[ 6403] = 1'b0;  addr_rom[ 6403]='h00002930;  wr_data_rom[ 6403]='h00000000;
    rd_cycle[ 6404] = 1'b0;  wr_cycle[ 6404] = 1'b1;  addr_rom[ 6404]='h00002e20;  wr_data_rom[ 6404]='h000022f1;
    rd_cycle[ 6405] = 1'b1;  wr_cycle[ 6405] = 1'b0;  addr_rom[ 6405]='h00001050;  wr_data_rom[ 6405]='h00000000;
    rd_cycle[ 6406] = 1'b0;  wr_cycle[ 6406] = 1'b1;  addr_rom[ 6406]='h00001c20;  wr_data_rom[ 6406]='h00000e59;
    rd_cycle[ 6407] = 1'b1;  wr_cycle[ 6407] = 1'b0;  addr_rom[ 6407]='h00003d88;  wr_data_rom[ 6407]='h00000000;
    rd_cycle[ 6408] = 1'b0;  wr_cycle[ 6408] = 1'b1;  addr_rom[ 6408]='h000039f8;  wr_data_rom[ 6408]='h000019fa;
    rd_cycle[ 6409] = 1'b0;  wr_cycle[ 6409] = 1'b1;  addr_rom[ 6409]='h00001350;  wr_data_rom[ 6409]='h00002167;
    rd_cycle[ 6410] = 1'b1;  wr_cycle[ 6410] = 1'b0;  addr_rom[ 6410]='h00000d54;  wr_data_rom[ 6410]='h00000000;
    rd_cycle[ 6411] = 1'b1;  wr_cycle[ 6411] = 1'b0;  addr_rom[ 6411]='h000037a4;  wr_data_rom[ 6411]='h00000000;
    rd_cycle[ 6412] = 1'b0;  wr_cycle[ 6412] = 1'b1;  addr_rom[ 6412]='h000035e0;  wr_data_rom[ 6412]='h00002fcb;
    rd_cycle[ 6413] = 1'b1;  wr_cycle[ 6413] = 1'b0;  addr_rom[ 6413]='h00002854;  wr_data_rom[ 6413]='h00000000;
    rd_cycle[ 6414] = 1'b1;  wr_cycle[ 6414] = 1'b0;  addr_rom[ 6414]='h000003dc;  wr_data_rom[ 6414]='h00000000;
    rd_cycle[ 6415] = 1'b1;  wr_cycle[ 6415] = 1'b0;  addr_rom[ 6415]='h0000350c;  wr_data_rom[ 6415]='h00000000;
    rd_cycle[ 6416] = 1'b1;  wr_cycle[ 6416] = 1'b0;  addr_rom[ 6416]='h00002fd4;  wr_data_rom[ 6416]='h00000000;
    rd_cycle[ 6417] = 1'b1;  wr_cycle[ 6417] = 1'b0;  addr_rom[ 6417]='h000037b8;  wr_data_rom[ 6417]='h00000000;
    rd_cycle[ 6418] = 1'b0;  wr_cycle[ 6418] = 1'b1;  addr_rom[ 6418]='h000017a4;  wr_data_rom[ 6418]='h00003a51;
    rd_cycle[ 6419] = 1'b1;  wr_cycle[ 6419] = 1'b0;  addr_rom[ 6419]='h000039b4;  wr_data_rom[ 6419]='h00000000;
    rd_cycle[ 6420] = 1'b1;  wr_cycle[ 6420] = 1'b0;  addr_rom[ 6420]='h0000106c;  wr_data_rom[ 6420]='h00000000;
    rd_cycle[ 6421] = 1'b1;  wr_cycle[ 6421] = 1'b0;  addr_rom[ 6421]='h000011b0;  wr_data_rom[ 6421]='h00000000;
    rd_cycle[ 6422] = 1'b0;  wr_cycle[ 6422] = 1'b1;  addr_rom[ 6422]='h00001fb0;  wr_data_rom[ 6422]='h00003868;
    rd_cycle[ 6423] = 1'b0;  wr_cycle[ 6423] = 1'b1;  addr_rom[ 6423]='h00002930;  wr_data_rom[ 6423]='h00001700;
    rd_cycle[ 6424] = 1'b1;  wr_cycle[ 6424] = 1'b0;  addr_rom[ 6424]='h00002940;  wr_data_rom[ 6424]='h00000000;
    rd_cycle[ 6425] = 1'b1;  wr_cycle[ 6425] = 1'b0;  addr_rom[ 6425]='h00000594;  wr_data_rom[ 6425]='h00000000;
    rd_cycle[ 6426] = 1'b1;  wr_cycle[ 6426] = 1'b0;  addr_rom[ 6426]='h00003654;  wr_data_rom[ 6426]='h00000000;
    rd_cycle[ 6427] = 1'b1;  wr_cycle[ 6427] = 1'b0;  addr_rom[ 6427]='h00001624;  wr_data_rom[ 6427]='h00000000;
    rd_cycle[ 6428] = 1'b0;  wr_cycle[ 6428] = 1'b1;  addr_rom[ 6428]='h000035d8;  wr_data_rom[ 6428]='h0000227b;
    rd_cycle[ 6429] = 1'b0;  wr_cycle[ 6429] = 1'b1;  addr_rom[ 6429]='h00000f44;  wr_data_rom[ 6429]='h00000b83;
    rd_cycle[ 6430] = 1'b1;  wr_cycle[ 6430] = 1'b0;  addr_rom[ 6430]='h000018f4;  wr_data_rom[ 6430]='h00000000;
    rd_cycle[ 6431] = 1'b1;  wr_cycle[ 6431] = 1'b0;  addr_rom[ 6431]='h00003ff0;  wr_data_rom[ 6431]='h00000000;
    rd_cycle[ 6432] = 1'b1;  wr_cycle[ 6432] = 1'b0;  addr_rom[ 6432]='h0000321c;  wr_data_rom[ 6432]='h00000000;
    rd_cycle[ 6433] = 1'b0;  wr_cycle[ 6433] = 1'b1;  addr_rom[ 6433]='h00002b10;  wr_data_rom[ 6433]='h00001ee2;
    rd_cycle[ 6434] = 1'b0;  wr_cycle[ 6434] = 1'b1;  addr_rom[ 6434]='h00000688;  wr_data_rom[ 6434]='h00001656;
    rd_cycle[ 6435] = 1'b0;  wr_cycle[ 6435] = 1'b1;  addr_rom[ 6435]='h00002e78;  wr_data_rom[ 6435]='h00002815;
    rd_cycle[ 6436] = 1'b1;  wr_cycle[ 6436] = 1'b0;  addr_rom[ 6436]='h00000a28;  wr_data_rom[ 6436]='h00000000;
    rd_cycle[ 6437] = 1'b0;  wr_cycle[ 6437] = 1'b1;  addr_rom[ 6437]='h00003e8c;  wr_data_rom[ 6437]='h00002486;
    rd_cycle[ 6438] = 1'b1;  wr_cycle[ 6438] = 1'b0;  addr_rom[ 6438]='h00002a88;  wr_data_rom[ 6438]='h00000000;
    rd_cycle[ 6439] = 1'b0;  wr_cycle[ 6439] = 1'b1;  addr_rom[ 6439]='h00003134;  wr_data_rom[ 6439]='h00001622;
    rd_cycle[ 6440] = 1'b1;  wr_cycle[ 6440] = 1'b0;  addr_rom[ 6440]='h00002efc;  wr_data_rom[ 6440]='h00000000;
    rd_cycle[ 6441] = 1'b1;  wr_cycle[ 6441] = 1'b0;  addr_rom[ 6441]='h00001c14;  wr_data_rom[ 6441]='h00000000;
    rd_cycle[ 6442] = 1'b1;  wr_cycle[ 6442] = 1'b0;  addr_rom[ 6442]='h00003a64;  wr_data_rom[ 6442]='h00000000;
    rd_cycle[ 6443] = 1'b1;  wr_cycle[ 6443] = 1'b0;  addr_rom[ 6443]='h000020ec;  wr_data_rom[ 6443]='h00000000;
    rd_cycle[ 6444] = 1'b1;  wr_cycle[ 6444] = 1'b0;  addr_rom[ 6444]='h00001a08;  wr_data_rom[ 6444]='h00000000;
    rd_cycle[ 6445] = 1'b0;  wr_cycle[ 6445] = 1'b1;  addr_rom[ 6445]='h0000369c;  wr_data_rom[ 6445]='h0000234b;
    rd_cycle[ 6446] = 1'b0;  wr_cycle[ 6446] = 1'b1;  addr_rom[ 6446]='h00002104;  wr_data_rom[ 6446]='h000007c9;
    rd_cycle[ 6447] = 1'b0;  wr_cycle[ 6447] = 1'b1;  addr_rom[ 6447]='h00003474;  wr_data_rom[ 6447]='h00002617;
    rd_cycle[ 6448] = 1'b1;  wr_cycle[ 6448] = 1'b0;  addr_rom[ 6448]='h000024c0;  wr_data_rom[ 6448]='h00000000;
    rd_cycle[ 6449] = 1'b0;  wr_cycle[ 6449] = 1'b1;  addr_rom[ 6449]='h00002ae4;  wr_data_rom[ 6449]='h000022a4;
    rd_cycle[ 6450] = 1'b0;  wr_cycle[ 6450] = 1'b1;  addr_rom[ 6450]='h00002488;  wr_data_rom[ 6450]='h0000325e;
    rd_cycle[ 6451] = 1'b1;  wr_cycle[ 6451] = 1'b0;  addr_rom[ 6451]='h00001a7c;  wr_data_rom[ 6451]='h00000000;
    rd_cycle[ 6452] = 1'b0;  wr_cycle[ 6452] = 1'b1;  addr_rom[ 6452]='h00000a98;  wr_data_rom[ 6452]='h00001730;
    rd_cycle[ 6453] = 1'b1;  wr_cycle[ 6453] = 1'b0;  addr_rom[ 6453]='h00002bc0;  wr_data_rom[ 6453]='h00000000;
    rd_cycle[ 6454] = 1'b1;  wr_cycle[ 6454] = 1'b0;  addr_rom[ 6454]='h00001ea4;  wr_data_rom[ 6454]='h00000000;
    rd_cycle[ 6455] = 1'b0;  wr_cycle[ 6455] = 1'b1;  addr_rom[ 6455]='h00001d60;  wr_data_rom[ 6455]='h00002b0a;
    rd_cycle[ 6456] = 1'b1;  wr_cycle[ 6456] = 1'b0;  addr_rom[ 6456]='h00001f44;  wr_data_rom[ 6456]='h00000000;
    rd_cycle[ 6457] = 1'b1;  wr_cycle[ 6457] = 1'b0;  addr_rom[ 6457]='h000039f4;  wr_data_rom[ 6457]='h00000000;
    rd_cycle[ 6458] = 1'b0;  wr_cycle[ 6458] = 1'b1;  addr_rom[ 6458]='h00000ad0;  wr_data_rom[ 6458]='h00002702;
    rd_cycle[ 6459] = 1'b0;  wr_cycle[ 6459] = 1'b1;  addr_rom[ 6459]='h00003698;  wr_data_rom[ 6459]='h00003fa0;
    rd_cycle[ 6460] = 1'b0;  wr_cycle[ 6460] = 1'b1;  addr_rom[ 6460]='h00000664;  wr_data_rom[ 6460]='h00000212;
    rd_cycle[ 6461] = 1'b1;  wr_cycle[ 6461] = 1'b0;  addr_rom[ 6461]='h00003594;  wr_data_rom[ 6461]='h00000000;
    rd_cycle[ 6462] = 1'b1;  wr_cycle[ 6462] = 1'b0;  addr_rom[ 6462]='h00003b64;  wr_data_rom[ 6462]='h00000000;
    rd_cycle[ 6463] = 1'b0;  wr_cycle[ 6463] = 1'b1;  addr_rom[ 6463]='h00001ce8;  wr_data_rom[ 6463]='h00001572;
    rd_cycle[ 6464] = 1'b0;  wr_cycle[ 6464] = 1'b1;  addr_rom[ 6464]='h0000084c;  wr_data_rom[ 6464]='h000013c5;
    rd_cycle[ 6465] = 1'b0;  wr_cycle[ 6465] = 1'b1;  addr_rom[ 6465]='h000001ac;  wr_data_rom[ 6465]='h00003649;
    rd_cycle[ 6466] = 1'b0;  wr_cycle[ 6466] = 1'b1;  addr_rom[ 6466]='h00000a10;  wr_data_rom[ 6466]='h00000682;
    rd_cycle[ 6467] = 1'b1;  wr_cycle[ 6467] = 1'b0;  addr_rom[ 6467]='h00000ef0;  wr_data_rom[ 6467]='h00000000;
    rd_cycle[ 6468] = 1'b1;  wr_cycle[ 6468] = 1'b0;  addr_rom[ 6468]='h0000376c;  wr_data_rom[ 6468]='h00000000;
    rd_cycle[ 6469] = 1'b0;  wr_cycle[ 6469] = 1'b1;  addr_rom[ 6469]='h000016d8;  wr_data_rom[ 6469]='h0000193f;
    rd_cycle[ 6470] = 1'b1;  wr_cycle[ 6470] = 1'b0;  addr_rom[ 6470]='h000002a0;  wr_data_rom[ 6470]='h00000000;
    rd_cycle[ 6471] = 1'b1;  wr_cycle[ 6471] = 1'b0;  addr_rom[ 6471]='h000032b8;  wr_data_rom[ 6471]='h00000000;
    rd_cycle[ 6472] = 1'b1;  wr_cycle[ 6472] = 1'b0;  addr_rom[ 6472]='h000022dc;  wr_data_rom[ 6472]='h00000000;
    rd_cycle[ 6473] = 1'b1;  wr_cycle[ 6473] = 1'b0;  addr_rom[ 6473]='h00000f0c;  wr_data_rom[ 6473]='h00000000;
    rd_cycle[ 6474] = 1'b1;  wr_cycle[ 6474] = 1'b0;  addr_rom[ 6474]='h00001d50;  wr_data_rom[ 6474]='h00000000;
    rd_cycle[ 6475] = 1'b0;  wr_cycle[ 6475] = 1'b1;  addr_rom[ 6475]='h00003d54;  wr_data_rom[ 6475]='h000033fc;
    rd_cycle[ 6476] = 1'b0;  wr_cycle[ 6476] = 1'b1;  addr_rom[ 6476]='h00000664;  wr_data_rom[ 6476]='h00001673;
    rd_cycle[ 6477] = 1'b0;  wr_cycle[ 6477] = 1'b1;  addr_rom[ 6477]='h00000c78;  wr_data_rom[ 6477]='h000000c3;
    rd_cycle[ 6478] = 1'b0;  wr_cycle[ 6478] = 1'b1;  addr_rom[ 6478]='h0000229c;  wr_data_rom[ 6478]='h00003770;
    rd_cycle[ 6479] = 1'b0;  wr_cycle[ 6479] = 1'b1;  addr_rom[ 6479]='h00000160;  wr_data_rom[ 6479]='h00003cc7;
    rd_cycle[ 6480] = 1'b1;  wr_cycle[ 6480] = 1'b0;  addr_rom[ 6480]='h00001504;  wr_data_rom[ 6480]='h00000000;
    rd_cycle[ 6481] = 1'b1;  wr_cycle[ 6481] = 1'b0;  addr_rom[ 6481]='h00002304;  wr_data_rom[ 6481]='h00000000;
    rd_cycle[ 6482] = 1'b1;  wr_cycle[ 6482] = 1'b0;  addr_rom[ 6482]='h0000018c;  wr_data_rom[ 6482]='h00000000;
    rd_cycle[ 6483] = 1'b1;  wr_cycle[ 6483] = 1'b0;  addr_rom[ 6483]='h00001b80;  wr_data_rom[ 6483]='h00000000;
    rd_cycle[ 6484] = 1'b1;  wr_cycle[ 6484] = 1'b0;  addr_rom[ 6484]='h00001784;  wr_data_rom[ 6484]='h00000000;
    rd_cycle[ 6485] = 1'b0;  wr_cycle[ 6485] = 1'b1;  addr_rom[ 6485]='h00001430;  wr_data_rom[ 6485]='h000015fe;
    rd_cycle[ 6486] = 1'b1;  wr_cycle[ 6486] = 1'b0;  addr_rom[ 6486]='h00003140;  wr_data_rom[ 6486]='h00000000;
    rd_cycle[ 6487] = 1'b1;  wr_cycle[ 6487] = 1'b0;  addr_rom[ 6487]='h00003750;  wr_data_rom[ 6487]='h00000000;
    rd_cycle[ 6488] = 1'b0;  wr_cycle[ 6488] = 1'b1;  addr_rom[ 6488]='h000009b0;  wr_data_rom[ 6488]='h00003375;
    rd_cycle[ 6489] = 1'b0;  wr_cycle[ 6489] = 1'b1;  addr_rom[ 6489]='h000027c8;  wr_data_rom[ 6489]='h000007ff;
    rd_cycle[ 6490] = 1'b0;  wr_cycle[ 6490] = 1'b1;  addr_rom[ 6490]='h00001390;  wr_data_rom[ 6490]='h00001682;
    rd_cycle[ 6491] = 1'b0;  wr_cycle[ 6491] = 1'b1;  addr_rom[ 6491]='h00000344;  wr_data_rom[ 6491]='h00002165;
    rd_cycle[ 6492] = 1'b0;  wr_cycle[ 6492] = 1'b1;  addr_rom[ 6492]='h00000490;  wr_data_rom[ 6492]='h00001bd6;
    rd_cycle[ 6493] = 1'b0;  wr_cycle[ 6493] = 1'b1;  addr_rom[ 6493]='h000006f8;  wr_data_rom[ 6493]='h00002f82;
    rd_cycle[ 6494] = 1'b1;  wr_cycle[ 6494] = 1'b0;  addr_rom[ 6494]='h00000438;  wr_data_rom[ 6494]='h00000000;
    rd_cycle[ 6495] = 1'b1;  wr_cycle[ 6495] = 1'b0;  addr_rom[ 6495]='h000018cc;  wr_data_rom[ 6495]='h00000000;
    rd_cycle[ 6496] = 1'b1;  wr_cycle[ 6496] = 1'b0;  addr_rom[ 6496]='h00000c80;  wr_data_rom[ 6496]='h00000000;
    rd_cycle[ 6497] = 1'b1;  wr_cycle[ 6497] = 1'b0;  addr_rom[ 6497]='h00000868;  wr_data_rom[ 6497]='h00000000;
    rd_cycle[ 6498] = 1'b1;  wr_cycle[ 6498] = 1'b0;  addr_rom[ 6498]='h00003380;  wr_data_rom[ 6498]='h00000000;
    rd_cycle[ 6499] = 1'b1;  wr_cycle[ 6499] = 1'b0;  addr_rom[ 6499]='h00002cb8;  wr_data_rom[ 6499]='h00000000;
    rd_cycle[ 6500] = 1'b0;  wr_cycle[ 6500] = 1'b1;  addr_rom[ 6500]='h00001d80;  wr_data_rom[ 6500]='h00000a62;
    rd_cycle[ 6501] = 1'b0;  wr_cycle[ 6501] = 1'b1;  addr_rom[ 6501]='h00003528;  wr_data_rom[ 6501]='h000003a6;
    rd_cycle[ 6502] = 1'b0;  wr_cycle[ 6502] = 1'b1;  addr_rom[ 6502]='h00001318;  wr_data_rom[ 6502]='h000008fb;
    rd_cycle[ 6503] = 1'b0;  wr_cycle[ 6503] = 1'b1;  addr_rom[ 6503]='h00000c64;  wr_data_rom[ 6503]='h0000002c;
    rd_cycle[ 6504] = 1'b1;  wr_cycle[ 6504] = 1'b0;  addr_rom[ 6504]='h0000039c;  wr_data_rom[ 6504]='h00000000;
    rd_cycle[ 6505] = 1'b0;  wr_cycle[ 6505] = 1'b1;  addr_rom[ 6505]='h000036b0;  wr_data_rom[ 6505]='h00002dd6;
    rd_cycle[ 6506] = 1'b1;  wr_cycle[ 6506] = 1'b0;  addr_rom[ 6506]='h00003634;  wr_data_rom[ 6506]='h00000000;
    rd_cycle[ 6507] = 1'b0;  wr_cycle[ 6507] = 1'b1;  addr_rom[ 6507]='h00000ce4;  wr_data_rom[ 6507]='h00003ff8;
    rd_cycle[ 6508] = 1'b1;  wr_cycle[ 6508] = 1'b0;  addr_rom[ 6508]='h0000032c;  wr_data_rom[ 6508]='h00000000;
    rd_cycle[ 6509] = 1'b1;  wr_cycle[ 6509] = 1'b0;  addr_rom[ 6509]='h00001d50;  wr_data_rom[ 6509]='h00000000;
    rd_cycle[ 6510] = 1'b1;  wr_cycle[ 6510] = 1'b0;  addr_rom[ 6510]='h00002a4c;  wr_data_rom[ 6510]='h00000000;
    rd_cycle[ 6511] = 1'b1;  wr_cycle[ 6511] = 1'b0;  addr_rom[ 6511]='h000021a0;  wr_data_rom[ 6511]='h00000000;
    rd_cycle[ 6512] = 1'b1;  wr_cycle[ 6512] = 1'b0;  addr_rom[ 6512]='h000011ac;  wr_data_rom[ 6512]='h00000000;
    rd_cycle[ 6513] = 1'b0;  wr_cycle[ 6513] = 1'b1;  addr_rom[ 6513]='h00002ac4;  wr_data_rom[ 6513]='h0000182a;
    rd_cycle[ 6514] = 1'b1;  wr_cycle[ 6514] = 1'b0;  addr_rom[ 6514]='h000007c0;  wr_data_rom[ 6514]='h00000000;
    rd_cycle[ 6515] = 1'b1;  wr_cycle[ 6515] = 1'b0;  addr_rom[ 6515]='h00003804;  wr_data_rom[ 6515]='h00000000;
    rd_cycle[ 6516] = 1'b0;  wr_cycle[ 6516] = 1'b1;  addr_rom[ 6516]='h00003208;  wr_data_rom[ 6516]='h000010f3;
    rd_cycle[ 6517] = 1'b1;  wr_cycle[ 6517] = 1'b0;  addr_rom[ 6517]='h000024fc;  wr_data_rom[ 6517]='h00000000;
    rd_cycle[ 6518] = 1'b0;  wr_cycle[ 6518] = 1'b1;  addr_rom[ 6518]='h000038d0;  wr_data_rom[ 6518]='h000028a5;
    rd_cycle[ 6519] = 1'b1;  wr_cycle[ 6519] = 1'b0;  addr_rom[ 6519]='h00002ac0;  wr_data_rom[ 6519]='h00000000;
    rd_cycle[ 6520] = 1'b0;  wr_cycle[ 6520] = 1'b1;  addr_rom[ 6520]='h000023d4;  wr_data_rom[ 6520]='h0000242e;
    rd_cycle[ 6521] = 1'b0;  wr_cycle[ 6521] = 1'b1;  addr_rom[ 6521]='h00001e7c;  wr_data_rom[ 6521]='h00000a87;
    rd_cycle[ 6522] = 1'b1;  wr_cycle[ 6522] = 1'b0;  addr_rom[ 6522]='h00001fa8;  wr_data_rom[ 6522]='h00000000;
    rd_cycle[ 6523] = 1'b0;  wr_cycle[ 6523] = 1'b1;  addr_rom[ 6523]='h0000017c;  wr_data_rom[ 6523]='h00001a0e;
    rd_cycle[ 6524] = 1'b0;  wr_cycle[ 6524] = 1'b1;  addr_rom[ 6524]='h000025d8;  wr_data_rom[ 6524]='h00002817;
    rd_cycle[ 6525] = 1'b1;  wr_cycle[ 6525] = 1'b0;  addr_rom[ 6525]='h00000c10;  wr_data_rom[ 6525]='h00000000;
    rd_cycle[ 6526] = 1'b1;  wr_cycle[ 6526] = 1'b0;  addr_rom[ 6526]='h000008c4;  wr_data_rom[ 6526]='h00000000;
    rd_cycle[ 6527] = 1'b1;  wr_cycle[ 6527] = 1'b0;  addr_rom[ 6527]='h000009a4;  wr_data_rom[ 6527]='h00000000;
    rd_cycle[ 6528] = 1'b1;  wr_cycle[ 6528] = 1'b0;  addr_rom[ 6528]='h00003bd8;  wr_data_rom[ 6528]='h00000000;
    rd_cycle[ 6529] = 1'b0;  wr_cycle[ 6529] = 1'b1;  addr_rom[ 6529]='h00000500;  wr_data_rom[ 6529]='h00002996;
    rd_cycle[ 6530] = 1'b0;  wr_cycle[ 6530] = 1'b1;  addr_rom[ 6530]='h000008d0;  wr_data_rom[ 6530]='h00001b51;
    rd_cycle[ 6531] = 1'b1;  wr_cycle[ 6531] = 1'b0;  addr_rom[ 6531]='h00001fc8;  wr_data_rom[ 6531]='h00000000;
    rd_cycle[ 6532] = 1'b1;  wr_cycle[ 6532] = 1'b0;  addr_rom[ 6532]='h00003590;  wr_data_rom[ 6532]='h00000000;
    rd_cycle[ 6533] = 1'b0;  wr_cycle[ 6533] = 1'b1;  addr_rom[ 6533]='h00003b54;  wr_data_rom[ 6533]='h00000bd5;
    rd_cycle[ 6534] = 1'b1;  wr_cycle[ 6534] = 1'b0;  addr_rom[ 6534]='h00002d78;  wr_data_rom[ 6534]='h00000000;
    rd_cycle[ 6535] = 1'b0;  wr_cycle[ 6535] = 1'b1;  addr_rom[ 6535]='h00002f84;  wr_data_rom[ 6535]='h00001191;
    rd_cycle[ 6536] = 1'b1;  wr_cycle[ 6536] = 1'b0;  addr_rom[ 6536]='h0000249c;  wr_data_rom[ 6536]='h00000000;
    rd_cycle[ 6537] = 1'b1;  wr_cycle[ 6537] = 1'b0;  addr_rom[ 6537]='h00002e44;  wr_data_rom[ 6537]='h00000000;
    rd_cycle[ 6538] = 1'b1;  wr_cycle[ 6538] = 1'b0;  addr_rom[ 6538]='h00001258;  wr_data_rom[ 6538]='h00000000;
    rd_cycle[ 6539] = 1'b1;  wr_cycle[ 6539] = 1'b0;  addr_rom[ 6539]='h0000344c;  wr_data_rom[ 6539]='h00000000;
    rd_cycle[ 6540] = 1'b0;  wr_cycle[ 6540] = 1'b1;  addr_rom[ 6540]='h00001fdc;  wr_data_rom[ 6540]='h0000002b;
    rd_cycle[ 6541] = 1'b0;  wr_cycle[ 6541] = 1'b1;  addr_rom[ 6541]='h00003d88;  wr_data_rom[ 6541]='h000004dc;
    rd_cycle[ 6542] = 1'b1;  wr_cycle[ 6542] = 1'b0;  addr_rom[ 6542]='h0000285c;  wr_data_rom[ 6542]='h00000000;
    rd_cycle[ 6543] = 1'b0;  wr_cycle[ 6543] = 1'b1;  addr_rom[ 6543]='h00001e84;  wr_data_rom[ 6543]='h0000267d;
    rd_cycle[ 6544] = 1'b1;  wr_cycle[ 6544] = 1'b0;  addr_rom[ 6544]='h00003fa8;  wr_data_rom[ 6544]='h00000000;
    rd_cycle[ 6545] = 1'b1;  wr_cycle[ 6545] = 1'b0;  addr_rom[ 6545]='h000000a0;  wr_data_rom[ 6545]='h00000000;
    rd_cycle[ 6546] = 1'b1;  wr_cycle[ 6546] = 1'b0;  addr_rom[ 6546]='h000029f4;  wr_data_rom[ 6546]='h00000000;
    rd_cycle[ 6547] = 1'b1;  wr_cycle[ 6547] = 1'b0;  addr_rom[ 6547]='h00002bb0;  wr_data_rom[ 6547]='h00000000;
    rd_cycle[ 6548] = 1'b1;  wr_cycle[ 6548] = 1'b0;  addr_rom[ 6548]='h000016f8;  wr_data_rom[ 6548]='h00000000;
    rd_cycle[ 6549] = 1'b0;  wr_cycle[ 6549] = 1'b1;  addr_rom[ 6549]='h00000338;  wr_data_rom[ 6549]='h00003be4;
    rd_cycle[ 6550] = 1'b0;  wr_cycle[ 6550] = 1'b1;  addr_rom[ 6550]='h00001cd4;  wr_data_rom[ 6550]='h00001b19;
    rd_cycle[ 6551] = 1'b0;  wr_cycle[ 6551] = 1'b1;  addr_rom[ 6551]='h000018d0;  wr_data_rom[ 6551]='h000006f2;
    rd_cycle[ 6552] = 1'b1;  wr_cycle[ 6552] = 1'b0;  addr_rom[ 6552]='h00002678;  wr_data_rom[ 6552]='h00000000;
    rd_cycle[ 6553] = 1'b1;  wr_cycle[ 6553] = 1'b0;  addr_rom[ 6553]='h000018d8;  wr_data_rom[ 6553]='h00000000;
    rd_cycle[ 6554] = 1'b1;  wr_cycle[ 6554] = 1'b0;  addr_rom[ 6554]='h00002c0c;  wr_data_rom[ 6554]='h00000000;
    rd_cycle[ 6555] = 1'b0;  wr_cycle[ 6555] = 1'b1;  addr_rom[ 6555]='h00000c00;  wr_data_rom[ 6555]='h0000273c;
    rd_cycle[ 6556] = 1'b0;  wr_cycle[ 6556] = 1'b1;  addr_rom[ 6556]='h00000074;  wr_data_rom[ 6556]='h00001f8d;
    rd_cycle[ 6557] = 1'b0;  wr_cycle[ 6557] = 1'b1;  addr_rom[ 6557]='h00001088;  wr_data_rom[ 6557]='h00000c9f;
    rd_cycle[ 6558] = 1'b0;  wr_cycle[ 6558] = 1'b1;  addr_rom[ 6558]='h00003d08;  wr_data_rom[ 6558]='h00002887;
    rd_cycle[ 6559] = 1'b0;  wr_cycle[ 6559] = 1'b1;  addr_rom[ 6559]='h0000359c;  wr_data_rom[ 6559]='h00001211;
    rd_cycle[ 6560] = 1'b0;  wr_cycle[ 6560] = 1'b1;  addr_rom[ 6560]='h000022d8;  wr_data_rom[ 6560]='h00000032;
    rd_cycle[ 6561] = 1'b1;  wr_cycle[ 6561] = 1'b0;  addr_rom[ 6561]='h00002458;  wr_data_rom[ 6561]='h00000000;
    rd_cycle[ 6562] = 1'b1;  wr_cycle[ 6562] = 1'b0;  addr_rom[ 6562]='h000027f0;  wr_data_rom[ 6562]='h00000000;
    rd_cycle[ 6563] = 1'b1;  wr_cycle[ 6563] = 1'b0;  addr_rom[ 6563]='h00000104;  wr_data_rom[ 6563]='h00000000;
    rd_cycle[ 6564] = 1'b1;  wr_cycle[ 6564] = 1'b0;  addr_rom[ 6564]='h00000978;  wr_data_rom[ 6564]='h00000000;
    rd_cycle[ 6565] = 1'b1;  wr_cycle[ 6565] = 1'b0;  addr_rom[ 6565]='h000015f0;  wr_data_rom[ 6565]='h00000000;
    rd_cycle[ 6566] = 1'b1;  wr_cycle[ 6566] = 1'b0;  addr_rom[ 6566]='h0000030c;  wr_data_rom[ 6566]='h00000000;
    rd_cycle[ 6567] = 1'b1;  wr_cycle[ 6567] = 1'b0;  addr_rom[ 6567]='h00003344;  wr_data_rom[ 6567]='h00000000;
    rd_cycle[ 6568] = 1'b1;  wr_cycle[ 6568] = 1'b0;  addr_rom[ 6568]='h00001ed4;  wr_data_rom[ 6568]='h00000000;
    rd_cycle[ 6569] = 1'b1;  wr_cycle[ 6569] = 1'b0;  addr_rom[ 6569]='h00001620;  wr_data_rom[ 6569]='h00000000;
    rd_cycle[ 6570] = 1'b1;  wr_cycle[ 6570] = 1'b0;  addr_rom[ 6570]='h000016f8;  wr_data_rom[ 6570]='h00000000;
    rd_cycle[ 6571] = 1'b0;  wr_cycle[ 6571] = 1'b1;  addr_rom[ 6571]='h00003c00;  wr_data_rom[ 6571]='h00000c75;
    rd_cycle[ 6572] = 1'b0;  wr_cycle[ 6572] = 1'b1;  addr_rom[ 6572]='h00000534;  wr_data_rom[ 6572]='h000006ae;
    rd_cycle[ 6573] = 1'b1;  wr_cycle[ 6573] = 1'b0;  addr_rom[ 6573]='h00002700;  wr_data_rom[ 6573]='h00000000;
    rd_cycle[ 6574] = 1'b1;  wr_cycle[ 6574] = 1'b0;  addr_rom[ 6574]='h00001594;  wr_data_rom[ 6574]='h00000000;
    rd_cycle[ 6575] = 1'b1;  wr_cycle[ 6575] = 1'b0;  addr_rom[ 6575]='h00002b98;  wr_data_rom[ 6575]='h00000000;
    rd_cycle[ 6576] = 1'b1;  wr_cycle[ 6576] = 1'b0;  addr_rom[ 6576]='h00000fa8;  wr_data_rom[ 6576]='h00000000;
    rd_cycle[ 6577] = 1'b1;  wr_cycle[ 6577] = 1'b0;  addr_rom[ 6577]='h00001bb0;  wr_data_rom[ 6577]='h00000000;
    rd_cycle[ 6578] = 1'b0;  wr_cycle[ 6578] = 1'b1;  addr_rom[ 6578]='h000030d0;  wr_data_rom[ 6578]='h000017ad;
    rd_cycle[ 6579] = 1'b1;  wr_cycle[ 6579] = 1'b0;  addr_rom[ 6579]='h00002a4c;  wr_data_rom[ 6579]='h00000000;
    rd_cycle[ 6580] = 1'b0;  wr_cycle[ 6580] = 1'b1;  addr_rom[ 6580]='h00002784;  wr_data_rom[ 6580]='h00000133;
    rd_cycle[ 6581] = 1'b0;  wr_cycle[ 6581] = 1'b1;  addr_rom[ 6581]='h000014c4;  wr_data_rom[ 6581]='h00001a18;
    rd_cycle[ 6582] = 1'b1;  wr_cycle[ 6582] = 1'b0;  addr_rom[ 6582]='h00002c1c;  wr_data_rom[ 6582]='h00000000;
    rd_cycle[ 6583] = 1'b1;  wr_cycle[ 6583] = 1'b0;  addr_rom[ 6583]='h00003c00;  wr_data_rom[ 6583]='h00000000;
    rd_cycle[ 6584] = 1'b1;  wr_cycle[ 6584] = 1'b0;  addr_rom[ 6584]='h00000640;  wr_data_rom[ 6584]='h00000000;
    rd_cycle[ 6585] = 1'b1;  wr_cycle[ 6585] = 1'b0;  addr_rom[ 6585]='h000039a8;  wr_data_rom[ 6585]='h00000000;
    rd_cycle[ 6586] = 1'b1;  wr_cycle[ 6586] = 1'b0;  addr_rom[ 6586]='h00001624;  wr_data_rom[ 6586]='h00000000;
    rd_cycle[ 6587] = 1'b0;  wr_cycle[ 6587] = 1'b1;  addr_rom[ 6587]='h000029e4;  wr_data_rom[ 6587]='h00000f5e;
    rd_cycle[ 6588] = 1'b1;  wr_cycle[ 6588] = 1'b0;  addr_rom[ 6588]='h00003d68;  wr_data_rom[ 6588]='h00000000;
    rd_cycle[ 6589] = 1'b1;  wr_cycle[ 6589] = 1'b0;  addr_rom[ 6589]='h000034f0;  wr_data_rom[ 6589]='h00000000;
    rd_cycle[ 6590] = 1'b1;  wr_cycle[ 6590] = 1'b0;  addr_rom[ 6590]='h000030c4;  wr_data_rom[ 6590]='h00000000;
    rd_cycle[ 6591] = 1'b1;  wr_cycle[ 6591] = 1'b0;  addr_rom[ 6591]='h00002174;  wr_data_rom[ 6591]='h00000000;
    rd_cycle[ 6592] = 1'b1;  wr_cycle[ 6592] = 1'b0;  addr_rom[ 6592]='h00000d68;  wr_data_rom[ 6592]='h00000000;
    rd_cycle[ 6593] = 1'b0;  wr_cycle[ 6593] = 1'b1;  addr_rom[ 6593]='h0000109c;  wr_data_rom[ 6593]='h0000164c;
    rd_cycle[ 6594] = 1'b1;  wr_cycle[ 6594] = 1'b0;  addr_rom[ 6594]='h00002898;  wr_data_rom[ 6594]='h00000000;
    rd_cycle[ 6595] = 1'b0;  wr_cycle[ 6595] = 1'b1;  addr_rom[ 6595]='h000034c0;  wr_data_rom[ 6595]='h000014b6;
    rd_cycle[ 6596] = 1'b1;  wr_cycle[ 6596] = 1'b0;  addr_rom[ 6596]='h000010c4;  wr_data_rom[ 6596]='h00000000;
    rd_cycle[ 6597] = 1'b1;  wr_cycle[ 6597] = 1'b0;  addr_rom[ 6597]='h0000255c;  wr_data_rom[ 6597]='h00000000;
    rd_cycle[ 6598] = 1'b0;  wr_cycle[ 6598] = 1'b1;  addr_rom[ 6598]='h00001024;  wr_data_rom[ 6598]='h000028d4;
    rd_cycle[ 6599] = 1'b0;  wr_cycle[ 6599] = 1'b1;  addr_rom[ 6599]='h00003ab0;  wr_data_rom[ 6599]='h00001653;
    rd_cycle[ 6600] = 1'b0;  wr_cycle[ 6600] = 1'b1;  addr_rom[ 6600]='h00001540;  wr_data_rom[ 6600]='h00002a40;
    rd_cycle[ 6601] = 1'b0;  wr_cycle[ 6601] = 1'b1;  addr_rom[ 6601]='h00000fc0;  wr_data_rom[ 6601]='h00000913;
    rd_cycle[ 6602] = 1'b1;  wr_cycle[ 6602] = 1'b0;  addr_rom[ 6602]='h00003e08;  wr_data_rom[ 6602]='h00000000;
    rd_cycle[ 6603] = 1'b0;  wr_cycle[ 6603] = 1'b1;  addr_rom[ 6603]='h00001210;  wr_data_rom[ 6603]='h00001a98;
    rd_cycle[ 6604] = 1'b0;  wr_cycle[ 6604] = 1'b1;  addr_rom[ 6604]='h00000f0c;  wr_data_rom[ 6604]='h00003004;
    rd_cycle[ 6605] = 1'b0;  wr_cycle[ 6605] = 1'b1;  addr_rom[ 6605]='h00001400;  wr_data_rom[ 6605]='h00002228;
    rd_cycle[ 6606] = 1'b0;  wr_cycle[ 6606] = 1'b1;  addr_rom[ 6606]='h00000a30;  wr_data_rom[ 6606]='h000016bb;
    rd_cycle[ 6607] = 1'b1;  wr_cycle[ 6607] = 1'b0;  addr_rom[ 6607]='h000025b8;  wr_data_rom[ 6607]='h00000000;
    rd_cycle[ 6608] = 1'b0;  wr_cycle[ 6608] = 1'b1;  addr_rom[ 6608]='h00002d0c;  wr_data_rom[ 6608]='h00002521;
    rd_cycle[ 6609] = 1'b0;  wr_cycle[ 6609] = 1'b1;  addr_rom[ 6609]='h00001350;  wr_data_rom[ 6609]='h00002113;
    rd_cycle[ 6610] = 1'b0;  wr_cycle[ 6610] = 1'b1;  addr_rom[ 6610]='h000024f4;  wr_data_rom[ 6610]='h000014dd;
    rd_cycle[ 6611] = 1'b0;  wr_cycle[ 6611] = 1'b1;  addr_rom[ 6611]='h00000598;  wr_data_rom[ 6611]='h000037b4;
    rd_cycle[ 6612] = 1'b0;  wr_cycle[ 6612] = 1'b1;  addr_rom[ 6612]='h000011f8;  wr_data_rom[ 6612]='h00001599;
    rd_cycle[ 6613] = 1'b0;  wr_cycle[ 6613] = 1'b1;  addr_rom[ 6613]='h000001e4;  wr_data_rom[ 6613]='h0000121b;
    rd_cycle[ 6614] = 1'b0;  wr_cycle[ 6614] = 1'b1;  addr_rom[ 6614]='h000012b4;  wr_data_rom[ 6614]='h00000965;
    rd_cycle[ 6615] = 1'b1;  wr_cycle[ 6615] = 1'b0;  addr_rom[ 6615]='h0000214c;  wr_data_rom[ 6615]='h00000000;
    rd_cycle[ 6616] = 1'b0;  wr_cycle[ 6616] = 1'b1;  addr_rom[ 6616]='h0000325c;  wr_data_rom[ 6616]='h000017b2;
    rd_cycle[ 6617] = 1'b0;  wr_cycle[ 6617] = 1'b1;  addr_rom[ 6617]='h0000157c;  wr_data_rom[ 6617]='h00002679;
    rd_cycle[ 6618] = 1'b0;  wr_cycle[ 6618] = 1'b1;  addr_rom[ 6618]='h0000043c;  wr_data_rom[ 6618]='h00001e5c;
    rd_cycle[ 6619] = 1'b0;  wr_cycle[ 6619] = 1'b1;  addr_rom[ 6619]='h000014b8;  wr_data_rom[ 6619]='h0000268e;
    rd_cycle[ 6620] = 1'b1;  wr_cycle[ 6620] = 1'b0;  addr_rom[ 6620]='h0000360c;  wr_data_rom[ 6620]='h00000000;
    rd_cycle[ 6621] = 1'b1;  wr_cycle[ 6621] = 1'b0;  addr_rom[ 6621]='h0000064c;  wr_data_rom[ 6621]='h00000000;
    rd_cycle[ 6622] = 1'b0;  wr_cycle[ 6622] = 1'b1;  addr_rom[ 6622]='h0000296c;  wr_data_rom[ 6622]='h00001412;
    rd_cycle[ 6623] = 1'b0;  wr_cycle[ 6623] = 1'b1;  addr_rom[ 6623]='h000038b8;  wr_data_rom[ 6623]='h000035dd;
    rd_cycle[ 6624] = 1'b1;  wr_cycle[ 6624] = 1'b0;  addr_rom[ 6624]='h00000398;  wr_data_rom[ 6624]='h00000000;
    rd_cycle[ 6625] = 1'b1;  wr_cycle[ 6625] = 1'b0;  addr_rom[ 6625]='h00000b60;  wr_data_rom[ 6625]='h00000000;
    rd_cycle[ 6626] = 1'b1;  wr_cycle[ 6626] = 1'b0;  addr_rom[ 6626]='h00003668;  wr_data_rom[ 6626]='h00000000;
    rd_cycle[ 6627] = 1'b1;  wr_cycle[ 6627] = 1'b0;  addr_rom[ 6627]='h00003ee4;  wr_data_rom[ 6627]='h00000000;
    rd_cycle[ 6628] = 1'b0;  wr_cycle[ 6628] = 1'b1;  addr_rom[ 6628]='h00000450;  wr_data_rom[ 6628]='h00002740;
    rd_cycle[ 6629] = 1'b0;  wr_cycle[ 6629] = 1'b1;  addr_rom[ 6629]='h00000fe0;  wr_data_rom[ 6629]='h00000eb8;
    rd_cycle[ 6630] = 1'b0;  wr_cycle[ 6630] = 1'b1;  addr_rom[ 6630]='h00003510;  wr_data_rom[ 6630]='h0000346a;
    rd_cycle[ 6631] = 1'b1;  wr_cycle[ 6631] = 1'b0;  addr_rom[ 6631]='h000023e0;  wr_data_rom[ 6631]='h00000000;
    rd_cycle[ 6632] = 1'b0;  wr_cycle[ 6632] = 1'b1;  addr_rom[ 6632]='h000031cc;  wr_data_rom[ 6632]='h000030fb;
    rd_cycle[ 6633] = 1'b1;  wr_cycle[ 6633] = 1'b0;  addr_rom[ 6633]='h000018b4;  wr_data_rom[ 6633]='h00000000;
    rd_cycle[ 6634] = 1'b1;  wr_cycle[ 6634] = 1'b0;  addr_rom[ 6634]='h00000ce0;  wr_data_rom[ 6634]='h00000000;
    rd_cycle[ 6635] = 1'b0;  wr_cycle[ 6635] = 1'b1;  addr_rom[ 6635]='h00000f04;  wr_data_rom[ 6635]='h00000b95;
    rd_cycle[ 6636] = 1'b0;  wr_cycle[ 6636] = 1'b1;  addr_rom[ 6636]='h00001d38;  wr_data_rom[ 6636]='h00000fcb;
    rd_cycle[ 6637] = 1'b0;  wr_cycle[ 6637] = 1'b1;  addr_rom[ 6637]='h00002058;  wr_data_rom[ 6637]='h00002b9d;
    rd_cycle[ 6638] = 1'b1;  wr_cycle[ 6638] = 1'b0;  addr_rom[ 6638]='h00002d9c;  wr_data_rom[ 6638]='h00000000;
    rd_cycle[ 6639] = 1'b0;  wr_cycle[ 6639] = 1'b1;  addr_rom[ 6639]='h000021a4;  wr_data_rom[ 6639]='h00001685;
    rd_cycle[ 6640] = 1'b1;  wr_cycle[ 6640] = 1'b0;  addr_rom[ 6640]='h00000574;  wr_data_rom[ 6640]='h00000000;
    rd_cycle[ 6641] = 1'b0;  wr_cycle[ 6641] = 1'b1;  addr_rom[ 6641]='h00003c80;  wr_data_rom[ 6641]='h0000179c;
    rd_cycle[ 6642] = 1'b0;  wr_cycle[ 6642] = 1'b1;  addr_rom[ 6642]='h00002e64;  wr_data_rom[ 6642]='h00001187;
    rd_cycle[ 6643] = 1'b1;  wr_cycle[ 6643] = 1'b0;  addr_rom[ 6643]='h00002d64;  wr_data_rom[ 6643]='h00000000;
    rd_cycle[ 6644] = 1'b1;  wr_cycle[ 6644] = 1'b0;  addr_rom[ 6644]='h0000151c;  wr_data_rom[ 6644]='h00000000;
    rd_cycle[ 6645] = 1'b1;  wr_cycle[ 6645] = 1'b0;  addr_rom[ 6645]='h00002fd4;  wr_data_rom[ 6645]='h00000000;
    rd_cycle[ 6646] = 1'b1;  wr_cycle[ 6646] = 1'b0;  addr_rom[ 6646]='h00002d0c;  wr_data_rom[ 6646]='h00000000;
    rd_cycle[ 6647] = 1'b0;  wr_cycle[ 6647] = 1'b1;  addr_rom[ 6647]='h00000048;  wr_data_rom[ 6647]='h00001eb8;
    rd_cycle[ 6648] = 1'b1;  wr_cycle[ 6648] = 1'b0;  addr_rom[ 6648]='h00002c14;  wr_data_rom[ 6648]='h00000000;
    rd_cycle[ 6649] = 1'b1;  wr_cycle[ 6649] = 1'b0;  addr_rom[ 6649]='h00000238;  wr_data_rom[ 6649]='h00000000;
    rd_cycle[ 6650] = 1'b1;  wr_cycle[ 6650] = 1'b0;  addr_rom[ 6650]='h00000d20;  wr_data_rom[ 6650]='h00000000;
    rd_cycle[ 6651] = 1'b0;  wr_cycle[ 6651] = 1'b1;  addr_rom[ 6651]='h00002a20;  wr_data_rom[ 6651]='h00000b36;
    rd_cycle[ 6652] = 1'b0;  wr_cycle[ 6652] = 1'b1;  addr_rom[ 6652]='h00003670;  wr_data_rom[ 6652]='h00002b1d;
    rd_cycle[ 6653] = 1'b1;  wr_cycle[ 6653] = 1'b0;  addr_rom[ 6653]='h00002b4c;  wr_data_rom[ 6653]='h00000000;
    rd_cycle[ 6654] = 1'b1;  wr_cycle[ 6654] = 1'b0;  addr_rom[ 6654]='h000011e4;  wr_data_rom[ 6654]='h00000000;
    rd_cycle[ 6655] = 1'b0;  wr_cycle[ 6655] = 1'b1;  addr_rom[ 6655]='h000027fc;  wr_data_rom[ 6655]='h000031b4;
    rd_cycle[ 6656] = 1'b1;  wr_cycle[ 6656] = 1'b0;  addr_rom[ 6656]='h00000fb0;  wr_data_rom[ 6656]='h00000000;
    rd_cycle[ 6657] = 1'b0;  wr_cycle[ 6657] = 1'b1;  addr_rom[ 6657]='h00003e64;  wr_data_rom[ 6657]='h00002e84;
    rd_cycle[ 6658] = 1'b1;  wr_cycle[ 6658] = 1'b0;  addr_rom[ 6658]='h00002250;  wr_data_rom[ 6658]='h00000000;
    rd_cycle[ 6659] = 1'b0;  wr_cycle[ 6659] = 1'b1;  addr_rom[ 6659]='h00002f40;  wr_data_rom[ 6659]='h000030f1;
    rd_cycle[ 6660] = 1'b0;  wr_cycle[ 6660] = 1'b1;  addr_rom[ 6660]='h0000344c;  wr_data_rom[ 6660]='h00003f55;
    rd_cycle[ 6661] = 1'b0;  wr_cycle[ 6661] = 1'b1;  addr_rom[ 6661]='h0000013c;  wr_data_rom[ 6661]='h0000397c;
    rd_cycle[ 6662] = 1'b0;  wr_cycle[ 6662] = 1'b1;  addr_rom[ 6662]='h00003004;  wr_data_rom[ 6662]='h00001900;
    rd_cycle[ 6663] = 1'b1;  wr_cycle[ 6663] = 1'b0;  addr_rom[ 6663]='h00002c1c;  wr_data_rom[ 6663]='h00000000;
    rd_cycle[ 6664] = 1'b1;  wr_cycle[ 6664] = 1'b0;  addr_rom[ 6664]='h00000844;  wr_data_rom[ 6664]='h00000000;
    rd_cycle[ 6665] = 1'b0;  wr_cycle[ 6665] = 1'b1;  addr_rom[ 6665]='h00001eac;  wr_data_rom[ 6665]='h000019da;
    rd_cycle[ 6666] = 1'b1;  wr_cycle[ 6666] = 1'b0;  addr_rom[ 6666]='h00003f78;  wr_data_rom[ 6666]='h00000000;
    rd_cycle[ 6667] = 1'b0;  wr_cycle[ 6667] = 1'b1;  addr_rom[ 6667]='h00002074;  wr_data_rom[ 6667]='h000015e5;
    rd_cycle[ 6668] = 1'b1;  wr_cycle[ 6668] = 1'b0;  addr_rom[ 6668]='h000022cc;  wr_data_rom[ 6668]='h00000000;
    rd_cycle[ 6669] = 1'b1;  wr_cycle[ 6669] = 1'b0;  addr_rom[ 6669]='h00000478;  wr_data_rom[ 6669]='h00000000;
    rd_cycle[ 6670] = 1'b1;  wr_cycle[ 6670] = 1'b0;  addr_rom[ 6670]='h000018ac;  wr_data_rom[ 6670]='h00000000;
    rd_cycle[ 6671] = 1'b0;  wr_cycle[ 6671] = 1'b1;  addr_rom[ 6671]='h00003fa8;  wr_data_rom[ 6671]='h000034d5;
    rd_cycle[ 6672] = 1'b1;  wr_cycle[ 6672] = 1'b0;  addr_rom[ 6672]='h0000379c;  wr_data_rom[ 6672]='h00000000;
    rd_cycle[ 6673] = 1'b0;  wr_cycle[ 6673] = 1'b1;  addr_rom[ 6673]='h000035e0;  wr_data_rom[ 6673]='h00002611;
    rd_cycle[ 6674] = 1'b1;  wr_cycle[ 6674] = 1'b0;  addr_rom[ 6674]='h000009b8;  wr_data_rom[ 6674]='h00000000;
    rd_cycle[ 6675] = 1'b1;  wr_cycle[ 6675] = 1'b0;  addr_rom[ 6675]='h00002878;  wr_data_rom[ 6675]='h00000000;
    rd_cycle[ 6676] = 1'b0;  wr_cycle[ 6676] = 1'b1;  addr_rom[ 6676]='h0000168c;  wr_data_rom[ 6676]='h000030ed;
    rd_cycle[ 6677] = 1'b1;  wr_cycle[ 6677] = 1'b0;  addr_rom[ 6677]='h00003264;  wr_data_rom[ 6677]='h00000000;
    rd_cycle[ 6678] = 1'b1;  wr_cycle[ 6678] = 1'b0;  addr_rom[ 6678]='h000012a4;  wr_data_rom[ 6678]='h00000000;
    rd_cycle[ 6679] = 1'b0;  wr_cycle[ 6679] = 1'b1;  addr_rom[ 6679]='h000033f4;  wr_data_rom[ 6679]='h00003880;
    rd_cycle[ 6680] = 1'b0;  wr_cycle[ 6680] = 1'b1;  addr_rom[ 6680]='h00003304;  wr_data_rom[ 6680]='h00000865;
    rd_cycle[ 6681] = 1'b1;  wr_cycle[ 6681] = 1'b0;  addr_rom[ 6681]='h00001380;  wr_data_rom[ 6681]='h00000000;
    rd_cycle[ 6682] = 1'b0;  wr_cycle[ 6682] = 1'b1;  addr_rom[ 6682]='h00000798;  wr_data_rom[ 6682]='h000005e8;
    rd_cycle[ 6683] = 1'b1;  wr_cycle[ 6683] = 1'b0;  addr_rom[ 6683]='h00002190;  wr_data_rom[ 6683]='h00000000;
    rd_cycle[ 6684] = 1'b1;  wr_cycle[ 6684] = 1'b0;  addr_rom[ 6684]='h000029e8;  wr_data_rom[ 6684]='h00000000;
    rd_cycle[ 6685] = 1'b0;  wr_cycle[ 6685] = 1'b1;  addr_rom[ 6685]='h00001694;  wr_data_rom[ 6685]='h00001df8;
    rd_cycle[ 6686] = 1'b1;  wr_cycle[ 6686] = 1'b0;  addr_rom[ 6686]='h000038b8;  wr_data_rom[ 6686]='h00000000;
    rd_cycle[ 6687] = 1'b0;  wr_cycle[ 6687] = 1'b1;  addr_rom[ 6687]='h00000810;  wr_data_rom[ 6687]='h00003b0f;
    rd_cycle[ 6688] = 1'b1;  wr_cycle[ 6688] = 1'b0;  addr_rom[ 6688]='h00000cdc;  wr_data_rom[ 6688]='h00000000;
    rd_cycle[ 6689] = 1'b1;  wr_cycle[ 6689] = 1'b0;  addr_rom[ 6689]='h00002d04;  wr_data_rom[ 6689]='h00000000;
    rd_cycle[ 6690] = 1'b0;  wr_cycle[ 6690] = 1'b1;  addr_rom[ 6690]='h0000047c;  wr_data_rom[ 6690]='h00002726;
    rd_cycle[ 6691] = 1'b0;  wr_cycle[ 6691] = 1'b1;  addr_rom[ 6691]='h00000d3c;  wr_data_rom[ 6691]='h00003cf8;
    rd_cycle[ 6692] = 1'b0;  wr_cycle[ 6692] = 1'b1;  addr_rom[ 6692]='h000008ec;  wr_data_rom[ 6692]='h000026e6;
    rd_cycle[ 6693] = 1'b0;  wr_cycle[ 6693] = 1'b1;  addr_rom[ 6693]='h00003c64;  wr_data_rom[ 6693]='h000033ca;
    rd_cycle[ 6694] = 1'b1;  wr_cycle[ 6694] = 1'b0;  addr_rom[ 6694]='h000039a4;  wr_data_rom[ 6694]='h00000000;
    rd_cycle[ 6695] = 1'b1;  wr_cycle[ 6695] = 1'b0;  addr_rom[ 6695]='h00002260;  wr_data_rom[ 6695]='h00000000;
    rd_cycle[ 6696] = 1'b1;  wr_cycle[ 6696] = 1'b0;  addr_rom[ 6696]='h0000307c;  wr_data_rom[ 6696]='h00000000;
    rd_cycle[ 6697] = 1'b0;  wr_cycle[ 6697] = 1'b1;  addr_rom[ 6697]='h000015f8;  wr_data_rom[ 6697]='h0000004a;
    rd_cycle[ 6698] = 1'b0;  wr_cycle[ 6698] = 1'b1;  addr_rom[ 6698]='h00000848;  wr_data_rom[ 6698]='h000022c8;
    rd_cycle[ 6699] = 1'b0;  wr_cycle[ 6699] = 1'b1;  addr_rom[ 6699]='h00002674;  wr_data_rom[ 6699]='h00001c70;
    rd_cycle[ 6700] = 1'b1;  wr_cycle[ 6700] = 1'b0;  addr_rom[ 6700]='h00001f8c;  wr_data_rom[ 6700]='h00000000;
    rd_cycle[ 6701] = 1'b0;  wr_cycle[ 6701] = 1'b1;  addr_rom[ 6701]='h00000c70;  wr_data_rom[ 6701]='h0000253b;
    rd_cycle[ 6702] = 1'b1;  wr_cycle[ 6702] = 1'b0;  addr_rom[ 6702]='h00000710;  wr_data_rom[ 6702]='h00000000;
    rd_cycle[ 6703] = 1'b0;  wr_cycle[ 6703] = 1'b1;  addr_rom[ 6703]='h000008fc;  wr_data_rom[ 6703]='h00002bdc;
    rd_cycle[ 6704] = 1'b0;  wr_cycle[ 6704] = 1'b1;  addr_rom[ 6704]='h000004d0;  wr_data_rom[ 6704]='h000025a7;
    rd_cycle[ 6705] = 1'b0;  wr_cycle[ 6705] = 1'b1;  addr_rom[ 6705]='h00000a74;  wr_data_rom[ 6705]='h000035e1;
    rd_cycle[ 6706] = 1'b0;  wr_cycle[ 6706] = 1'b1;  addr_rom[ 6706]='h00002450;  wr_data_rom[ 6706]='h000038cb;
    rd_cycle[ 6707] = 1'b1;  wr_cycle[ 6707] = 1'b0;  addr_rom[ 6707]='h000012b8;  wr_data_rom[ 6707]='h00000000;
    rd_cycle[ 6708] = 1'b0;  wr_cycle[ 6708] = 1'b1;  addr_rom[ 6708]='h000002e4;  wr_data_rom[ 6708]='h00000979;
    rd_cycle[ 6709] = 1'b0;  wr_cycle[ 6709] = 1'b1;  addr_rom[ 6709]='h000007fc;  wr_data_rom[ 6709]='h0000064b;
    rd_cycle[ 6710] = 1'b0;  wr_cycle[ 6710] = 1'b1;  addr_rom[ 6710]='h00001274;  wr_data_rom[ 6710]='h0000274e;
    rd_cycle[ 6711] = 1'b1;  wr_cycle[ 6711] = 1'b0;  addr_rom[ 6711]='h00003ae8;  wr_data_rom[ 6711]='h00000000;
    rd_cycle[ 6712] = 1'b1;  wr_cycle[ 6712] = 1'b0;  addr_rom[ 6712]='h0000038c;  wr_data_rom[ 6712]='h00000000;
    rd_cycle[ 6713] = 1'b1;  wr_cycle[ 6713] = 1'b0;  addr_rom[ 6713]='h0000263c;  wr_data_rom[ 6713]='h00000000;
    rd_cycle[ 6714] = 1'b0;  wr_cycle[ 6714] = 1'b1;  addr_rom[ 6714]='h00000734;  wr_data_rom[ 6714]='h000024d1;
    rd_cycle[ 6715] = 1'b1;  wr_cycle[ 6715] = 1'b0;  addr_rom[ 6715]='h0000060c;  wr_data_rom[ 6715]='h00000000;
    rd_cycle[ 6716] = 1'b0;  wr_cycle[ 6716] = 1'b1;  addr_rom[ 6716]='h00003c28;  wr_data_rom[ 6716]='h000022bf;
    rd_cycle[ 6717] = 1'b0;  wr_cycle[ 6717] = 1'b1;  addr_rom[ 6717]='h00003d40;  wr_data_rom[ 6717]='h000027ad;
    rd_cycle[ 6718] = 1'b0;  wr_cycle[ 6718] = 1'b1;  addr_rom[ 6718]='h00002c58;  wr_data_rom[ 6718]='h000035bf;
    rd_cycle[ 6719] = 1'b0;  wr_cycle[ 6719] = 1'b1;  addr_rom[ 6719]='h00002cb8;  wr_data_rom[ 6719]='h000014b4;
    rd_cycle[ 6720] = 1'b0;  wr_cycle[ 6720] = 1'b1;  addr_rom[ 6720]='h00000ab8;  wr_data_rom[ 6720]='h00003494;
    rd_cycle[ 6721] = 1'b0;  wr_cycle[ 6721] = 1'b1;  addr_rom[ 6721]='h00001984;  wr_data_rom[ 6721]='h000006df;
    rd_cycle[ 6722] = 1'b1;  wr_cycle[ 6722] = 1'b0;  addr_rom[ 6722]='h00000a20;  wr_data_rom[ 6722]='h00000000;
    rd_cycle[ 6723] = 1'b1;  wr_cycle[ 6723] = 1'b0;  addr_rom[ 6723]='h00003230;  wr_data_rom[ 6723]='h00000000;
    rd_cycle[ 6724] = 1'b1;  wr_cycle[ 6724] = 1'b0;  addr_rom[ 6724]='h000010fc;  wr_data_rom[ 6724]='h00000000;
    rd_cycle[ 6725] = 1'b1;  wr_cycle[ 6725] = 1'b0;  addr_rom[ 6725]='h00002f00;  wr_data_rom[ 6725]='h00000000;
    rd_cycle[ 6726] = 1'b1;  wr_cycle[ 6726] = 1'b0;  addr_rom[ 6726]='h00002758;  wr_data_rom[ 6726]='h00000000;
    rd_cycle[ 6727] = 1'b1;  wr_cycle[ 6727] = 1'b0;  addr_rom[ 6727]='h000037e0;  wr_data_rom[ 6727]='h00000000;
    rd_cycle[ 6728] = 1'b0;  wr_cycle[ 6728] = 1'b1;  addr_rom[ 6728]='h000009d4;  wr_data_rom[ 6728]='h00002bee;
    rd_cycle[ 6729] = 1'b1;  wr_cycle[ 6729] = 1'b0;  addr_rom[ 6729]='h00002160;  wr_data_rom[ 6729]='h00000000;
    rd_cycle[ 6730] = 1'b1;  wr_cycle[ 6730] = 1'b0;  addr_rom[ 6730]='h00002ee8;  wr_data_rom[ 6730]='h00000000;
    rd_cycle[ 6731] = 1'b1;  wr_cycle[ 6731] = 1'b0;  addr_rom[ 6731]='h00001984;  wr_data_rom[ 6731]='h00000000;
    rd_cycle[ 6732] = 1'b1;  wr_cycle[ 6732] = 1'b0;  addr_rom[ 6732]='h00002ae0;  wr_data_rom[ 6732]='h00000000;
    rd_cycle[ 6733] = 1'b0;  wr_cycle[ 6733] = 1'b1;  addr_rom[ 6733]='h000031d8;  wr_data_rom[ 6733]='h00000a3e;
    rd_cycle[ 6734] = 1'b1;  wr_cycle[ 6734] = 1'b0;  addr_rom[ 6734]='h00001a64;  wr_data_rom[ 6734]='h00000000;
    rd_cycle[ 6735] = 1'b0;  wr_cycle[ 6735] = 1'b1;  addr_rom[ 6735]='h00003fc0;  wr_data_rom[ 6735]='h00003d80;
    rd_cycle[ 6736] = 1'b1;  wr_cycle[ 6736] = 1'b0;  addr_rom[ 6736]='h000003c8;  wr_data_rom[ 6736]='h00000000;
    rd_cycle[ 6737] = 1'b0;  wr_cycle[ 6737] = 1'b1;  addr_rom[ 6737]='h00001d40;  wr_data_rom[ 6737]='h00002d2e;
    rd_cycle[ 6738] = 1'b0;  wr_cycle[ 6738] = 1'b1;  addr_rom[ 6738]='h00002830;  wr_data_rom[ 6738]='h0000084d;
    rd_cycle[ 6739] = 1'b1;  wr_cycle[ 6739] = 1'b0;  addr_rom[ 6739]='h00003a04;  wr_data_rom[ 6739]='h00000000;
    rd_cycle[ 6740] = 1'b1;  wr_cycle[ 6740] = 1'b0;  addr_rom[ 6740]='h00003350;  wr_data_rom[ 6740]='h00000000;
    rd_cycle[ 6741] = 1'b0;  wr_cycle[ 6741] = 1'b1;  addr_rom[ 6741]='h000016c0;  wr_data_rom[ 6741]='h00000a42;
    rd_cycle[ 6742] = 1'b0;  wr_cycle[ 6742] = 1'b1;  addr_rom[ 6742]='h000026d4;  wr_data_rom[ 6742]='h00003bba;
    rd_cycle[ 6743] = 1'b0;  wr_cycle[ 6743] = 1'b1;  addr_rom[ 6743]='h000001f4;  wr_data_rom[ 6743]='h00003bc9;
    rd_cycle[ 6744] = 1'b0;  wr_cycle[ 6744] = 1'b1;  addr_rom[ 6744]='h00000de0;  wr_data_rom[ 6744]='h00001968;
    rd_cycle[ 6745] = 1'b1;  wr_cycle[ 6745] = 1'b0;  addr_rom[ 6745]='h00002c18;  wr_data_rom[ 6745]='h00000000;
    rd_cycle[ 6746] = 1'b0;  wr_cycle[ 6746] = 1'b1;  addr_rom[ 6746]='h00000398;  wr_data_rom[ 6746]='h00001e11;
    rd_cycle[ 6747] = 1'b0;  wr_cycle[ 6747] = 1'b1;  addr_rom[ 6747]='h00000db8;  wr_data_rom[ 6747]='h00000597;
    rd_cycle[ 6748] = 1'b1;  wr_cycle[ 6748] = 1'b0;  addr_rom[ 6748]='h000039d0;  wr_data_rom[ 6748]='h00000000;
    rd_cycle[ 6749] = 1'b1;  wr_cycle[ 6749] = 1'b0;  addr_rom[ 6749]='h000021f4;  wr_data_rom[ 6749]='h00000000;
    rd_cycle[ 6750] = 1'b1;  wr_cycle[ 6750] = 1'b0;  addr_rom[ 6750]='h0000021c;  wr_data_rom[ 6750]='h00000000;
    rd_cycle[ 6751] = 1'b0;  wr_cycle[ 6751] = 1'b1;  addr_rom[ 6751]='h00001fb0;  wr_data_rom[ 6751]='h0000037f;
    rd_cycle[ 6752] = 1'b1;  wr_cycle[ 6752] = 1'b0;  addr_rom[ 6752]='h0000112c;  wr_data_rom[ 6752]='h00000000;
    rd_cycle[ 6753] = 1'b0;  wr_cycle[ 6753] = 1'b1;  addr_rom[ 6753]='h00003128;  wr_data_rom[ 6753]='h00000601;
    rd_cycle[ 6754] = 1'b1;  wr_cycle[ 6754] = 1'b0;  addr_rom[ 6754]='h00002fa0;  wr_data_rom[ 6754]='h00000000;
    rd_cycle[ 6755] = 1'b1;  wr_cycle[ 6755] = 1'b0;  addr_rom[ 6755]='h00003834;  wr_data_rom[ 6755]='h00000000;
    rd_cycle[ 6756] = 1'b1;  wr_cycle[ 6756] = 1'b0;  addr_rom[ 6756]='h000001f8;  wr_data_rom[ 6756]='h00000000;
    rd_cycle[ 6757] = 1'b1;  wr_cycle[ 6757] = 1'b0;  addr_rom[ 6757]='h00000ddc;  wr_data_rom[ 6757]='h00000000;
    rd_cycle[ 6758] = 1'b1;  wr_cycle[ 6758] = 1'b0;  addr_rom[ 6758]='h00003410;  wr_data_rom[ 6758]='h00000000;
    rd_cycle[ 6759] = 1'b0;  wr_cycle[ 6759] = 1'b1;  addr_rom[ 6759]='h00001908;  wr_data_rom[ 6759]='h0000241a;
    rd_cycle[ 6760] = 1'b1;  wr_cycle[ 6760] = 1'b0;  addr_rom[ 6760]='h00001b9c;  wr_data_rom[ 6760]='h00000000;
    rd_cycle[ 6761] = 1'b1;  wr_cycle[ 6761] = 1'b0;  addr_rom[ 6761]='h00003540;  wr_data_rom[ 6761]='h00000000;
    rd_cycle[ 6762] = 1'b1;  wr_cycle[ 6762] = 1'b0;  addr_rom[ 6762]='h00001eec;  wr_data_rom[ 6762]='h00000000;
    rd_cycle[ 6763] = 1'b1;  wr_cycle[ 6763] = 1'b0;  addr_rom[ 6763]='h000006c0;  wr_data_rom[ 6763]='h00000000;
    rd_cycle[ 6764] = 1'b0;  wr_cycle[ 6764] = 1'b1;  addr_rom[ 6764]='h00000024;  wr_data_rom[ 6764]='h0000146b;
    rd_cycle[ 6765] = 1'b1;  wr_cycle[ 6765] = 1'b0;  addr_rom[ 6765]='h000039a4;  wr_data_rom[ 6765]='h00000000;
    rd_cycle[ 6766] = 1'b0;  wr_cycle[ 6766] = 1'b1;  addr_rom[ 6766]='h00000710;  wr_data_rom[ 6766]='h00002528;
    rd_cycle[ 6767] = 1'b1;  wr_cycle[ 6767] = 1'b0;  addr_rom[ 6767]='h00001168;  wr_data_rom[ 6767]='h00000000;
    rd_cycle[ 6768] = 1'b1;  wr_cycle[ 6768] = 1'b0;  addr_rom[ 6768]='h000025bc;  wr_data_rom[ 6768]='h00000000;
    rd_cycle[ 6769] = 1'b0;  wr_cycle[ 6769] = 1'b1;  addr_rom[ 6769]='h000030b8;  wr_data_rom[ 6769]='h00003481;
    rd_cycle[ 6770] = 1'b0;  wr_cycle[ 6770] = 1'b1;  addr_rom[ 6770]='h00002bc0;  wr_data_rom[ 6770]='h00000880;
    rd_cycle[ 6771] = 1'b0;  wr_cycle[ 6771] = 1'b1;  addr_rom[ 6771]='h000008fc;  wr_data_rom[ 6771]='h00000013;
    rd_cycle[ 6772] = 1'b0;  wr_cycle[ 6772] = 1'b1;  addr_rom[ 6772]='h00002288;  wr_data_rom[ 6772]='h00000cf6;
    rd_cycle[ 6773] = 1'b1;  wr_cycle[ 6773] = 1'b0;  addr_rom[ 6773]='h0000202c;  wr_data_rom[ 6773]='h00000000;
    rd_cycle[ 6774] = 1'b0;  wr_cycle[ 6774] = 1'b1;  addr_rom[ 6774]='h00002aa0;  wr_data_rom[ 6774]='h0000220d;
    rd_cycle[ 6775] = 1'b0;  wr_cycle[ 6775] = 1'b1;  addr_rom[ 6775]='h00000508;  wr_data_rom[ 6775]='h0000009d;
    rd_cycle[ 6776] = 1'b1;  wr_cycle[ 6776] = 1'b0;  addr_rom[ 6776]='h00001e08;  wr_data_rom[ 6776]='h00000000;
    rd_cycle[ 6777] = 1'b0;  wr_cycle[ 6777] = 1'b1;  addr_rom[ 6777]='h00001c9c;  wr_data_rom[ 6777]='h00003a93;
    rd_cycle[ 6778] = 1'b1;  wr_cycle[ 6778] = 1'b0;  addr_rom[ 6778]='h000015d0;  wr_data_rom[ 6778]='h00000000;
    rd_cycle[ 6779] = 1'b0;  wr_cycle[ 6779] = 1'b1;  addr_rom[ 6779]='h000035bc;  wr_data_rom[ 6779]='h0000049f;
    rd_cycle[ 6780] = 1'b1;  wr_cycle[ 6780] = 1'b0;  addr_rom[ 6780]='h00003390;  wr_data_rom[ 6780]='h00000000;
    rd_cycle[ 6781] = 1'b0;  wr_cycle[ 6781] = 1'b1;  addr_rom[ 6781]='h00001160;  wr_data_rom[ 6781]='h00001c5b;
    rd_cycle[ 6782] = 1'b0;  wr_cycle[ 6782] = 1'b1;  addr_rom[ 6782]='h00003708;  wr_data_rom[ 6782]='h00003250;
    rd_cycle[ 6783] = 1'b1;  wr_cycle[ 6783] = 1'b0;  addr_rom[ 6783]='h00001b30;  wr_data_rom[ 6783]='h00000000;
    rd_cycle[ 6784] = 1'b1;  wr_cycle[ 6784] = 1'b0;  addr_rom[ 6784]='h00003400;  wr_data_rom[ 6784]='h00000000;
    rd_cycle[ 6785] = 1'b1;  wr_cycle[ 6785] = 1'b0;  addr_rom[ 6785]='h00001d64;  wr_data_rom[ 6785]='h00000000;
    rd_cycle[ 6786] = 1'b0;  wr_cycle[ 6786] = 1'b1;  addr_rom[ 6786]='h000037c8;  wr_data_rom[ 6786]='h00002e25;
    rd_cycle[ 6787] = 1'b1;  wr_cycle[ 6787] = 1'b0;  addr_rom[ 6787]='h00003284;  wr_data_rom[ 6787]='h00000000;
    rd_cycle[ 6788] = 1'b0;  wr_cycle[ 6788] = 1'b1;  addr_rom[ 6788]='h00002fd0;  wr_data_rom[ 6788]='h000034dc;
    rd_cycle[ 6789] = 1'b0;  wr_cycle[ 6789] = 1'b1;  addr_rom[ 6789]='h0000126c;  wr_data_rom[ 6789]='h000037ed;
    rd_cycle[ 6790] = 1'b1;  wr_cycle[ 6790] = 1'b0;  addr_rom[ 6790]='h00000474;  wr_data_rom[ 6790]='h00000000;
    rd_cycle[ 6791] = 1'b0;  wr_cycle[ 6791] = 1'b1;  addr_rom[ 6791]='h000025ec;  wr_data_rom[ 6791]='h00003da8;
    rd_cycle[ 6792] = 1'b1;  wr_cycle[ 6792] = 1'b0;  addr_rom[ 6792]='h00003db8;  wr_data_rom[ 6792]='h00000000;
    rd_cycle[ 6793] = 1'b1;  wr_cycle[ 6793] = 1'b0;  addr_rom[ 6793]='h000031bc;  wr_data_rom[ 6793]='h00000000;
    rd_cycle[ 6794] = 1'b0;  wr_cycle[ 6794] = 1'b1;  addr_rom[ 6794]='h00002950;  wr_data_rom[ 6794]='h0000321b;
    rd_cycle[ 6795] = 1'b1;  wr_cycle[ 6795] = 1'b0;  addr_rom[ 6795]='h00002470;  wr_data_rom[ 6795]='h00000000;
    rd_cycle[ 6796] = 1'b1;  wr_cycle[ 6796] = 1'b0;  addr_rom[ 6796]='h000029c8;  wr_data_rom[ 6796]='h00000000;
    rd_cycle[ 6797] = 1'b0;  wr_cycle[ 6797] = 1'b1;  addr_rom[ 6797]='h0000246c;  wr_data_rom[ 6797]='h0000399b;
    rd_cycle[ 6798] = 1'b1;  wr_cycle[ 6798] = 1'b0;  addr_rom[ 6798]='h00002b68;  wr_data_rom[ 6798]='h00000000;
    rd_cycle[ 6799] = 1'b1;  wr_cycle[ 6799] = 1'b0;  addr_rom[ 6799]='h00003528;  wr_data_rom[ 6799]='h00000000;
    rd_cycle[ 6800] = 1'b0;  wr_cycle[ 6800] = 1'b1;  addr_rom[ 6800]='h00003fd0;  wr_data_rom[ 6800]='h00001884;
    rd_cycle[ 6801] = 1'b0;  wr_cycle[ 6801] = 1'b1;  addr_rom[ 6801]='h00003d14;  wr_data_rom[ 6801]='h0000268f;
    rd_cycle[ 6802] = 1'b1;  wr_cycle[ 6802] = 1'b0;  addr_rom[ 6802]='h0000155c;  wr_data_rom[ 6802]='h00000000;
    rd_cycle[ 6803] = 1'b1;  wr_cycle[ 6803] = 1'b0;  addr_rom[ 6803]='h000029d4;  wr_data_rom[ 6803]='h00000000;
    rd_cycle[ 6804] = 1'b0;  wr_cycle[ 6804] = 1'b1;  addr_rom[ 6804]='h000014f4;  wr_data_rom[ 6804]='h00003054;
    rd_cycle[ 6805] = 1'b1;  wr_cycle[ 6805] = 1'b0;  addr_rom[ 6805]='h000026cc;  wr_data_rom[ 6805]='h00000000;
    rd_cycle[ 6806] = 1'b0;  wr_cycle[ 6806] = 1'b1;  addr_rom[ 6806]='h0000250c;  wr_data_rom[ 6806]='h00000625;
    rd_cycle[ 6807] = 1'b1;  wr_cycle[ 6807] = 1'b0;  addr_rom[ 6807]='h00001758;  wr_data_rom[ 6807]='h00000000;
    rd_cycle[ 6808] = 1'b1;  wr_cycle[ 6808] = 1'b0;  addr_rom[ 6808]='h000016a4;  wr_data_rom[ 6808]='h00000000;
    rd_cycle[ 6809] = 1'b0;  wr_cycle[ 6809] = 1'b1;  addr_rom[ 6809]='h00003f8c;  wr_data_rom[ 6809]='h00002696;
    rd_cycle[ 6810] = 1'b0;  wr_cycle[ 6810] = 1'b1;  addr_rom[ 6810]='h000012d4;  wr_data_rom[ 6810]='h0000371b;
    rd_cycle[ 6811] = 1'b0;  wr_cycle[ 6811] = 1'b1;  addr_rom[ 6811]='h00001f40;  wr_data_rom[ 6811]='h000010c5;
    rd_cycle[ 6812] = 1'b1;  wr_cycle[ 6812] = 1'b0;  addr_rom[ 6812]='h00001260;  wr_data_rom[ 6812]='h00000000;
    rd_cycle[ 6813] = 1'b1;  wr_cycle[ 6813] = 1'b0;  addr_rom[ 6813]='h00000ae8;  wr_data_rom[ 6813]='h00000000;
    rd_cycle[ 6814] = 1'b1;  wr_cycle[ 6814] = 1'b0;  addr_rom[ 6814]='h00000ab8;  wr_data_rom[ 6814]='h00000000;
    rd_cycle[ 6815] = 1'b0;  wr_cycle[ 6815] = 1'b1;  addr_rom[ 6815]='h0000193c;  wr_data_rom[ 6815]='h0000052f;
    rd_cycle[ 6816] = 1'b1;  wr_cycle[ 6816] = 1'b0;  addr_rom[ 6816]='h00002d1c;  wr_data_rom[ 6816]='h00000000;
    rd_cycle[ 6817] = 1'b1;  wr_cycle[ 6817] = 1'b0;  addr_rom[ 6817]='h0000022c;  wr_data_rom[ 6817]='h00000000;
    rd_cycle[ 6818] = 1'b0;  wr_cycle[ 6818] = 1'b1;  addr_rom[ 6818]='h00003c4c;  wr_data_rom[ 6818]='h00003f13;
    rd_cycle[ 6819] = 1'b0;  wr_cycle[ 6819] = 1'b1;  addr_rom[ 6819]='h00000684;  wr_data_rom[ 6819]='h0000215c;
    rd_cycle[ 6820] = 1'b0;  wr_cycle[ 6820] = 1'b1;  addr_rom[ 6820]='h00000fa4;  wr_data_rom[ 6820]='h000037ba;
    rd_cycle[ 6821] = 1'b0;  wr_cycle[ 6821] = 1'b1;  addr_rom[ 6821]='h00001060;  wr_data_rom[ 6821]='h000006c1;
    rd_cycle[ 6822] = 1'b1;  wr_cycle[ 6822] = 1'b0;  addr_rom[ 6822]='h00001464;  wr_data_rom[ 6822]='h00000000;
    rd_cycle[ 6823] = 1'b0;  wr_cycle[ 6823] = 1'b1;  addr_rom[ 6823]='h0000210c;  wr_data_rom[ 6823]='h00001865;
    rd_cycle[ 6824] = 1'b0;  wr_cycle[ 6824] = 1'b1;  addr_rom[ 6824]='h00003cfc;  wr_data_rom[ 6824]='h000003f9;
    rd_cycle[ 6825] = 1'b0;  wr_cycle[ 6825] = 1'b1;  addr_rom[ 6825]='h00002c9c;  wr_data_rom[ 6825]='h00001311;
    rd_cycle[ 6826] = 1'b1;  wr_cycle[ 6826] = 1'b0;  addr_rom[ 6826]='h00003478;  wr_data_rom[ 6826]='h00000000;
    rd_cycle[ 6827] = 1'b1;  wr_cycle[ 6827] = 1'b0;  addr_rom[ 6827]='h0000182c;  wr_data_rom[ 6827]='h00000000;
    rd_cycle[ 6828] = 1'b0;  wr_cycle[ 6828] = 1'b1;  addr_rom[ 6828]='h00000f6c;  wr_data_rom[ 6828]='h0000162b;
    rd_cycle[ 6829] = 1'b0;  wr_cycle[ 6829] = 1'b1;  addr_rom[ 6829]='h000003bc;  wr_data_rom[ 6829]='h00003033;
    rd_cycle[ 6830] = 1'b1;  wr_cycle[ 6830] = 1'b0;  addr_rom[ 6830]='h00002974;  wr_data_rom[ 6830]='h00000000;
    rd_cycle[ 6831] = 1'b1;  wr_cycle[ 6831] = 1'b0;  addr_rom[ 6831]='h00001514;  wr_data_rom[ 6831]='h00000000;
    rd_cycle[ 6832] = 1'b0;  wr_cycle[ 6832] = 1'b1;  addr_rom[ 6832]='h00002054;  wr_data_rom[ 6832]='h00002523;
    rd_cycle[ 6833] = 1'b0;  wr_cycle[ 6833] = 1'b1;  addr_rom[ 6833]='h00000f64;  wr_data_rom[ 6833]='h000017fe;
    rd_cycle[ 6834] = 1'b1;  wr_cycle[ 6834] = 1'b0;  addr_rom[ 6834]='h00003774;  wr_data_rom[ 6834]='h00000000;
    rd_cycle[ 6835] = 1'b0;  wr_cycle[ 6835] = 1'b1;  addr_rom[ 6835]='h00000374;  wr_data_rom[ 6835]='h00000d0c;
    rd_cycle[ 6836] = 1'b0;  wr_cycle[ 6836] = 1'b1;  addr_rom[ 6836]='h00000798;  wr_data_rom[ 6836]='h00002b52;
    rd_cycle[ 6837] = 1'b1;  wr_cycle[ 6837] = 1'b0;  addr_rom[ 6837]='h00003394;  wr_data_rom[ 6837]='h00000000;
    rd_cycle[ 6838] = 1'b1;  wr_cycle[ 6838] = 1'b0;  addr_rom[ 6838]='h00002014;  wr_data_rom[ 6838]='h00000000;
    rd_cycle[ 6839] = 1'b1;  wr_cycle[ 6839] = 1'b0;  addr_rom[ 6839]='h00002760;  wr_data_rom[ 6839]='h00000000;
    rd_cycle[ 6840] = 1'b1;  wr_cycle[ 6840] = 1'b0;  addr_rom[ 6840]='h0000331c;  wr_data_rom[ 6840]='h00000000;
    rd_cycle[ 6841] = 1'b1;  wr_cycle[ 6841] = 1'b0;  addr_rom[ 6841]='h00003814;  wr_data_rom[ 6841]='h00000000;
    rd_cycle[ 6842] = 1'b1;  wr_cycle[ 6842] = 1'b0;  addr_rom[ 6842]='h00000278;  wr_data_rom[ 6842]='h00000000;
    rd_cycle[ 6843] = 1'b1;  wr_cycle[ 6843] = 1'b0;  addr_rom[ 6843]='h00000770;  wr_data_rom[ 6843]='h00000000;
    rd_cycle[ 6844] = 1'b0;  wr_cycle[ 6844] = 1'b1;  addr_rom[ 6844]='h00003720;  wr_data_rom[ 6844]='h0000092c;
    rd_cycle[ 6845] = 1'b1;  wr_cycle[ 6845] = 1'b0;  addr_rom[ 6845]='h0000284c;  wr_data_rom[ 6845]='h00000000;
    rd_cycle[ 6846] = 1'b1;  wr_cycle[ 6846] = 1'b0;  addr_rom[ 6846]='h00000f54;  wr_data_rom[ 6846]='h00000000;
    rd_cycle[ 6847] = 1'b1;  wr_cycle[ 6847] = 1'b0;  addr_rom[ 6847]='h00003084;  wr_data_rom[ 6847]='h00000000;
    rd_cycle[ 6848] = 1'b1;  wr_cycle[ 6848] = 1'b0;  addr_rom[ 6848]='h00000e78;  wr_data_rom[ 6848]='h00000000;
    rd_cycle[ 6849] = 1'b0;  wr_cycle[ 6849] = 1'b1;  addr_rom[ 6849]='h00002ec4;  wr_data_rom[ 6849]='h000013ac;
    rd_cycle[ 6850] = 1'b0;  wr_cycle[ 6850] = 1'b1;  addr_rom[ 6850]='h00003b30;  wr_data_rom[ 6850]='h00000dcb;
    rd_cycle[ 6851] = 1'b1;  wr_cycle[ 6851] = 1'b0;  addr_rom[ 6851]='h00003e8c;  wr_data_rom[ 6851]='h00000000;
    rd_cycle[ 6852] = 1'b0;  wr_cycle[ 6852] = 1'b1;  addr_rom[ 6852]='h00002768;  wr_data_rom[ 6852]='h00000b25;
    rd_cycle[ 6853] = 1'b1;  wr_cycle[ 6853] = 1'b0;  addr_rom[ 6853]='h0000345c;  wr_data_rom[ 6853]='h00000000;
    rd_cycle[ 6854] = 1'b0;  wr_cycle[ 6854] = 1'b1;  addr_rom[ 6854]='h000012f4;  wr_data_rom[ 6854]='h0000114e;
    rd_cycle[ 6855] = 1'b1;  wr_cycle[ 6855] = 1'b0;  addr_rom[ 6855]='h00000fe4;  wr_data_rom[ 6855]='h00000000;
    rd_cycle[ 6856] = 1'b0;  wr_cycle[ 6856] = 1'b1;  addr_rom[ 6856]='h00002548;  wr_data_rom[ 6856]='h000023d2;
    rd_cycle[ 6857] = 1'b0;  wr_cycle[ 6857] = 1'b1;  addr_rom[ 6857]='h0000185c;  wr_data_rom[ 6857]='h00001f25;
    rd_cycle[ 6858] = 1'b0;  wr_cycle[ 6858] = 1'b1;  addr_rom[ 6858]='h000016e8;  wr_data_rom[ 6858]='h00000532;
    rd_cycle[ 6859] = 1'b0;  wr_cycle[ 6859] = 1'b1;  addr_rom[ 6859]='h000007d4;  wr_data_rom[ 6859]='h0000025c;
    rd_cycle[ 6860] = 1'b0;  wr_cycle[ 6860] = 1'b1;  addr_rom[ 6860]='h000039f4;  wr_data_rom[ 6860]='h00002905;
    rd_cycle[ 6861] = 1'b1;  wr_cycle[ 6861] = 1'b0;  addr_rom[ 6861]='h00002988;  wr_data_rom[ 6861]='h00000000;
    rd_cycle[ 6862] = 1'b0;  wr_cycle[ 6862] = 1'b1;  addr_rom[ 6862]='h000035c0;  wr_data_rom[ 6862]='h00002428;
    rd_cycle[ 6863] = 1'b0;  wr_cycle[ 6863] = 1'b1;  addr_rom[ 6863]='h00002694;  wr_data_rom[ 6863]='h0000214a;
    rd_cycle[ 6864] = 1'b0;  wr_cycle[ 6864] = 1'b1;  addr_rom[ 6864]='h00003000;  wr_data_rom[ 6864]='h00000eec;
    rd_cycle[ 6865] = 1'b0;  wr_cycle[ 6865] = 1'b1;  addr_rom[ 6865]='h00000af4;  wr_data_rom[ 6865]='h00002356;
    rd_cycle[ 6866] = 1'b1;  wr_cycle[ 6866] = 1'b0;  addr_rom[ 6866]='h00000b68;  wr_data_rom[ 6866]='h00000000;
    rd_cycle[ 6867] = 1'b1;  wr_cycle[ 6867] = 1'b0;  addr_rom[ 6867]='h000020dc;  wr_data_rom[ 6867]='h00000000;
    rd_cycle[ 6868] = 1'b0;  wr_cycle[ 6868] = 1'b1;  addr_rom[ 6868]='h00001584;  wr_data_rom[ 6868]='h00003e20;
    rd_cycle[ 6869] = 1'b0;  wr_cycle[ 6869] = 1'b1;  addr_rom[ 6869]='h000027d8;  wr_data_rom[ 6869]='h00003416;
    rd_cycle[ 6870] = 1'b1;  wr_cycle[ 6870] = 1'b0;  addr_rom[ 6870]='h00000c38;  wr_data_rom[ 6870]='h00000000;
    rd_cycle[ 6871] = 1'b1;  wr_cycle[ 6871] = 1'b0;  addr_rom[ 6871]='h0000365c;  wr_data_rom[ 6871]='h00000000;
    rd_cycle[ 6872] = 1'b0;  wr_cycle[ 6872] = 1'b1;  addr_rom[ 6872]='h00003104;  wr_data_rom[ 6872]='h00003e6d;
    rd_cycle[ 6873] = 1'b0;  wr_cycle[ 6873] = 1'b1;  addr_rom[ 6873]='h000011a8;  wr_data_rom[ 6873]='h000036d2;
    rd_cycle[ 6874] = 1'b1;  wr_cycle[ 6874] = 1'b0;  addr_rom[ 6874]='h000008c8;  wr_data_rom[ 6874]='h00000000;
    rd_cycle[ 6875] = 1'b0;  wr_cycle[ 6875] = 1'b1;  addr_rom[ 6875]='h00000c2c;  wr_data_rom[ 6875]='h000014cf;
    rd_cycle[ 6876] = 1'b1;  wr_cycle[ 6876] = 1'b0;  addr_rom[ 6876]='h00001188;  wr_data_rom[ 6876]='h00000000;
    rd_cycle[ 6877] = 1'b1;  wr_cycle[ 6877] = 1'b0;  addr_rom[ 6877]='h00000c9c;  wr_data_rom[ 6877]='h00000000;
    rd_cycle[ 6878] = 1'b0;  wr_cycle[ 6878] = 1'b1;  addr_rom[ 6878]='h000026ec;  wr_data_rom[ 6878]='h00001141;
    rd_cycle[ 6879] = 1'b0;  wr_cycle[ 6879] = 1'b1;  addr_rom[ 6879]='h000031a4;  wr_data_rom[ 6879]='h000010a7;
    rd_cycle[ 6880] = 1'b0;  wr_cycle[ 6880] = 1'b1;  addr_rom[ 6880]='h00003288;  wr_data_rom[ 6880]='h00002484;
    rd_cycle[ 6881] = 1'b0;  wr_cycle[ 6881] = 1'b1;  addr_rom[ 6881]='h00002470;  wr_data_rom[ 6881]='h00000976;
    rd_cycle[ 6882] = 1'b0;  wr_cycle[ 6882] = 1'b1;  addr_rom[ 6882]='h0000186c;  wr_data_rom[ 6882]='h00002f20;
    rd_cycle[ 6883] = 1'b1;  wr_cycle[ 6883] = 1'b0;  addr_rom[ 6883]='h000024f4;  wr_data_rom[ 6883]='h00000000;
    rd_cycle[ 6884] = 1'b1;  wr_cycle[ 6884] = 1'b0;  addr_rom[ 6884]='h00000200;  wr_data_rom[ 6884]='h00000000;
    rd_cycle[ 6885] = 1'b0;  wr_cycle[ 6885] = 1'b1;  addr_rom[ 6885]='h00001d50;  wr_data_rom[ 6885]='h0000364c;
    rd_cycle[ 6886] = 1'b1;  wr_cycle[ 6886] = 1'b0;  addr_rom[ 6886]='h00003744;  wr_data_rom[ 6886]='h00000000;
    rd_cycle[ 6887] = 1'b0;  wr_cycle[ 6887] = 1'b1;  addr_rom[ 6887]='h00003eb8;  wr_data_rom[ 6887]='h000015a2;
    rd_cycle[ 6888] = 1'b1;  wr_cycle[ 6888] = 1'b0;  addr_rom[ 6888]='h00000dcc;  wr_data_rom[ 6888]='h00000000;
    rd_cycle[ 6889] = 1'b0;  wr_cycle[ 6889] = 1'b1;  addr_rom[ 6889]='h000009f0;  wr_data_rom[ 6889]='h00002296;
    rd_cycle[ 6890] = 1'b1;  wr_cycle[ 6890] = 1'b0;  addr_rom[ 6890]='h00002f34;  wr_data_rom[ 6890]='h00000000;
    rd_cycle[ 6891] = 1'b1;  wr_cycle[ 6891] = 1'b0;  addr_rom[ 6891]='h00003eb0;  wr_data_rom[ 6891]='h00000000;
    rd_cycle[ 6892] = 1'b1;  wr_cycle[ 6892] = 1'b0;  addr_rom[ 6892]='h0000306c;  wr_data_rom[ 6892]='h00000000;
    rd_cycle[ 6893] = 1'b1;  wr_cycle[ 6893] = 1'b0;  addr_rom[ 6893]='h00002cd0;  wr_data_rom[ 6893]='h00000000;
    rd_cycle[ 6894] = 1'b0;  wr_cycle[ 6894] = 1'b1;  addr_rom[ 6894]='h00000f78;  wr_data_rom[ 6894]='h0000304d;
    rd_cycle[ 6895] = 1'b0;  wr_cycle[ 6895] = 1'b1;  addr_rom[ 6895]='h00000388;  wr_data_rom[ 6895]='h00000936;
    rd_cycle[ 6896] = 1'b0;  wr_cycle[ 6896] = 1'b1;  addr_rom[ 6896]='h00000bc8;  wr_data_rom[ 6896]='h000009f4;
    rd_cycle[ 6897] = 1'b1;  wr_cycle[ 6897] = 1'b0;  addr_rom[ 6897]='h00001b0c;  wr_data_rom[ 6897]='h00000000;
    rd_cycle[ 6898] = 1'b1;  wr_cycle[ 6898] = 1'b0;  addr_rom[ 6898]='h00000d00;  wr_data_rom[ 6898]='h00000000;
    rd_cycle[ 6899] = 1'b0;  wr_cycle[ 6899] = 1'b1;  addr_rom[ 6899]='h00001c9c;  wr_data_rom[ 6899]='h00001d46;
    rd_cycle[ 6900] = 1'b0;  wr_cycle[ 6900] = 1'b1;  addr_rom[ 6900]='h00000470;  wr_data_rom[ 6900]='h0000090f;
    rd_cycle[ 6901] = 1'b0;  wr_cycle[ 6901] = 1'b1;  addr_rom[ 6901]='h00001538;  wr_data_rom[ 6901]='h00001888;
    rd_cycle[ 6902] = 1'b1;  wr_cycle[ 6902] = 1'b0;  addr_rom[ 6902]='h00001470;  wr_data_rom[ 6902]='h00000000;
    rd_cycle[ 6903] = 1'b1;  wr_cycle[ 6903] = 1'b0;  addr_rom[ 6903]='h00003400;  wr_data_rom[ 6903]='h00000000;
    rd_cycle[ 6904] = 1'b1;  wr_cycle[ 6904] = 1'b0;  addr_rom[ 6904]='h000034c4;  wr_data_rom[ 6904]='h00000000;
    rd_cycle[ 6905] = 1'b0;  wr_cycle[ 6905] = 1'b1;  addr_rom[ 6905]='h000037a8;  wr_data_rom[ 6905]='h00001e55;
    rd_cycle[ 6906] = 1'b0;  wr_cycle[ 6906] = 1'b1;  addr_rom[ 6906]='h000002c4;  wr_data_rom[ 6906]='h0000397b;
    rd_cycle[ 6907] = 1'b1;  wr_cycle[ 6907] = 1'b0;  addr_rom[ 6907]='h00003528;  wr_data_rom[ 6907]='h00000000;
    rd_cycle[ 6908] = 1'b1;  wr_cycle[ 6908] = 1'b0;  addr_rom[ 6908]='h000018f4;  wr_data_rom[ 6908]='h00000000;
    rd_cycle[ 6909] = 1'b1;  wr_cycle[ 6909] = 1'b0;  addr_rom[ 6909]='h00001a04;  wr_data_rom[ 6909]='h00000000;
    rd_cycle[ 6910] = 1'b1;  wr_cycle[ 6910] = 1'b0;  addr_rom[ 6910]='h00001788;  wr_data_rom[ 6910]='h00000000;
    rd_cycle[ 6911] = 1'b1;  wr_cycle[ 6911] = 1'b0;  addr_rom[ 6911]='h00000b14;  wr_data_rom[ 6911]='h00000000;
    rd_cycle[ 6912] = 1'b1;  wr_cycle[ 6912] = 1'b0;  addr_rom[ 6912]='h00003d0c;  wr_data_rom[ 6912]='h00000000;
    rd_cycle[ 6913] = 1'b0;  wr_cycle[ 6913] = 1'b1;  addr_rom[ 6913]='h000007ac;  wr_data_rom[ 6913]='h000008f3;
    rd_cycle[ 6914] = 1'b0;  wr_cycle[ 6914] = 1'b1;  addr_rom[ 6914]='h000027b0;  wr_data_rom[ 6914]='h00001d8f;
    rd_cycle[ 6915] = 1'b0;  wr_cycle[ 6915] = 1'b1;  addr_rom[ 6915]='h00002fcc;  wr_data_rom[ 6915]='h000016c7;
    rd_cycle[ 6916] = 1'b1;  wr_cycle[ 6916] = 1'b0;  addr_rom[ 6916]='h00001eb8;  wr_data_rom[ 6916]='h00000000;
    rd_cycle[ 6917] = 1'b1;  wr_cycle[ 6917] = 1'b0;  addr_rom[ 6917]='h00002ec0;  wr_data_rom[ 6917]='h00000000;
    rd_cycle[ 6918] = 1'b0;  wr_cycle[ 6918] = 1'b1;  addr_rom[ 6918]='h00001278;  wr_data_rom[ 6918]='h00002047;
    rd_cycle[ 6919] = 1'b1;  wr_cycle[ 6919] = 1'b0;  addr_rom[ 6919]='h00003824;  wr_data_rom[ 6919]='h00000000;
    rd_cycle[ 6920] = 1'b1;  wr_cycle[ 6920] = 1'b0;  addr_rom[ 6920]='h00003c08;  wr_data_rom[ 6920]='h00000000;
    rd_cycle[ 6921] = 1'b0;  wr_cycle[ 6921] = 1'b1;  addr_rom[ 6921]='h00002750;  wr_data_rom[ 6921]='h00001c82;
    rd_cycle[ 6922] = 1'b1;  wr_cycle[ 6922] = 1'b0;  addr_rom[ 6922]='h00001820;  wr_data_rom[ 6922]='h00000000;
    rd_cycle[ 6923] = 1'b0;  wr_cycle[ 6923] = 1'b1;  addr_rom[ 6923]='h0000001c;  wr_data_rom[ 6923]='h00003287;
    rd_cycle[ 6924] = 1'b0;  wr_cycle[ 6924] = 1'b1;  addr_rom[ 6924]='h000009f4;  wr_data_rom[ 6924]='h00002e54;
    rd_cycle[ 6925] = 1'b0;  wr_cycle[ 6925] = 1'b1;  addr_rom[ 6925]='h0000342c;  wr_data_rom[ 6925]='h0000057c;
    rd_cycle[ 6926] = 1'b1;  wr_cycle[ 6926] = 1'b0;  addr_rom[ 6926]='h000013c8;  wr_data_rom[ 6926]='h00000000;
    rd_cycle[ 6927] = 1'b0;  wr_cycle[ 6927] = 1'b1;  addr_rom[ 6927]='h0000364c;  wr_data_rom[ 6927]='h0000036b;
    rd_cycle[ 6928] = 1'b1;  wr_cycle[ 6928] = 1'b0;  addr_rom[ 6928]='h00002968;  wr_data_rom[ 6928]='h00000000;
    rd_cycle[ 6929] = 1'b0;  wr_cycle[ 6929] = 1'b1;  addr_rom[ 6929]='h00000918;  wr_data_rom[ 6929]='h00002533;
    rd_cycle[ 6930] = 1'b0;  wr_cycle[ 6930] = 1'b1;  addr_rom[ 6930]='h00001880;  wr_data_rom[ 6930]='h00002df3;
    rd_cycle[ 6931] = 1'b1;  wr_cycle[ 6931] = 1'b0;  addr_rom[ 6931]='h00002b3c;  wr_data_rom[ 6931]='h00000000;
    rd_cycle[ 6932] = 1'b1;  wr_cycle[ 6932] = 1'b0;  addr_rom[ 6932]='h00003a5c;  wr_data_rom[ 6932]='h00000000;
    rd_cycle[ 6933] = 1'b1;  wr_cycle[ 6933] = 1'b0;  addr_rom[ 6933]='h00001bd0;  wr_data_rom[ 6933]='h00000000;
    rd_cycle[ 6934] = 1'b1;  wr_cycle[ 6934] = 1'b0;  addr_rom[ 6934]='h00001afc;  wr_data_rom[ 6934]='h00000000;
    rd_cycle[ 6935] = 1'b1;  wr_cycle[ 6935] = 1'b0;  addr_rom[ 6935]='h0000268c;  wr_data_rom[ 6935]='h00000000;
    rd_cycle[ 6936] = 1'b1;  wr_cycle[ 6936] = 1'b0;  addr_rom[ 6936]='h000000a0;  wr_data_rom[ 6936]='h00000000;
    rd_cycle[ 6937] = 1'b0;  wr_cycle[ 6937] = 1'b1;  addr_rom[ 6937]='h00003ab4;  wr_data_rom[ 6937]='h00003ff3;
    rd_cycle[ 6938] = 1'b0;  wr_cycle[ 6938] = 1'b1;  addr_rom[ 6938]='h00003b94;  wr_data_rom[ 6938]='h00002a02;
    rd_cycle[ 6939] = 1'b0;  wr_cycle[ 6939] = 1'b1;  addr_rom[ 6939]='h00001de8;  wr_data_rom[ 6939]='h00003112;
    rd_cycle[ 6940] = 1'b0;  wr_cycle[ 6940] = 1'b1;  addr_rom[ 6940]='h000009d8;  wr_data_rom[ 6940]='h000025f4;
    rd_cycle[ 6941] = 1'b1;  wr_cycle[ 6941] = 1'b0;  addr_rom[ 6941]='h0000012c;  wr_data_rom[ 6941]='h00000000;
    rd_cycle[ 6942] = 1'b0;  wr_cycle[ 6942] = 1'b1;  addr_rom[ 6942]='h00000e58;  wr_data_rom[ 6942]='h00002491;
    rd_cycle[ 6943] = 1'b0;  wr_cycle[ 6943] = 1'b1;  addr_rom[ 6943]='h00003a7c;  wr_data_rom[ 6943]='h00002575;
    rd_cycle[ 6944] = 1'b1;  wr_cycle[ 6944] = 1'b0;  addr_rom[ 6944]='h00000e78;  wr_data_rom[ 6944]='h00000000;
    rd_cycle[ 6945] = 1'b0;  wr_cycle[ 6945] = 1'b1;  addr_rom[ 6945]='h0000166c;  wr_data_rom[ 6945]='h00002f4a;
    rd_cycle[ 6946] = 1'b1;  wr_cycle[ 6946] = 1'b0;  addr_rom[ 6946]='h00003660;  wr_data_rom[ 6946]='h00000000;
    rd_cycle[ 6947] = 1'b0;  wr_cycle[ 6947] = 1'b1;  addr_rom[ 6947]='h0000040c;  wr_data_rom[ 6947]='h0000171a;
    rd_cycle[ 6948] = 1'b1;  wr_cycle[ 6948] = 1'b0;  addr_rom[ 6948]='h00001b8c;  wr_data_rom[ 6948]='h00000000;
    rd_cycle[ 6949] = 1'b1;  wr_cycle[ 6949] = 1'b0;  addr_rom[ 6949]='h000024f8;  wr_data_rom[ 6949]='h00000000;
    rd_cycle[ 6950] = 1'b0;  wr_cycle[ 6950] = 1'b1;  addr_rom[ 6950]='h000013c0;  wr_data_rom[ 6950]='h000037db;
    rd_cycle[ 6951] = 1'b0;  wr_cycle[ 6951] = 1'b1;  addr_rom[ 6951]='h00000b10;  wr_data_rom[ 6951]='h000036a8;
    rd_cycle[ 6952] = 1'b1;  wr_cycle[ 6952] = 1'b0;  addr_rom[ 6952]='h00000334;  wr_data_rom[ 6952]='h00000000;
    rd_cycle[ 6953] = 1'b1;  wr_cycle[ 6953] = 1'b0;  addr_rom[ 6953]='h00000498;  wr_data_rom[ 6953]='h00000000;
    rd_cycle[ 6954] = 1'b0;  wr_cycle[ 6954] = 1'b1;  addr_rom[ 6954]='h0000238c;  wr_data_rom[ 6954]='h00002901;
    rd_cycle[ 6955] = 1'b1;  wr_cycle[ 6955] = 1'b0;  addr_rom[ 6955]='h000006a0;  wr_data_rom[ 6955]='h00000000;
    rd_cycle[ 6956] = 1'b0;  wr_cycle[ 6956] = 1'b1;  addr_rom[ 6956]='h0000385c;  wr_data_rom[ 6956]='h00001526;
    rd_cycle[ 6957] = 1'b1;  wr_cycle[ 6957] = 1'b0;  addr_rom[ 6957]='h00003ad4;  wr_data_rom[ 6957]='h00000000;
    rd_cycle[ 6958] = 1'b0;  wr_cycle[ 6958] = 1'b1;  addr_rom[ 6958]='h00003890;  wr_data_rom[ 6958]='h00001690;
    rd_cycle[ 6959] = 1'b0;  wr_cycle[ 6959] = 1'b1;  addr_rom[ 6959]='h00002b54;  wr_data_rom[ 6959]='h00001114;
    rd_cycle[ 6960] = 1'b1;  wr_cycle[ 6960] = 1'b0;  addr_rom[ 6960]='h000031c8;  wr_data_rom[ 6960]='h00000000;
    rd_cycle[ 6961] = 1'b1;  wr_cycle[ 6961] = 1'b0;  addr_rom[ 6961]='h00001ffc;  wr_data_rom[ 6961]='h00000000;
    rd_cycle[ 6962] = 1'b1;  wr_cycle[ 6962] = 1'b0;  addr_rom[ 6962]='h00001f3c;  wr_data_rom[ 6962]='h00000000;
    rd_cycle[ 6963] = 1'b1;  wr_cycle[ 6963] = 1'b0;  addr_rom[ 6963]='h000025d8;  wr_data_rom[ 6963]='h00000000;
    rd_cycle[ 6964] = 1'b0;  wr_cycle[ 6964] = 1'b1;  addr_rom[ 6964]='h00001e10;  wr_data_rom[ 6964]='h00000bef;
    rd_cycle[ 6965] = 1'b1;  wr_cycle[ 6965] = 1'b0;  addr_rom[ 6965]='h00003808;  wr_data_rom[ 6965]='h00000000;
    rd_cycle[ 6966] = 1'b0;  wr_cycle[ 6966] = 1'b1;  addr_rom[ 6966]='h00002624;  wr_data_rom[ 6966]='h00002eb0;
    rd_cycle[ 6967] = 1'b0;  wr_cycle[ 6967] = 1'b1;  addr_rom[ 6967]='h00003944;  wr_data_rom[ 6967]='h000013ab;
    rd_cycle[ 6968] = 1'b1;  wr_cycle[ 6968] = 1'b0;  addr_rom[ 6968]='h00002160;  wr_data_rom[ 6968]='h00000000;
    rd_cycle[ 6969] = 1'b1;  wr_cycle[ 6969] = 1'b0;  addr_rom[ 6969]='h00003398;  wr_data_rom[ 6969]='h00000000;
    rd_cycle[ 6970] = 1'b1;  wr_cycle[ 6970] = 1'b0;  addr_rom[ 6970]='h00001570;  wr_data_rom[ 6970]='h00000000;
    rd_cycle[ 6971] = 1'b0;  wr_cycle[ 6971] = 1'b1;  addr_rom[ 6971]='h0000315c;  wr_data_rom[ 6971]='h00001a2d;
    rd_cycle[ 6972] = 1'b0;  wr_cycle[ 6972] = 1'b1;  addr_rom[ 6972]='h00003398;  wr_data_rom[ 6972]='h00002d94;
    rd_cycle[ 6973] = 1'b0;  wr_cycle[ 6973] = 1'b1;  addr_rom[ 6973]='h0000263c;  wr_data_rom[ 6973]='h00000641;
    rd_cycle[ 6974] = 1'b0;  wr_cycle[ 6974] = 1'b1;  addr_rom[ 6974]='h00002c94;  wr_data_rom[ 6974]='h00000f44;
    rd_cycle[ 6975] = 1'b1;  wr_cycle[ 6975] = 1'b0;  addr_rom[ 6975]='h00001304;  wr_data_rom[ 6975]='h00000000;
    rd_cycle[ 6976] = 1'b1;  wr_cycle[ 6976] = 1'b0;  addr_rom[ 6976]='h00001ba0;  wr_data_rom[ 6976]='h00000000;
    rd_cycle[ 6977] = 1'b0;  wr_cycle[ 6977] = 1'b1;  addr_rom[ 6977]='h00003d10;  wr_data_rom[ 6977]='h000037b6;
    rd_cycle[ 6978] = 1'b0;  wr_cycle[ 6978] = 1'b1;  addr_rom[ 6978]='h00003768;  wr_data_rom[ 6978]='h00000f22;
    rd_cycle[ 6979] = 1'b1;  wr_cycle[ 6979] = 1'b0;  addr_rom[ 6979]='h00000ab8;  wr_data_rom[ 6979]='h00000000;
    rd_cycle[ 6980] = 1'b0;  wr_cycle[ 6980] = 1'b1;  addr_rom[ 6980]='h00000588;  wr_data_rom[ 6980]='h00002d23;
    rd_cycle[ 6981] = 1'b1;  wr_cycle[ 6981] = 1'b0;  addr_rom[ 6981]='h00002e20;  wr_data_rom[ 6981]='h00000000;
    rd_cycle[ 6982] = 1'b1;  wr_cycle[ 6982] = 1'b0;  addr_rom[ 6982]='h00000130;  wr_data_rom[ 6982]='h00000000;
    rd_cycle[ 6983] = 1'b1;  wr_cycle[ 6983] = 1'b0;  addr_rom[ 6983]='h00000dac;  wr_data_rom[ 6983]='h00000000;
    rd_cycle[ 6984] = 1'b1;  wr_cycle[ 6984] = 1'b0;  addr_rom[ 6984]='h000016fc;  wr_data_rom[ 6984]='h00000000;
    rd_cycle[ 6985] = 1'b0;  wr_cycle[ 6985] = 1'b1;  addr_rom[ 6985]='h00003bcc;  wr_data_rom[ 6985]='h00000696;
    rd_cycle[ 6986] = 1'b0;  wr_cycle[ 6986] = 1'b1;  addr_rom[ 6986]='h0000161c;  wr_data_rom[ 6986]='h0000071f;
    rd_cycle[ 6987] = 1'b1;  wr_cycle[ 6987] = 1'b0;  addr_rom[ 6987]='h000001dc;  wr_data_rom[ 6987]='h00000000;
    rd_cycle[ 6988] = 1'b1;  wr_cycle[ 6988] = 1'b0;  addr_rom[ 6988]='h000016a8;  wr_data_rom[ 6988]='h00000000;
    rd_cycle[ 6989] = 1'b1;  wr_cycle[ 6989] = 1'b0;  addr_rom[ 6989]='h00000a90;  wr_data_rom[ 6989]='h00000000;
    rd_cycle[ 6990] = 1'b1;  wr_cycle[ 6990] = 1'b0;  addr_rom[ 6990]='h0000168c;  wr_data_rom[ 6990]='h00000000;
    rd_cycle[ 6991] = 1'b1;  wr_cycle[ 6991] = 1'b0;  addr_rom[ 6991]='h000017d8;  wr_data_rom[ 6991]='h00000000;
    rd_cycle[ 6992] = 1'b1;  wr_cycle[ 6992] = 1'b0;  addr_rom[ 6992]='h00003170;  wr_data_rom[ 6992]='h00000000;
    rd_cycle[ 6993] = 1'b1;  wr_cycle[ 6993] = 1'b0;  addr_rom[ 6993]='h0000120c;  wr_data_rom[ 6993]='h00000000;
    rd_cycle[ 6994] = 1'b0;  wr_cycle[ 6994] = 1'b1;  addr_rom[ 6994]='h00002c04;  wr_data_rom[ 6994]='h0000223b;
    rd_cycle[ 6995] = 1'b0;  wr_cycle[ 6995] = 1'b1;  addr_rom[ 6995]='h000004a0;  wr_data_rom[ 6995]='h00000169;
    rd_cycle[ 6996] = 1'b1;  wr_cycle[ 6996] = 1'b0;  addr_rom[ 6996]='h00001f5c;  wr_data_rom[ 6996]='h00000000;
    rd_cycle[ 6997] = 1'b0;  wr_cycle[ 6997] = 1'b1;  addr_rom[ 6997]='h00003e64;  wr_data_rom[ 6997]='h0000155c;
    rd_cycle[ 6998] = 1'b0;  wr_cycle[ 6998] = 1'b1;  addr_rom[ 6998]='h000009b4;  wr_data_rom[ 6998]='h00002126;
    rd_cycle[ 6999] = 1'b0;  wr_cycle[ 6999] = 1'b1;  addr_rom[ 6999]='h00002168;  wr_data_rom[ 6999]='h00001f88;
    rd_cycle[ 7000] = 1'b0;  wr_cycle[ 7000] = 1'b1;  addr_rom[ 7000]='h00003eec;  wr_data_rom[ 7000]='h00002269;
    rd_cycle[ 7001] = 1'b0;  wr_cycle[ 7001] = 1'b1;  addr_rom[ 7001]='h00003a10;  wr_data_rom[ 7001]='h00003973;
    rd_cycle[ 7002] = 1'b1;  wr_cycle[ 7002] = 1'b0;  addr_rom[ 7002]='h0000232c;  wr_data_rom[ 7002]='h00000000;
    rd_cycle[ 7003] = 1'b0;  wr_cycle[ 7003] = 1'b1;  addr_rom[ 7003]='h000007b8;  wr_data_rom[ 7003]='h00001666;
    rd_cycle[ 7004] = 1'b1;  wr_cycle[ 7004] = 1'b0;  addr_rom[ 7004]='h00002e10;  wr_data_rom[ 7004]='h00000000;
    rd_cycle[ 7005] = 1'b0;  wr_cycle[ 7005] = 1'b1;  addr_rom[ 7005]='h000023b8;  wr_data_rom[ 7005]='h000036be;
    rd_cycle[ 7006] = 1'b0;  wr_cycle[ 7006] = 1'b1;  addr_rom[ 7006]='h00000c9c;  wr_data_rom[ 7006]='h0000003a;
    rd_cycle[ 7007] = 1'b0;  wr_cycle[ 7007] = 1'b1;  addr_rom[ 7007]='h00003cc0;  wr_data_rom[ 7007]='h00000f12;
    rd_cycle[ 7008] = 1'b1;  wr_cycle[ 7008] = 1'b0;  addr_rom[ 7008]='h00003cbc;  wr_data_rom[ 7008]='h00000000;
    rd_cycle[ 7009] = 1'b1;  wr_cycle[ 7009] = 1'b0;  addr_rom[ 7009]='h000006f4;  wr_data_rom[ 7009]='h00000000;
    rd_cycle[ 7010] = 1'b1;  wr_cycle[ 7010] = 1'b0;  addr_rom[ 7010]='h00001d70;  wr_data_rom[ 7010]='h00000000;
    rd_cycle[ 7011] = 1'b0;  wr_cycle[ 7011] = 1'b1;  addr_rom[ 7011]='h00003684;  wr_data_rom[ 7011]='h000033af;
    rd_cycle[ 7012] = 1'b0;  wr_cycle[ 7012] = 1'b1;  addr_rom[ 7012]='h000022bc;  wr_data_rom[ 7012]='h00003d4a;
    rd_cycle[ 7013] = 1'b0;  wr_cycle[ 7013] = 1'b1;  addr_rom[ 7013]='h00001168;  wr_data_rom[ 7013]='h00000ecc;
    rd_cycle[ 7014] = 1'b1;  wr_cycle[ 7014] = 1'b0;  addr_rom[ 7014]='h000000d4;  wr_data_rom[ 7014]='h00000000;
    rd_cycle[ 7015] = 1'b1;  wr_cycle[ 7015] = 1'b0;  addr_rom[ 7015]='h000039bc;  wr_data_rom[ 7015]='h00000000;
    rd_cycle[ 7016] = 1'b1;  wr_cycle[ 7016] = 1'b0;  addr_rom[ 7016]='h00002c48;  wr_data_rom[ 7016]='h00000000;
    rd_cycle[ 7017] = 1'b0;  wr_cycle[ 7017] = 1'b1;  addr_rom[ 7017]='h00003e8c;  wr_data_rom[ 7017]='h00000874;
    rd_cycle[ 7018] = 1'b0;  wr_cycle[ 7018] = 1'b1;  addr_rom[ 7018]='h0000042c;  wr_data_rom[ 7018]='h0000138b;
    rd_cycle[ 7019] = 1'b0;  wr_cycle[ 7019] = 1'b1;  addr_rom[ 7019]='h00002e40;  wr_data_rom[ 7019]='h00003dd2;
    rd_cycle[ 7020] = 1'b0;  wr_cycle[ 7020] = 1'b1;  addr_rom[ 7020]='h0000337c;  wr_data_rom[ 7020]='h000019bd;
    rd_cycle[ 7021] = 1'b1;  wr_cycle[ 7021] = 1'b0;  addr_rom[ 7021]='h00000e3c;  wr_data_rom[ 7021]='h00000000;
    rd_cycle[ 7022] = 1'b1;  wr_cycle[ 7022] = 1'b0;  addr_rom[ 7022]='h00000a10;  wr_data_rom[ 7022]='h00000000;
    rd_cycle[ 7023] = 1'b0;  wr_cycle[ 7023] = 1'b1;  addr_rom[ 7023]='h00003178;  wr_data_rom[ 7023]='h00001997;
    rd_cycle[ 7024] = 1'b1;  wr_cycle[ 7024] = 1'b0;  addr_rom[ 7024]='h000012dc;  wr_data_rom[ 7024]='h00000000;
    rd_cycle[ 7025] = 1'b1;  wr_cycle[ 7025] = 1'b0;  addr_rom[ 7025]='h00003200;  wr_data_rom[ 7025]='h00000000;
    rd_cycle[ 7026] = 1'b0;  wr_cycle[ 7026] = 1'b1;  addr_rom[ 7026]='h00000af4;  wr_data_rom[ 7026]='h0000302d;
    rd_cycle[ 7027] = 1'b1;  wr_cycle[ 7027] = 1'b0;  addr_rom[ 7027]='h00002ac8;  wr_data_rom[ 7027]='h00000000;
    rd_cycle[ 7028] = 1'b1;  wr_cycle[ 7028] = 1'b0;  addr_rom[ 7028]='h00000bac;  wr_data_rom[ 7028]='h00000000;
    rd_cycle[ 7029] = 1'b0;  wr_cycle[ 7029] = 1'b1;  addr_rom[ 7029]='h000019a0;  wr_data_rom[ 7029]='h00002e79;
    rd_cycle[ 7030] = 1'b0;  wr_cycle[ 7030] = 1'b1;  addr_rom[ 7030]='h000011b4;  wr_data_rom[ 7030]='h000036e9;
    rd_cycle[ 7031] = 1'b0;  wr_cycle[ 7031] = 1'b1;  addr_rom[ 7031]='h000033f0;  wr_data_rom[ 7031]='h00001834;
    rd_cycle[ 7032] = 1'b1;  wr_cycle[ 7032] = 1'b0;  addr_rom[ 7032]='h00001684;  wr_data_rom[ 7032]='h00000000;
    rd_cycle[ 7033] = 1'b1;  wr_cycle[ 7033] = 1'b0;  addr_rom[ 7033]='h00003b64;  wr_data_rom[ 7033]='h00000000;
    rd_cycle[ 7034] = 1'b1;  wr_cycle[ 7034] = 1'b0;  addr_rom[ 7034]='h00003afc;  wr_data_rom[ 7034]='h00000000;
    rd_cycle[ 7035] = 1'b1;  wr_cycle[ 7035] = 1'b0;  addr_rom[ 7035]='h00000bec;  wr_data_rom[ 7035]='h00000000;
    rd_cycle[ 7036] = 1'b0;  wr_cycle[ 7036] = 1'b1;  addr_rom[ 7036]='h00003670;  wr_data_rom[ 7036]='h00000adf;
    rd_cycle[ 7037] = 1'b0;  wr_cycle[ 7037] = 1'b1;  addr_rom[ 7037]='h00000980;  wr_data_rom[ 7037]='h0000000d;
    rd_cycle[ 7038] = 1'b1;  wr_cycle[ 7038] = 1'b0;  addr_rom[ 7038]='h00002f80;  wr_data_rom[ 7038]='h00000000;
    rd_cycle[ 7039] = 1'b0;  wr_cycle[ 7039] = 1'b1;  addr_rom[ 7039]='h00001ad8;  wr_data_rom[ 7039]='h00000c43;
    rd_cycle[ 7040] = 1'b1;  wr_cycle[ 7040] = 1'b0;  addr_rom[ 7040]='h00000888;  wr_data_rom[ 7040]='h00000000;
    rd_cycle[ 7041] = 1'b1;  wr_cycle[ 7041] = 1'b0;  addr_rom[ 7041]='h000021a4;  wr_data_rom[ 7041]='h00000000;
    rd_cycle[ 7042] = 1'b1;  wr_cycle[ 7042] = 1'b0;  addr_rom[ 7042]='h00001758;  wr_data_rom[ 7042]='h00000000;
    rd_cycle[ 7043] = 1'b0;  wr_cycle[ 7043] = 1'b1;  addr_rom[ 7043]='h000005c4;  wr_data_rom[ 7043]='h0000259d;
    rd_cycle[ 7044] = 1'b1;  wr_cycle[ 7044] = 1'b0;  addr_rom[ 7044]='h00001608;  wr_data_rom[ 7044]='h00000000;
    rd_cycle[ 7045] = 1'b0;  wr_cycle[ 7045] = 1'b1;  addr_rom[ 7045]='h000030e4;  wr_data_rom[ 7045]='h0000287e;
    rd_cycle[ 7046] = 1'b0;  wr_cycle[ 7046] = 1'b1;  addr_rom[ 7046]='h00003720;  wr_data_rom[ 7046]='h00002079;
    rd_cycle[ 7047] = 1'b1;  wr_cycle[ 7047] = 1'b0;  addr_rom[ 7047]='h00000e00;  wr_data_rom[ 7047]='h00000000;
    rd_cycle[ 7048] = 1'b1;  wr_cycle[ 7048] = 1'b0;  addr_rom[ 7048]='h00001db8;  wr_data_rom[ 7048]='h00000000;
    rd_cycle[ 7049] = 1'b0;  wr_cycle[ 7049] = 1'b1;  addr_rom[ 7049]='h000001ac;  wr_data_rom[ 7049]='h00000ab8;
    rd_cycle[ 7050] = 1'b0;  wr_cycle[ 7050] = 1'b1;  addr_rom[ 7050]='h00001e60;  wr_data_rom[ 7050]='h000034c7;
    rd_cycle[ 7051] = 1'b1;  wr_cycle[ 7051] = 1'b0;  addr_rom[ 7051]='h00003254;  wr_data_rom[ 7051]='h00000000;
    rd_cycle[ 7052] = 1'b0;  wr_cycle[ 7052] = 1'b1;  addr_rom[ 7052]='h00001590;  wr_data_rom[ 7052]='h000000b7;
    rd_cycle[ 7053] = 1'b1;  wr_cycle[ 7053] = 1'b0;  addr_rom[ 7053]='h000009a8;  wr_data_rom[ 7053]='h00000000;
    rd_cycle[ 7054] = 1'b1;  wr_cycle[ 7054] = 1'b0;  addr_rom[ 7054]='h00000b34;  wr_data_rom[ 7054]='h00000000;
    rd_cycle[ 7055] = 1'b1;  wr_cycle[ 7055] = 1'b0;  addr_rom[ 7055]='h0000060c;  wr_data_rom[ 7055]='h00000000;
    rd_cycle[ 7056] = 1'b1;  wr_cycle[ 7056] = 1'b0;  addr_rom[ 7056]='h00000508;  wr_data_rom[ 7056]='h00000000;
    rd_cycle[ 7057] = 1'b0;  wr_cycle[ 7057] = 1'b1;  addr_rom[ 7057]='h00003874;  wr_data_rom[ 7057]='h00000f4e;
    rd_cycle[ 7058] = 1'b0;  wr_cycle[ 7058] = 1'b1;  addr_rom[ 7058]='h00000ae8;  wr_data_rom[ 7058]='h00001690;
    rd_cycle[ 7059] = 1'b1;  wr_cycle[ 7059] = 1'b0;  addr_rom[ 7059]='h000003d0;  wr_data_rom[ 7059]='h00000000;
    rd_cycle[ 7060] = 1'b1;  wr_cycle[ 7060] = 1'b0;  addr_rom[ 7060]='h00002508;  wr_data_rom[ 7060]='h00000000;
    rd_cycle[ 7061] = 1'b1;  wr_cycle[ 7061] = 1'b0;  addr_rom[ 7061]='h00003a34;  wr_data_rom[ 7061]='h00000000;
    rd_cycle[ 7062] = 1'b1;  wr_cycle[ 7062] = 1'b0;  addr_rom[ 7062]='h00003bac;  wr_data_rom[ 7062]='h00000000;
    rd_cycle[ 7063] = 1'b0;  wr_cycle[ 7063] = 1'b1;  addr_rom[ 7063]='h000028fc;  wr_data_rom[ 7063]='h00001da2;
    rd_cycle[ 7064] = 1'b1;  wr_cycle[ 7064] = 1'b0;  addr_rom[ 7064]='h00000ba4;  wr_data_rom[ 7064]='h00000000;
    rd_cycle[ 7065] = 1'b1;  wr_cycle[ 7065] = 1'b0;  addr_rom[ 7065]='h000035bc;  wr_data_rom[ 7065]='h00000000;
    rd_cycle[ 7066] = 1'b1;  wr_cycle[ 7066] = 1'b0;  addr_rom[ 7066]='h00003690;  wr_data_rom[ 7066]='h00000000;
    rd_cycle[ 7067] = 1'b0;  wr_cycle[ 7067] = 1'b1;  addr_rom[ 7067]='h00003368;  wr_data_rom[ 7067]='h000017c8;
    rd_cycle[ 7068] = 1'b0;  wr_cycle[ 7068] = 1'b1;  addr_rom[ 7068]='h00003ba0;  wr_data_rom[ 7068]='h000012b6;
    rd_cycle[ 7069] = 1'b1;  wr_cycle[ 7069] = 1'b0;  addr_rom[ 7069]='h00002634;  wr_data_rom[ 7069]='h00000000;
    rd_cycle[ 7070] = 1'b0;  wr_cycle[ 7070] = 1'b1;  addr_rom[ 7070]='h0000380c;  wr_data_rom[ 7070]='h00000ef3;
    rd_cycle[ 7071] = 1'b1;  wr_cycle[ 7071] = 1'b0;  addr_rom[ 7071]='h000023ac;  wr_data_rom[ 7071]='h00000000;
    rd_cycle[ 7072] = 1'b0;  wr_cycle[ 7072] = 1'b1;  addr_rom[ 7072]='h00003014;  wr_data_rom[ 7072]='h00002ba9;
    rd_cycle[ 7073] = 1'b0;  wr_cycle[ 7073] = 1'b1;  addr_rom[ 7073]='h00003998;  wr_data_rom[ 7073]='h00003d1c;
    rd_cycle[ 7074] = 1'b1;  wr_cycle[ 7074] = 1'b0;  addr_rom[ 7074]='h00001008;  wr_data_rom[ 7074]='h00000000;
    rd_cycle[ 7075] = 1'b1;  wr_cycle[ 7075] = 1'b0;  addr_rom[ 7075]='h0000132c;  wr_data_rom[ 7075]='h00000000;
    rd_cycle[ 7076] = 1'b1;  wr_cycle[ 7076] = 1'b0;  addr_rom[ 7076]='h00001b50;  wr_data_rom[ 7076]='h00000000;
    rd_cycle[ 7077] = 1'b1;  wr_cycle[ 7077] = 1'b0;  addr_rom[ 7077]='h000001a0;  wr_data_rom[ 7077]='h00000000;
    rd_cycle[ 7078] = 1'b0;  wr_cycle[ 7078] = 1'b1;  addr_rom[ 7078]='h00003c0c;  wr_data_rom[ 7078]='h00001d86;
    rd_cycle[ 7079] = 1'b0;  wr_cycle[ 7079] = 1'b1;  addr_rom[ 7079]='h00002f78;  wr_data_rom[ 7079]='h00000dc0;
    rd_cycle[ 7080] = 1'b0;  wr_cycle[ 7080] = 1'b1;  addr_rom[ 7080]='h000004b0;  wr_data_rom[ 7080]='h00001d2e;
    rd_cycle[ 7081] = 1'b0;  wr_cycle[ 7081] = 1'b1;  addr_rom[ 7081]='h00001edc;  wr_data_rom[ 7081]='h00002d6a;
    rd_cycle[ 7082] = 1'b1;  wr_cycle[ 7082] = 1'b0;  addr_rom[ 7082]='h00000cb8;  wr_data_rom[ 7082]='h00000000;
    rd_cycle[ 7083] = 1'b1;  wr_cycle[ 7083] = 1'b0;  addr_rom[ 7083]='h000006cc;  wr_data_rom[ 7083]='h00000000;
    rd_cycle[ 7084] = 1'b1;  wr_cycle[ 7084] = 1'b0;  addr_rom[ 7084]='h00000ea4;  wr_data_rom[ 7084]='h00000000;
    rd_cycle[ 7085] = 1'b1;  wr_cycle[ 7085] = 1'b0;  addr_rom[ 7085]='h000017f8;  wr_data_rom[ 7085]='h00000000;
    rd_cycle[ 7086] = 1'b1;  wr_cycle[ 7086] = 1'b0;  addr_rom[ 7086]='h000024d8;  wr_data_rom[ 7086]='h00000000;
    rd_cycle[ 7087] = 1'b0;  wr_cycle[ 7087] = 1'b1;  addr_rom[ 7087]='h0000345c;  wr_data_rom[ 7087]='h00001199;
    rd_cycle[ 7088] = 1'b0;  wr_cycle[ 7088] = 1'b1;  addr_rom[ 7088]='h000006c4;  wr_data_rom[ 7088]='h00003986;
    rd_cycle[ 7089] = 1'b0;  wr_cycle[ 7089] = 1'b1;  addr_rom[ 7089]='h00001a70;  wr_data_rom[ 7089]='h00002245;
    rd_cycle[ 7090] = 1'b1;  wr_cycle[ 7090] = 1'b0;  addr_rom[ 7090]='h000017c0;  wr_data_rom[ 7090]='h00000000;
    rd_cycle[ 7091] = 1'b1;  wr_cycle[ 7091] = 1'b0;  addr_rom[ 7091]='h0000245c;  wr_data_rom[ 7091]='h00000000;
    rd_cycle[ 7092] = 1'b1;  wr_cycle[ 7092] = 1'b0;  addr_rom[ 7092]='h00003c74;  wr_data_rom[ 7092]='h00000000;
    rd_cycle[ 7093] = 1'b1;  wr_cycle[ 7093] = 1'b0;  addr_rom[ 7093]='h00000234;  wr_data_rom[ 7093]='h00000000;
    rd_cycle[ 7094] = 1'b1;  wr_cycle[ 7094] = 1'b0;  addr_rom[ 7094]='h000018bc;  wr_data_rom[ 7094]='h00000000;
    rd_cycle[ 7095] = 1'b1;  wr_cycle[ 7095] = 1'b0;  addr_rom[ 7095]='h00000b1c;  wr_data_rom[ 7095]='h00000000;
    rd_cycle[ 7096] = 1'b0;  wr_cycle[ 7096] = 1'b1;  addr_rom[ 7096]='h00001d54;  wr_data_rom[ 7096]='h00001f4c;
    rd_cycle[ 7097] = 1'b0;  wr_cycle[ 7097] = 1'b1;  addr_rom[ 7097]='h000013fc;  wr_data_rom[ 7097]='h0000121f;
    rd_cycle[ 7098] = 1'b1;  wr_cycle[ 7098] = 1'b0;  addr_rom[ 7098]='h0000121c;  wr_data_rom[ 7098]='h00000000;
    rd_cycle[ 7099] = 1'b1;  wr_cycle[ 7099] = 1'b0;  addr_rom[ 7099]='h00000714;  wr_data_rom[ 7099]='h00000000;
    rd_cycle[ 7100] = 1'b0;  wr_cycle[ 7100] = 1'b1;  addr_rom[ 7100]='h000034d8;  wr_data_rom[ 7100]='h00000529;
    rd_cycle[ 7101] = 1'b0;  wr_cycle[ 7101] = 1'b1;  addr_rom[ 7101]='h000027bc;  wr_data_rom[ 7101]='h000013d3;
    rd_cycle[ 7102] = 1'b1;  wr_cycle[ 7102] = 1'b0;  addr_rom[ 7102]='h000025b4;  wr_data_rom[ 7102]='h00000000;
    rd_cycle[ 7103] = 1'b0;  wr_cycle[ 7103] = 1'b1;  addr_rom[ 7103]='h000013b0;  wr_data_rom[ 7103]='h00002c47;
    rd_cycle[ 7104] = 1'b1;  wr_cycle[ 7104] = 1'b0;  addr_rom[ 7104]='h0000319c;  wr_data_rom[ 7104]='h00000000;
    rd_cycle[ 7105] = 1'b0;  wr_cycle[ 7105] = 1'b1;  addr_rom[ 7105]='h000033b0;  wr_data_rom[ 7105]='h00003a1b;
    rd_cycle[ 7106] = 1'b0;  wr_cycle[ 7106] = 1'b1;  addr_rom[ 7106]='h00000504;  wr_data_rom[ 7106]='h000024d7;
    rd_cycle[ 7107] = 1'b0;  wr_cycle[ 7107] = 1'b1;  addr_rom[ 7107]='h00000e90;  wr_data_rom[ 7107]='h000028b5;
    rd_cycle[ 7108] = 1'b1;  wr_cycle[ 7108] = 1'b0;  addr_rom[ 7108]='h000016c0;  wr_data_rom[ 7108]='h00000000;
    rd_cycle[ 7109] = 1'b1;  wr_cycle[ 7109] = 1'b0;  addr_rom[ 7109]='h00001434;  wr_data_rom[ 7109]='h00000000;
    rd_cycle[ 7110] = 1'b0;  wr_cycle[ 7110] = 1'b1;  addr_rom[ 7110]='h00003d94;  wr_data_rom[ 7110]='h00003172;
    rd_cycle[ 7111] = 1'b0;  wr_cycle[ 7111] = 1'b1;  addr_rom[ 7111]='h000006bc;  wr_data_rom[ 7111]='h000018b4;
    rd_cycle[ 7112] = 1'b1;  wr_cycle[ 7112] = 1'b0;  addr_rom[ 7112]='h00003e88;  wr_data_rom[ 7112]='h00000000;
    rd_cycle[ 7113] = 1'b1;  wr_cycle[ 7113] = 1'b0;  addr_rom[ 7113]='h000026a8;  wr_data_rom[ 7113]='h00000000;
    rd_cycle[ 7114] = 1'b0;  wr_cycle[ 7114] = 1'b1;  addr_rom[ 7114]='h00002e28;  wr_data_rom[ 7114]='h0000324f;
    rd_cycle[ 7115] = 1'b1;  wr_cycle[ 7115] = 1'b0;  addr_rom[ 7115]='h000010c4;  wr_data_rom[ 7115]='h00000000;
    rd_cycle[ 7116] = 1'b1;  wr_cycle[ 7116] = 1'b0;  addr_rom[ 7116]='h000009d0;  wr_data_rom[ 7116]='h00000000;
    rd_cycle[ 7117] = 1'b1;  wr_cycle[ 7117] = 1'b0;  addr_rom[ 7117]='h00002828;  wr_data_rom[ 7117]='h00000000;
    rd_cycle[ 7118] = 1'b0;  wr_cycle[ 7118] = 1'b1;  addr_rom[ 7118]='h00000d78;  wr_data_rom[ 7118]='h000027e6;
    rd_cycle[ 7119] = 1'b1;  wr_cycle[ 7119] = 1'b0;  addr_rom[ 7119]='h00003e64;  wr_data_rom[ 7119]='h00000000;
    rd_cycle[ 7120] = 1'b1;  wr_cycle[ 7120] = 1'b0;  addr_rom[ 7120]='h000016a4;  wr_data_rom[ 7120]='h00000000;
    rd_cycle[ 7121] = 1'b1;  wr_cycle[ 7121] = 1'b0;  addr_rom[ 7121]='h00001bf8;  wr_data_rom[ 7121]='h00000000;
    rd_cycle[ 7122] = 1'b0;  wr_cycle[ 7122] = 1'b1;  addr_rom[ 7122]='h00003238;  wr_data_rom[ 7122]='h00002875;
    rd_cycle[ 7123] = 1'b1;  wr_cycle[ 7123] = 1'b0;  addr_rom[ 7123]='h00003474;  wr_data_rom[ 7123]='h00000000;
    rd_cycle[ 7124] = 1'b1;  wr_cycle[ 7124] = 1'b0;  addr_rom[ 7124]='h0000010c;  wr_data_rom[ 7124]='h00000000;
    rd_cycle[ 7125] = 1'b0;  wr_cycle[ 7125] = 1'b1;  addr_rom[ 7125]='h0000352c;  wr_data_rom[ 7125]='h00001510;
    rd_cycle[ 7126] = 1'b0;  wr_cycle[ 7126] = 1'b1;  addr_rom[ 7126]='h00002708;  wr_data_rom[ 7126]='h00003394;
    rd_cycle[ 7127] = 1'b1;  wr_cycle[ 7127] = 1'b0;  addr_rom[ 7127]='h0000096c;  wr_data_rom[ 7127]='h00000000;
    rd_cycle[ 7128] = 1'b0;  wr_cycle[ 7128] = 1'b1;  addr_rom[ 7128]='h00000d24;  wr_data_rom[ 7128]='h00001fb4;
    rd_cycle[ 7129] = 1'b1;  wr_cycle[ 7129] = 1'b0;  addr_rom[ 7129]='h00002b08;  wr_data_rom[ 7129]='h00000000;
    rd_cycle[ 7130] = 1'b1;  wr_cycle[ 7130] = 1'b0;  addr_rom[ 7130]='h0000019c;  wr_data_rom[ 7130]='h00000000;
    rd_cycle[ 7131] = 1'b1;  wr_cycle[ 7131] = 1'b0;  addr_rom[ 7131]='h00003514;  wr_data_rom[ 7131]='h00000000;
    rd_cycle[ 7132] = 1'b0;  wr_cycle[ 7132] = 1'b1;  addr_rom[ 7132]='h00003480;  wr_data_rom[ 7132]='h0000278a;
    rd_cycle[ 7133] = 1'b1;  wr_cycle[ 7133] = 1'b0;  addr_rom[ 7133]='h000019a8;  wr_data_rom[ 7133]='h00000000;
    rd_cycle[ 7134] = 1'b1;  wr_cycle[ 7134] = 1'b0;  addr_rom[ 7134]='h000032a4;  wr_data_rom[ 7134]='h00000000;
    rd_cycle[ 7135] = 1'b0;  wr_cycle[ 7135] = 1'b1;  addr_rom[ 7135]='h0000221c;  wr_data_rom[ 7135]='h00000a48;
    rd_cycle[ 7136] = 1'b0;  wr_cycle[ 7136] = 1'b1;  addr_rom[ 7136]='h000039b8;  wr_data_rom[ 7136]='h0000060c;
    rd_cycle[ 7137] = 1'b0;  wr_cycle[ 7137] = 1'b1;  addr_rom[ 7137]='h000025d0;  wr_data_rom[ 7137]='h000001f8;
    rd_cycle[ 7138] = 1'b0;  wr_cycle[ 7138] = 1'b1;  addr_rom[ 7138]='h00002b58;  wr_data_rom[ 7138]='h0000366f;
    rd_cycle[ 7139] = 1'b0;  wr_cycle[ 7139] = 1'b1;  addr_rom[ 7139]='h00001e90;  wr_data_rom[ 7139]='h00001d4d;
    rd_cycle[ 7140] = 1'b0;  wr_cycle[ 7140] = 1'b1;  addr_rom[ 7140]='h000009f0;  wr_data_rom[ 7140]='h00000ce7;
    rd_cycle[ 7141] = 1'b0;  wr_cycle[ 7141] = 1'b1;  addr_rom[ 7141]='h00000d6c;  wr_data_rom[ 7141]='h0000209c;
    rd_cycle[ 7142] = 1'b1;  wr_cycle[ 7142] = 1'b0;  addr_rom[ 7142]='h00002758;  wr_data_rom[ 7142]='h00000000;
    rd_cycle[ 7143] = 1'b0;  wr_cycle[ 7143] = 1'b1;  addr_rom[ 7143]='h00003fa4;  wr_data_rom[ 7143]='h00003798;
    rd_cycle[ 7144] = 1'b0;  wr_cycle[ 7144] = 1'b1;  addr_rom[ 7144]='h00002700;  wr_data_rom[ 7144]='h00001298;
    rd_cycle[ 7145] = 1'b0;  wr_cycle[ 7145] = 1'b1;  addr_rom[ 7145]='h00000a04;  wr_data_rom[ 7145]='h00000807;
    rd_cycle[ 7146] = 1'b1;  wr_cycle[ 7146] = 1'b0;  addr_rom[ 7146]='h00002db0;  wr_data_rom[ 7146]='h00000000;
    rd_cycle[ 7147] = 1'b1;  wr_cycle[ 7147] = 1'b0;  addr_rom[ 7147]='h00000d04;  wr_data_rom[ 7147]='h00000000;
    rd_cycle[ 7148] = 1'b0;  wr_cycle[ 7148] = 1'b1;  addr_rom[ 7148]='h00001ee4;  wr_data_rom[ 7148]='h00002853;
    rd_cycle[ 7149] = 1'b0;  wr_cycle[ 7149] = 1'b1;  addr_rom[ 7149]='h00000f88;  wr_data_rom[ 7149]='h00001f9d;
    rd_cycle[ 7150] = 1'b1;  wr_cycle[ 7150] = 1'b0;  addr_rom[ 7150]='h0000254c;  wr_data_rom[ 7150]='h00000000;
    rd_cycle[ 7151] = 1'b0;  wr_cycle[ 7151] = 1'b1;  addr_rom[ 7151]='h0000099c;  wr_data_rom[ 7151]='h000026c8;
    rd_cycle[ 7152] = 1'b0;  wr_cycle[ 7152] = 1'b1;  addr_rom[ 7152]='h000038c8;  wr_data_rom[ 7152]='h00002961;
    rd_cycle[ 7153] = 1'b1;  wr_cycle[ 7153] = 1'b0;  addr_rom[ 7153]='h00002fe4;  wr_data_rom[ 7153]='h00000000;
    rd_cycle[ 7154] = 1'b0;  wr_cycle[ 7154] = 1'b1;  addr_rom[ 7154]='h00003318;  wr_data_rom[ 7154]='h00002fca;
    rd_cycle[ 7155] = 1'b1;  wr_cycle[ 7155] = 1'b0;  addr_rom[ 7155]='h00003730;  wr_data_rom[ 7155]='h00000000;
    rd_cycle[ 7156] = 1'b1;  wr_cycle[ 7156] = 1'b0;  addr_rom[ 7156]='h00001474;  wr_data_rom[ 7156]='h00000000;
    rd_cycle[ 7157] = 1'b0;  wr_cycle[ 7157] = 1'b1;  addr_rom[ 7157]='h000019e8;  wr_data_rom[ 7157]='h00001eca;
    rd_cycle[ 7158] = 1'b0;  wr_cycle[ 7158] = 1'b1;  addr_rom[ 7158]='h00003120;  wr_data_rom[ 7158]='h00001582;
    rd_cycle[ 7159] = 1'b0;  wr_cycle[ 7159] = 1'b1;  addr_rom[ 7159]='h00003980;  wr_data_rom[ 7159]='h00002b9b;
    rd_cycle[ 7160] = 1'b0;  wr_cycle[ 7160] = 1'b1;  addr_rom[ 7160]='h00002b2c;  wr_data_rom[ 7160]='h0000175a;
    rd_cycle[ 7161] = 1'b1;  wr_cycle[ 7161] = 1'b0;  addr_rom[ 7161]='h00001208;  wr_data_rom[ 7161]='h00000000;
    rd_cycle[ 7162] = 1'b0;  wr_cycle[ 7162] = 1'b1;  addr_rom[ 7162]='h00002a30;  wr_data_rom[ 7162]='h00003d8e;
    rd_cycle[ 7163] = 1'b0;  wr_cycle[ 7163] = 1'b1;  addr_rom[ 7163]='h000019f8;  wr_data_rom[ 7163]='h0000051d;
    rd_cycle[ 7164] = 1'b1;  wr_cycle[ 7164] = 1'b0;  addr_rom[ 7164]='h000030ec;  wr_data_rom[ 7164]='h00000000;
    rd_cycle[ 7165] = 1'b0;  wr_cycle[ 7165] = 1'b1;  addr_rom[ 7165]='h00000c58;  wr_data_rom[ 7165]='h000006eb;
    rd_cycle[ 7166] = 1'b1;  wr_cycle[ 7166] = 1'b0;  addr_rom[ 7166]='h00001aa4;  wr_data_rom[ 7166]='h00000000;
    rd_cycle[ 7167] = 1'b0;  wr_cycle[ 7167] = 1'b1;  addr_rom[ 7167]='h00003394;  wr_data_rom[ 7167]='h00002ae6;
    rd_cycle[ 7168] = 1'b0;  wr_cycle[ 7168] = 1'b1;  addr_rom[ 7168]='h000027b0;  wr_data_rom[ 7168]='h00003f5a;
    rd_cycle[ 7169] = 1'b0;  wr_cycle[ 7169] = 1'b1;  addr_rom[ 7169]='h00003104;  wr_data_rom[ 7169]='h000013f6;
    rd_cycle[ 7170] = 1'b0;  wr_cycle[ 7170] = 1'b1;  addr_rom[ 7170]='h00003058;  wr_data_rom[ 7170]='h000020be;
    rd_cycle[ 7171] = 1'b1;  wr_cycle[ 7171] = 1'b0;  addr_rom[ 7171]='h00003c74;  wr_data_rom[ 7171]='h00000000;
    rd_cycle[ 7172] = 1'b0;  wr_cycle[ 7172] = 1'b1;  addr_rom[ 7172]='h0000046c;  wr_data_rom[ 7172]='h00003c0e;
    rd_cycle[ 7173] = 1'b1;  wr_cycle[ 7173] = 1'b0;  addr_rom[ 7173]='h00003118;  wr_data_rom[ 7173]='h00000000;
    rd_cycle[ 7174] = 1'b0;  wr_cycle[ 7174] = 1'b1;  addr_rom[ 7174]='h00000c5c;  wr_data_rom[ 7174]='h00002b32;
    rd_cycle[ 7175] = 1'b0;  wr_cycle[ 7175] = 1'b1;  addr_rom[ 7175]='h00001890;  wr_data_rom[ 7175]='h00000a6c;
    rd_cycle[ 7176] = 1'b0;  wr_cycle[ 7176] = 1'b1;  addr_rom[ 7176]='h00001e44;  wr_data_rom[ 7176]='h00003157;
    rd_cycle[ 7177] = 1'b0;  wr_cycle[ 7177] = 1'b1;  addr_rom[ 7177]='h00000df0;  wr_data_rom[ 7177]='h0000193b;
    rd_cycle[ 7178] = 1'b1;  wr_cycle[ 7178] = 1'b0;  addr_rom[ 7178]='h000009fc;  wr_data_rom[ 7178]='h00000000;
    rd_cycle[ 7179] = 1'b1;  wr_cycle[ 7179] = 1'b0;  addr_rom[ 7179]='h000018a4;  wr_data_rom[ 7179]='h00000000;
    rd_cycle[ 7180] = 1'b1;  wr_cycle[ 7180] = 1'b0;  addr_rom[ 7180]='h0000113c;  wr_data_rom[ 7180]='h00000000;
    rd_cycle[ 7181] = 1'b1;  wr_cycle[ 7181] = 1'b0;  addr_rom[ 7181]='h00001850;  wr_data_rom[ 7181]='h00000000;
    rd_cycle[ 7182] = 1'b1;  wr_cycle[ 7182] = 1'b0;  addr_rom[ 7182]='h00003abc;  wr_data_rom[ 7182]='h00000000;
    rd_cycle[ 7183] = 1'b1;  wr_cycle[ 7183] = 1'b0;  addr_rom[ 7183]='h00000ab8;  wr_data_rom[ 7183]='h00000000;
    rd_cycle[ 7184] = 1'b1;  wr_cycle[ 7184] = 1'b0;  addr_rom[ 7184]='h000036a0;  wr_data_rom[ 7184]='h00000000;
    rd_cycle[ 7185] = 1'b1;  wr_cycle[ 7185] = 1'b0;  addr_rom[ 7185]='h00000230;  wr_data_rom[ 7185]='h00000000;
    rd_cycle[ 7186] = 1'b1;  wr_cycle[ 7186] = 1'b0;  addr_rom[ 7186]='h0000031c;  wr_data_rom[ 7186]='h00000000;
    rd_cycle[ 7187] = 1'b0;  wr_cycle[ 7187] = 1'b1;  addr_rom[ 7187]='h00000dc4;  wr_data_rom[ 7187]='h00001717;
    rd_cycle[ 7188] = 1'b1;  wr_cycle[ 7188] = 1'b0;  addr_rom[ 7188]='h000010d8;  wr_data_rom[ 7188]='h00000000;
    rd_cycle[ 7189] = 1'b1;  wr_cycle[ 7189] = 1'b0;  addr_rom[ 7189]='h0000345c;  wr_data_rom[ 7189]='h00000000;
    rd_cycle[ 7190] = 1'b0;  wr_cycle[ 7190] = 1'b1;  addr_rom[ 7190]='h000003b4;  wr_data_rom[ 7190]='h000016fb;
    rd_cycle[ 7191] = 1'b1;  wr_cycle[ 7191] = 1'b0;  addr_rom[ 7191]='h00000170;  wr_data_rom[ 7191]='h00000000;
    rd_cycle[ 7192] = 1'b0;  wr_cycle[ 7192] = 1'b1;  addr_rom[ 7192]='h00002650;  wr_data_rom[ 7192]='h00001685;
    rd_cycle[ 7193] = 1'b1;  wr_cycle[ 7193] = 1'b0;  addr_rom[ 7193]='h0000296c;  wr_data_rom[ 7193]='h00000000;
    rd_cycle[ 7194] = 1'b0;  wr_cycle[ 7194] = 1'b1;  addr_rom[ 7194]='h00002680;  wr_data_rom[ 7194]='h00002c49;
    rd_cycle[ 7195] = 1'b0;  wr_cycle[ 7195] = 1'b1;  addr_rom[ 7195]='h00000638;  wr_data_rom[ 7195]='h0000219f;
    rd_cycle[ 7196] = 1'b0;  wr_cycle[ 7196] = 1'b1;  addr_rom[ 7196]='h00003954;  wr_data_rom[ 7196]='h0000057c;
    rd_cycle[ 7197] = 1'b0;  wr_cycle[ 7197] = 1'b1;  addr_rom[ 7197]='h00003208;  wr_data_rom[ 7197]='h00003127;
    rd_cycle[ 7198] = 1'b1;  wr_cycle[ 7198] = 1'b0;  addr_rom[ 7198]='h00003518;  wr_data_rom[ 7198]='h00000000;
    rd_cycle[ 7199] = 1'b1;  wr_cycle[ 7199] = 1'b0;  addr_rom[ 7199]='h000027c4;  wr_data_rom[ 7199]='h00000000;
    rd_cycle[ 7200] = 1'b1;  wr_cycle[ 7200] = 1'b0;  addr_rom[ 7200]='h00001864;  wr_data_rom[ 7200]='h00000000;
    rd_cycle[ 7201] = 1'b0;  wr_cycle[ 7201] = 1'b1;  addr_rom[ 7201]='h00002558;  wr_data_rom[ 7201]='h00003594;
    rd_cycle[ 7202] = 1'b0;  wr_cycle[ 7202] = 1'b1;  addr_rom[ 7202]='h0000060c;  wr_data_rom[ 7202]='h000014bf;
    rd_cycle[ 7203] = 1'b1;  wr_cycle[ 7203] = 1'b0;  addr_rom[ 7203]='h00000230;  wr_data_rom[ 7203]='h00000000;
    rd_cycle[ 7204] = 1'b0;  wr_cycle[ 7204] = 1'b1;  addr_rom[ 7204]='h00003f14;  wr_data_rom[ 7204]='h000015a4;
    rd_cycle[ 7205] = 1'b1;  wr_cycle[ 7205] = 1'b0;  addr_rom[ 7205]='h0000158c;  wr_data_rom[ 7205]='h00000000;
    rd_cycle[ 7206] = 1'b0;  wr_cycle[ 7206] = 1'b1;  addr_rom[ 7206]='h00001200;  wr_data_rom[ 7206]='h00000919;
    rd_cycle[ 7207] = 1'b1;  wr_cycle[ 7207] = 1'b0;  addr_rom[ 7207]='h00001840;  wr_data_rom[ 7207]='h00000000;
    rd_cycle[ 7208] = 1'b0;  wr_cycle[ 7208] = 1'b1;  addr_rom[ 7208]='h000020d8;  wr_data_rom[ 7208]='h000018d4;
    rd_cycle[ 7209] = 1'b0;  wr_cycle[ 7209] = 1'b1;  addr_rom[ 7209]='h00000468;  wr_data_rom[ 7209]='h00003b01;
    rd_cycle[ 7210] = 1'b0;  wr_cycle[ 7210] = 1'b1;  addr_rom[ 7210]='h00002330;  wr_data_rom[ 7210]='h000011d9;
    rd_cycle[ 7211] = 1'b1;  wr_cycle[ 7211] = 1'b0;  addr_rom[ 7211]='h000033a0;  wr_data_rom[ 7211]='h00000000;
    rd_cycle[ 7212] = 1'b0;  wr_cycle[ 7212] = 1'b1;  addr_rom[ 7212]='h00000c94;  wr_data_rom[ 7212]='h00002880;
    rd_cycle[ 7213] = 1'b1;  wr_cycle[ 7213] = 1'b0;  addr_rom[ 7213]='h00002414;  wr_data_rom[ 7213]='h00000000;
    rd_cycle[ 7214] = 1'b1;  wr_cycle[ 7214] = 1'b0;  addr_rom[ 7214]='h000022e8;  wr_data_rom[ 7214]='h00000000;
    rd_cycle[ 7215] = 1'b1;  wr_cycle[ 7215] = 1'b0;  addr_rom[ 7215]='h000010ec;  wr_data_rom[ 7215]='h00000000;
    rd_cycle[ 7216] = 1'b0;  wr_cycle[ 7216] = 1'b1;  addr_rom[ 7216]='h00003778;  wr_data_rom[ 7216]='h0000055d;
    rd_cycle[ 7217] = 1'b0;  wr_cycle[ 7217] = 1'b1;  addr_rom[ 7217]='h00000a08;  wr_data_rom[ 7217]='h000007b9;
    rd_cycle[ 7218] = 1'b0;  wr_cycle[ 7218] = 1'b1;  addr_rom[ 7218]='h00003678;  wr_data_rom[ 7218]='h000029a7;
    rd_cycle[ 7219] = 1'b1;  wr_cycle[ 7219] = 1'b0;  addr_rom[ 7219]='h00000078;  wr_data_rom[ 7219]='h00000000;
    rd_cycle[ 7220] = 1'b0;  wr_cycle[ 7220] = 1'b1;  addr_rom[ 7220]='h00002e60;  wr_data_rom[ 7220]='h00003762;
    rd_cycle[ 7221] = 1'b0;  wr_cycle[ 7221] = 1'b1;  addr_rom[ 7221]='h00003ea4;  wr_data_rom[ 7221]='h00001b0d;
    rd_cycle[ 7222] = 1'b1;  wr_cycle[ 7222] = 1'b0;  addr_rom[ 7222]='h00002074;  wr_data_rom[ 7222]='h00000000;
    rd_cycle[ 7223] = 1'b0;  wr_cycle[ 7223] = 1'b1;  addr_rom[ 7223]='h00003368;  wr_data_rom[ 7223]='h00003292;
    rd_cycle[ 7224] = 1'b0;  wr_cycle[ 7224] = 1'b1;  addr_rom[ 7224]='h0000155c;  wr_data_rom[ 7224]='h00003b39;
    rd_cycle[ 7225] = 1'b0;  wr_cycle[ 7225] = 1'b1;  addr_rom[ 7225]='h00000ec8;  wr_data_rom[ 7225]='h00003413;
    rd_cycle[ 7226] = 1'b0;  wr_cycle[ 7226] = 1'b1;  addr_rom[ 7226]='h00003bc4;  wr_data_rom[ 7226]='h00001aaf;
    rd_cycle[ 7227] = 1'b1;  wr_cycle[ 7227] = 1'b0;  addr_rom[ 7227]='h000033c0;  wr_data_rom[ 7227]='h00000000;
    rd_cycle[ 7228] = 1'b0;  wr_cycle[ 7228] = 1'b1;  addr_rom[ 7228]='h00003250;  wr_data_rom[ 7228]='h00003d8d;
    rd_cycle[ 7229] = 1'b0;  wr_cycle[ 7229] = 1'b1;  addr_rom[ 7229]='h00000bc4;  wr_data_rom[ 7229]='h00001584;
    rd_cycle[ 7230] = 1'b1;  wr_cycle[ 7230] = 1'b0;  addr_rom[ 7230]='h000028e8;  wr_data_rom[ 7230]='h00000000;
    rd_cycle[ 7231] = 1'b0;  wr_cycle[ 7231] = 1'b1;  addr_rom[ 7231]='h000009b4;  wr_data_rom[ 7231]='h00001f03;
    rd_cycle[ 7232] = 1'b0;  wr_cycle[ 7232] = 1'b1;  addr_rom[ 7232]='h00000dc4;  wr_data_rom[ 7232]='h000012b1;
    rd_cycle[ 7233] = 1'b1;  wr_cycle[ 7233] = 1'b0;  addr_rom[ 7233]='h00001350;  wr_data_rom[ 7233]='h00000000;
    rd_cycle[ 7234] = 1'b0;  wr_cycle[ 7234] = 1'b1;  addr_rom[ 7234]='h000005d4;  wr_data_rom[ 7234]='h00002be3;
    rd_cycle[ 7235] = 1'b1;  wr_cycle[ 7235] = 1'b0;  addr_rom[ 7235]='h000020c0;  wr_data_rom[ 7235]='h00000000;
    rd_cycle[ 7236] = 1'b1;  wr_cycle[ 7236] = 1'b0;  addr_rom[ 7236]='h000031ec;  wr_data_rom[ 7236]='h00000000;
    rd_cycle[ 7237] = 1'b1;  wr_cycle[ 7237] = 1'b0;  addr_rom[ 7237]='h00000d4c;  wr_data_rom[ 7237]='h00000000;
    rd_cycle[ 7238] = 1'b1;  wr_cycle[ 7238] = 1'b0;  addr_rom[ 7238]='h00003ea8;  wr_data_rom[ 7238]='h00000000;
    rd_cycle[ 7239] = 1'b0;  wr_cycle[ 7239] = 1'b1;  addr_rom[ 7239]='h00001300;  wr_data_rom[ 7239]='h00000f9a;
    rd_cycle[ 7240] = 1'b1;  wr_cycle[ 7240] = 1'b0;  addr_rom[ 7240]='h00000bbc;  wr_data_rom[ 7240]='h00000000;
    rd_cycle[ 7241] = 1'b1;  wr_cycle[ 7241] = 1'b0;  addr_rom[ 7241]='h000035f4;  wr_data_rom[ 7241]='h00000000;
    rd_cycle[ 7242] = 1'b1;  wr_cycle[ 7242] = 1'b0;  addr_rom[ 7242]='h00001308;  wr_data_rom[ 7242]='h00000000;
    rd_cycle[ 7243] = 1'b0;  wr_cycle[ 7243] = 1'b1;  addr_rom[ 7243]='h000012a8;  wr_data_rom[ 7243]='h0000150a;
    rd_cycle[ 7244] = 1'b1;  wr_cycle[ 7244] = 1'b0;  addr_rom[ 7244]='h00000508;  wr_data_rom[ 7244]='h00000000;
    rd_cycle[ 7245] = 1'b0;  wr_cycle[ 7245] = 1'b1;  addr_rom[ 7245]='h00000884;  wr_data_rom[ 7245]='h00001100;
    rd_cycle[ 7246] = 1'b0;  wr_cycle[ 7246] = 1'b1;  addr_rom[ 7246]='h00001ac8;  wr_data_rom[ 7246]='h00003930;
    rd_cycle[ 7247] = 1'b0;  wr_cycle[ 7247] = 1'b1;  addr_rom[ 7247]='h000027fc;  wr_data_rom[ 7247]='h000007c4;
    rd_cycle[ 7248] = 1'b0;  wr_cycle[ 7248] = 1'b1;  addr_rom[ 7248]='h0000350c;  wr_data_rom[ 7248]='h00003688;
    rd_cycle[ 7249] = 1'b1;  wr_cycle[ 7249] = 1'b0;  addr_rom[ 7249]='h00003618;  wr_data_rom[ 7249]='h00000000;
    rd_cycle[ 7250] = 1'b0;  wr_cycle[ 7250] = 1'b1;  addr_rom[ 7250]='h000026c0;  wr_data_rom[ 7250]='h00000edc;
    rd_cycle[ 7251] = 1'b1;  wr_cycle[ 7251] = 1'b0;  addr_rom[ 7251]='h000021e4;  wr_data_rom[ 7251]='h00000000;
    rd_cycle[ 7252] = 1'b0;  wr_cycle[ 7252] = 1'b1;  addr_rom[ 7252]='h00000788;  wr_data_rom[ 7252]='h00000e1f;
    rd_cycle[ 7253] = 1'b1;  wr_cycle[ 7253] = 1'b0;  addr_rom[ 7253]='h000011d0;  wr_data_rom[ 7253]='h00000000;
    rd_cycle[ 7254] = 1'b0;  wr_cycle[ 7254] = 1'b1;  addr_rom[ 7254]='h00000948;  wr_data_rom[ 7254]='h00001b63;
    rd_cycle[ 7255] = 1'b0;  wr_cycle[ 7255] = 1'b1;  addr_rom[ 7255]='h000030a8;  wr_data_rom[ 7255]='h00001540;
    rd_cycle[ 7256] = 1'b0;  wr_cycle[ 7256] = 1'b1;  addr_rom[ 7256]='h00002e14;  wr_data_rom[ 7256]='h0000070e;
    rd_cycle[ 7257] = 1'b0;  wr_cycle[ 7257] = 1'b1;  addr_rom[ 7257]='h0000290c;  wr_data_rom[ 7257]='h00002111;
    rd_cycle[ 7258] = 1'b1;  wr_cycle[ 7258] = 1'b0;  addr_rom[ 7258]='h00001030;  wr_data_rom[ 7258]='h00000000;
    rd_cycle[ 7259] = 1'b1;  wr_cycle[ 7259] = 1'b0;  addr_rom[ 7259]='h00000870;  wr_data_rom[ 7259]='h00000000;
    rd_cycle[ 7260] = 1'b0;  wr_cycle[ 7260] = 1'b1;  addr_rom[ 7260]='h00000810;  wr_data_rom[ 7260]='h00002da2;
    rd_cycle[ 7261] = 1'b0;  wr_cycle[ 7261] = 1'b1;  addr_rom[ 7261]='h00003d88;  wr_data_rom[ 7261]='h0000244e;
    rd_cycle[ 7262] = 1'b1;  wr_cycle[ 7262] = 1'b0;  addr_rom[ 7262]='h000022bc;  wr_data_rom[ 7262]='h00000000;
    rd_cycle[ 7263] = 1'b0;  wr_cycle[ 7263] = 1'b1;  addr_rom[ 7263]='h00002280;  wr_data_rom[ 7263]='h000019f4;
    rd_cycle[ 7264] = 1'b1;  wr_cycle[ 7264] = 1'b0;  addr_rom[ 7264]='h00000528;  wr_data_rom[ 7264]='h00000000;
    rd_cycle[ 7265] = 1'b0;  wr_cycle[ 7265] = 1'b1;  addr_rom[ 7265]='h00003948;  wr_data_rom[ 7265]='h00003e55;
    rd_cycle[ 7266] = 1'b0;  wr_cycle[ 7266] = 1'b1;  addr_rom[ 7266]='h000005ec;  wr_data_rom[ 7266]='h00001700;
    rd_cycle[ 7267] = 1'b0;  wr_cycle[ 7267] = 1'b1;  addr_rom[ 7267]='h00000678;  wr_data_rom[ 7267]='h00000735;
    rd_cycle[ 7268] = 1'b0;  wr_cycle[ 7268] = 1'b1;  addr_rom[ 7268]='h00002488;  wr_data_rom[ 7268]='h0000216b;
    rd_cycle[ 7269] = 1'b0;  wr_cycle[ 7269] = 1'b1;  addr_rom[ 7269]='h000003b8;  wr_data_rom[ 7269]='h00002b45;
    rd_cycle[ 7270] = 1'b0;  wr_cycle[ 7270] = 1'b1;  addr_rom[ 7270]='h00001b1c;  wr_data_rom[ 7270]='h00003f45;
    rd_cycle[ 7271] = 1'b0;  wr_cycle[ 7271] = 1'b1;  addr_rom[ 7271]='h000034cc;  wr_data_rom[ 7271]='h0000079d;
    rd_cycle[ 7272] = 1'b0;  wr_cycle[ 7272] = 1'b1;  addr_rom[ 7272]='h00003c54;  wr_data_rom[ 7272]='h00000a19;
    rd_cycle[ 7273] = 1'b1;  wr_cycle[ 7273] = 1'b0;  addr_rom[ 7273]='h00000688;  wr_data_rom[ 7273]='h00000000;
    rd_cycle[ 7274] = 1'b1;  wr_cycle[ 7274] = 1'b0;  addr_rom[ 7274]='h00003a40;  wr_data_rom[ 7274]='h00000000;
    rd_cycle[ 7275] = 1'b1;  wr_cycle[ 7275] = 1'b0;  addr_rom[ 7275]='h000033e4;  wr_data_rom[ 7275]='h00000000;
    rd_cycle[ 7276] = 1'b0;  wr_cycle[ 7276] = 1'b1;  addr_rom[ 7276]='h00003ba4;  wr_data_rom[ 7276]='h0000321a;
    rd_cycle[ 7277] = 1'b0;  wr_cycle[ 7277] = 1'b1;  addr_rom[ 7277]='h0000397c;  wr_data_rom[ 7277]='h00001c09;
    rd_cycle[ 7278] = 1'b1;  wr_cycle[ 7278] = 1'b0;  addr_rom[ 7278]='h00000b0c;  wr_data_rom[ 7278]='h00000000;
    rd_cycle[ 7279] = 1'b1;  wr_cycle[ 7279] = 1'b0;  addr_rom[ 7279]='h00001c88;  wr_data_rom[ 7279]='h00000000;
    rd_cycle[ 7280] = 1'b0;  wr_cycle[ 7280] = 1'b1;  addr_rom[ 7280]='h00003424;  wr_data_rom[ 7280]='h00001e13;
    rd_cycle[ 7281] = 1'b0;  wr_cycle[ 7281] = 1'b1;  addr_rom[ 7281]='h00003ca4;  wr_data_rom[ 7281]='h00002426;
    rd_cycle[ 7282] = 1'b0;  wr_cycle[ 7282] = 1'b1;  addr_rom[ 7282]='h00000d48;  wr_data_rom[ 7282]='h00002e24;
    rd_cycle[ 7283] = 1'b1;  wr_cycle[ 7283] = 1'b0;  addr_rom[ 7283]='h00000d10;  wr_data_rom[ 7283]='h00000000;
    rd_cycle[ 7284] = 1'b0;  wr_cycle[ 7284] = 1'b1;  addr_rom[ 7284]='h00000b98;  wr_data_rom[ 7284]='h00000355;
    rd_cycle[ 7285] = 1'b0;  wr_cycle[ 7285] = 1'b1;  addr_rom[ 7285]='h00001d28;  wr_data_rom[ 7285]='h00003a92;
    rd_cycle[ 7286] = 1'b1;  wr_cycle[ 7286] = 1'b0;  addr_rom[ 7286]='h000015f0;  wr_data_rom[ 7286]='h00000000;
    rd_cycle[ 7287] = 1'b1;  wr_cycle[ 7287] = 1'b0;  addr_rom[ 7287]='h000036ec;  wr_data_rom[ 7287]='h00000000;
    rd_cycle[ 7288] = 1'b1;  wr_cycle[ 7288] = 1'b0;  addr_rom[ 7288]='h00003284;  wr_data_rom[ 7288]='h00000000;
    rd_cycle[ 7289] = 1'b1;  wr_cycle[ 7289] = 1'b0;  addr_rom[ 7289]='h00001148;  wr_data_rom[ 7289]='h00000000;
    rd_cycle[ 7290] = 1'b1;  wr_cycle[ 7290] = 1'b0;  addr_rom[ 7290]='h00001ca4;  wr_data_rom[ 7290]='h00000000;
    rd_cycle[ 7291] = 1'b1;  wr_cycle[ 7291] = 1'b0;  addr_rom[ 7291]='h000032e8;  wr_data_rom[ 7291]='h00000000;
    rd_cycle[ 7292] = 1'b0;  wr_cycle[ 7292] = 1'b1;  addr_rom[ 7292]='h000035b0;  wr_data_rom[ 7292]='h0000254b;
    rd_cycle[ 7293] = 1'b0;  wr_cycle[ 7293] = 1'b1;  addr_rom[ 7293]='h00002a3c;  wr_data_rom[ 7293]='h00002928;
    rd_cycle[ 7294] = 1'b0;  wr_cycle[ 7294] = 1'b1;  addr_rom[ 7294]='h0000242c;  wr_data_rom[ 7294]='h00001b6c;
    rd_cycle[ 7295] = 1'b0;  wr_cycle[ 7295] = 1'b1;  addr_rom[ 7295]='h00001b18;  wr_data_rom[ 7295]='h0000196e;
    rd_cycle[ 7296] = 1'b0;  wr_cycle[ 7296] = 1'b1;  addr_rom[ 7296]='h00001f48;  wr_data_rom[ 7296]='h00002208;
    rd_cycle[ 7297] = 1'b0;  wr_cycle[ 7297] = 1'b1;  addr_rom[ 7297]='h00000e78;  wr_data_rom[ 7297]='h00001749;
    rd_cycle[ 7298] = 1'b1;  wr_cycle[ 7298] = 1'b0;  addr_rom[ 7298]='h00000ce4;  wr_data_rom[ 7298]='h00000000;
    rd_cycle[ 7299] = 1'b1;  wr_cycle[ 7299] = 1'b0;  addr_rom[ 7299]='h00003eb8;  wr_data_rom[ 7299]='h00000000;
    rd_cycle[ 7300] = 1'b0;  wr_cycle[ 7300] = 1'b1;  addr_rom[ 7300]='h00001b1c;  wr_data_rom[ 7300]='h00001916;
    rd_cycle[ 7301] = 1'b0;  wr_cycle[ 7301] = 1'b1;  addr_rom[ 7301]='h00001b44;  wr_data_rom[ 7301]='h0000041b;
    rd_cycle[ 7302] = 1'b0;  wr_cycle[ 7302] = 1'b1;  addr_rom[ 7302]='h00000618;  wr_data_rom[ 7302]='h0000216f;
    rd_cycle[ 7303] = 1'b1;  wr_cycle[ 7303] = 1'b0;  addr_rom[ 7303]='h0000382c;  wr_data_rom[ 7303]='h00000000;
    rd_cycle[ 7304] = 1'b1;  wr_cycle[ 7304] = 1'b0;  addr_rom[ 7304]='h000021d8;  wr_data_rom[ 7304]='h00000000;
    rd_cycle[ 7305] = 1'b0;  wr_cycle[ 7305] = 1'b1;  addr_rom[ 7305]='h00000dd4;  wr_data_rom[ 7305]='h00001183;
    rd_cycle[ 7306] = 1'b0;  wr_cycle[ 7306] = 1'b1;  addr_rom[ 7306]='h000020ac;  wr_data_rom[ 7306]='h0000055d;
    rd_cycle[ 7307] = 1'b0;  wr_cycle[ 7307] = 1'b1;  addr_rom[ 7307]='h00002a5c;  wr_data_rom[ 7307]='h00000d33;
    rd_cycle[ 7308] = 1'b1;  wr_cycle[ 7308] = 1'b0;  addr_rom[ 7308]='h000024f0;  wr_data_rom[ 7308]='h00000000;
    rd_cycle[ 7309] = 1'b1;  wr_cycle[ 7309] = 1'b0;  addr_rom[ 7309]='h000027a4;  wr_data_rom[ 7309]='h00000000;
    rd_cycle[ 7310] = 1'b1;  wr_cycle[ 7310] = 1'b0;  addr_rom[ 7310]='h00003cb4;  wr_data_rom[ 7310]='h00000000;
    rd_cycle[ 7311] = 1'b0;  wr_cycle[ 7311] = 1'b1;  addr_rom[ 7311]='h000010a4;  wr_data_rom[ 7311]='h00001f95;
    rd_cycle[ 7312] = 1'b1;  wr_cycle[ 7312] = 1'b0;  addr_rom[ 7312]='h00001dac;  wr_data_rom[ 7312]='h00000000;
    rd_cycle[ 7313] = 1'b0;  wr_cycle[ 7313] = 1'b1;  addr_rom[ 7313]='h000027a0;  wr_data_rom[ 7313]='h000018df;
    rd_cycle[ 7314] = 1'b1;  wr_cycle[ 7314] = 1'b0;  addr_rom[ 7314]='h00000620;  wr_data_rom[ 7314]='h00000000;
    rd_cycle[ 7315] = 1'b0;  wr_cycle[ 7315] = 1'b1;  addr_rom[ 7315]='h00000340;  wr_data_rom[ 7315]='h00003c34;
    rd_cycle[ 7316] = 1'b1;  wr_cycle[ 7316] = 1'b0;  addr_rom[ 7316]='h00002e40;  wr_data_rom[ 7316]='h00000000;
    rd_cycle[ 7317] = 1'b0;  wr_cycle[ 7317] = 1'b1;  addr_rom[ 7317]='h00002424;  wr_data_rom[ 7317]='h000011de;
    rd_cycle[ 7318] = 1'b1;  wr_cycle[ 7318] = 1'b0;  addr_rom[ 7318]='h00002360;  wr_data_rom[ 7318]='h00000000;
    rd_cycle[ 7319] = 1'b1;  wr_cycle[ 7319] = 1'b0;  addr_rom[ 7319]='h00000990;  wr_data_rom[ 7319]='h00000000;
    rd_cycle[ 7320] = 1'b1;  wr_cycle[ 7320] = 1'b0;  addr_rom[ 7320]='h00000554;  wr_data_rom[ 7320]='h00000000;
    rd_cycle[ 7321] = 1'b1;  wr_cycle[ 7321] = 1'b0;  addr_rom[ 7321]='h00002e20;  wr_data_rom[ 7321]='h00000000;
    rd_cycle[ 7322] = 1'b0;  wr_cycle[ 7322] = 1'b1;  addr_rom[ 7322]='h00003374;  wr_data_rom[ 7322]='h00001a21;
    rd_cycle[ 7323] = 1'b0;  wr_cycle[ 7323] = 1'b1;  addr_rom[ 7323]='h00003e20;  wr_data_rom[ 7323]='h00002784;
    rd_cycle[ 7324] = 1'b0;  wr_cycle[ 7324] = 1'b1;  addr_rom[ 7324]='h000030c8;  wr_data_rom[ 7324]='h00001524;
    rd_cycle[ 7325] = 1'b0;  wr_cycle[ 7325] = 1'b1;  addr_rom[ 7325]='h000010ec;  wr_data_rom[ 7325]='h00001f91;
    rd_cycle[ 7326] = 1'b0;  wr_cycle[ 7326] = 1'b1;  addr_rom[ 7326]='h00000894;  wr_data_rom[ 7326]='h000001bf;
    rd_cycle[ 7327] = 1'b1;  wr_cycle[ 7327] = 1'b0;  addr_rom[ 7327]='h000022ac;  wr_data_rom[ 7327]='h00000000;
    rd_cycle[ 7328] = 1'b0;  wr_cycle[ 7328] = 1'b1;  addr_rom[ 7328]='h00001fa4;  wr_data_rom[ 7328]='h00000595;
    rd_cycle[ 7329] = 1'b1;  wr_cycle[ 7329] = 1'b0;  addr_rom[ 7329]='h0000232c;  wr_data_rom[ 7329]='h00000000;
    rd_cycle[ 7330] = 1'b1;  wr_cycle[ 7330] = 1'b0;  addr_rom[ 7330]='h000021a4;  wr_data_rom[ 7330]='h00000000;
    rd_cycle[ 7331] = 1'b0;  wr_cycle[ 7331] = 1'b1;  addr_rom[ 7331]='h00003d80;  wr_data_rom[ 7331]='h00000f7e;
    rd_cycle[ 7332] = 1'b0;  wr_cycle[ 7332] = 1'b1;  addr_rom[ 7332]='h00000ee8;  wr_data_rom[ 7332]='h00003118;
    rd_cycle[ 7333] = 1'b0;  wr_cycle[ 7333] = 1'b1;  addr_rom[ 7333]='h00000068;  wr_data_rom[ 7333]='h00002f6d;
    rd_cycle[ 7334] = 1'b1;  wr_cycle[ 7334] = 1'b0;  addr_rom[ 7334]='h00001918;  wr_data_rom[ 7334]='h00000000;
    rd_cycle[ 7335] = 1'b0;  wr_cycle[ 7335] = 1'b1;  addr_rom[ 7335]='h00001fd0;  wr_data_rom[ 7335]='h00000361;
    rd_cycle[ 7336] = 1'b1;  wr_cycle[ 7336] = 1'b0;  addr_rom[ 7336]='h000003e4;  wr_data_rom[ 7336]='h00000000;
    rd_cycle[ 7337] = 1'b1;  wr_cycle[ 7337] = 1'b0;  addr_rom[ 7337]='h00001cec;  wr_data_rom[ 7337]='h00000000;
    rd_cycle[ 7338] = 1'b0;  wr_cycle[ 7338] = 1'b1;  addr_rom[ 7338]='h00000b24;  wr_data_rom[ 7338]='h00003f34;
    rd_cycle[ 7339] = 1'b1;  wr_cycle[ 7339] = 1'b0;  addr_rom[ 7339]='h00001bb4;  wr_data_rom[ 7339]='h00000000;
    rd_cycle[ 7340] = 1'b1;  wr_cycle[ 7340] = 1'b0;  addr_rom[ 7340]='h00001f10;  wr_data_rom[ 7340]='h00000000;
    rd_cycle[ 7341] = 1'b0;  wr_cycle[ 7341] = 1'b1;  addr_rom[ 7341]='h00003e88;  wr_data_rom[ 7341]='h000016c5;
    rd_cycle[ 7342] = 1'b1;  wr_cycle[ 7342] = 1'b0;  addr_rom[ 7342]='h00001164;  wr_data_rom[ 7342]='h00000000;
    rd_cycle[ 7343] = 1'b1;  wr_cycle[ 7343] = 1'b0;  addr_rom[ 7343]='h000009e4;  wr_data_rom[ 7343]='h00000000;
    rd_cycle[ 7344] = 1'b1;  wr_cycle[ 7344] = 1'b0;  addr_rom[ 7344]='h00003b34;  wr_data_rom[ 7344]='h00000000;
    rd_cycle[ 7345] = 1'b0;  wr_cycle[ 7345] = 1'b1;  addr_rom[ 7345]='h000009d0;  wr_data_rom[ 7345]='h00002f71;
    rd_cycle[ 7346] = 1'b0;  wr_cycle[ 7346] = 1'b1;  addr_rom[ 7346]='h00000550;  wr_data_rom[ 7346]='h00003fc5;
    rd_cycle[ 7347] = 1'b0;  wr_cycle[ 7347] = 1'b1;  addr_rom[ 7347]='h0000104c;  wr_data_rom[ 7347]='h00002361;
    rd_cycle[ 7348] = 1'b1;  wr_cycle[ 7348] = 1'b0;  addr_rom[ 7348]='h00001fdc;  wr_data_rom[ 7348]='h00000000;
    rd_cycle[ 7349] = 1'b1;  wr_cycle[ 7349] = 1'b0;  addr_rom[ 7349]='h00002430;  wr_data_rom[ 7349]='h00000000;
    rd_cycle[ 7350] = 1'b1;  wr_cycle[ 7350] = 1'b0;  addr_rom[ 7350]='h0000278c;  wr_data_rom[ 7350]='h00000000;
    rd_cycle[ 7351] = 1'b1;  wr_cycle[ 7351] = 1'b0;  addr_rom[ 7351]='h00003f50;  wr_data_rom[ 7351]='h00000000;
    rd_cycle[ 7352] = 1'b1;  wr_cycle[ 7352] = 1'b0;  addr_rom[ 7352]='h00000668;  wr_data_rom[ 7352]='h00000000;
    rd_cycle[ 7353] = 1'b0;  wr_cycle[ 7353] = 1'b1;  addr_rom[ 7353]='h000003ec;  wr_data_rom[ 7353]='h00001025;
    rd_cycle[ 7354] = 1'b0;  wr_cycle[ 7354] = 1'b1;  addr_rom[ 7354]='h000030a0;  wr_data_rom[ 7354]='h00000b86;
    rd_cycle[ 7355] = 1'b0;  wr_cycle[ 7355] = 1'b1;  addr_rom[ 7355]='h00001714;  wr_data_rom[ 7355]='h000025d3;
    rd_cycle[ 7356] = 1'b0;  wr_cycle[ 7356] = 1'b1;  addr_rom[ 7356]='h00000898;  wr_data_rom[ 7356]='h00000b7b;
    rd_cycle[ 7357] = 1'b0;  wr_cycle[ 7357] = 1'b1;  addr_rom[ 7357]='h00001ac4;  wr_data_rom[ 7357]='h00001ad4;
    rd_cycle[ 7358] = 1'b1;  wr_cycle[ 7358] = 1'b0;  addr_rom[ 7358]='h000005e8;  wr_data_rom[ 7358]='h00000000;
    rd_cycle[ 7359] = 1'b0;  wr_cycle[ 7359] = 1'b1;  addr_rom[ 7359]='h00000548;  wr_data_rom[ 7359]='h00002366;
    rd_cycle[ 7360] = 1'b1;  wr_cycle[ 7360] = 1'b0;  addr_rom[ 7360]='h00001ea0;  wr_data_rom[ 7360]='h00000000;
    rd_cycle[ 7361] = 1'b0;  wr_cycle[ 7361] = 1'b1;  addr_rom[ 7361]='h00002758;  wr_data_rom[ 7361]='h00001017;
    rd_cycle[ 7362] = 1'b0;  wr_cycle[ 7362] = 1'b1;  addr_rom[ 7362]='h0000088c;  wr_data_rom[ 7362]='h00000d30;
    rd_cycle[ 7363] = 1'b1;  wr_cycle[ 7363] = 1'b0;  addr_rom[ 7363]='h00001a64;  wr_data_rom[ 7363]='h00000000;
    rd_cycle[ 7364] = 1'b1;  wr_cycle[ 7364] = 1'b0;  addr_rom[ 7364]='h00002c28;  wr_data_rom[ 7364]='h00000000;
    rd_cycle[ 7365] = 1'b1;  wr_cycle[ 7365] = 1'b0;  addr_rom[ 7365]='h0000336c;  wr_data_rom[ 7365]='h00000000;
    rd_cycle[ 7366] = 1'b0;  wr_cycle[ 7366] = 1'b1;  addr_rom[ 7366]='h00003718;  wr_data_rom[ 7366]='h00001132;
    rd_cycle[ 7367] = 1'b0;  wr_cycle[ 7367] = 1'b1;  addr_rom[ 7367]='h00000fd0;  wr_data_rom[ 7367]='h00001b3f;
    rd_cycle[ 7368] = 1'b1;  wr_cycle[ 7368] = 1'b0;  addr_rom[ 7368]='h00002c6c;  wr_data_rom[ 7368]='h00000000;
    rd_cycle[ 7369] = 1'b0;  wr_cycle[ 7369] = 1'b1;  addr_rom[ 7369]='h000022e0;  wr_data_rom[ 7369]='h00002cb0;
    rd_cycle[ 7370] = 1'b1;  wr_cycle[ 7370] = 1'b0;  addr_rom[ 7370]='h00001b78;  wr_data_rom[ 7370]='h00000000;
    rd_cycle[ 7371] = 1'b0;  wr_cycle[ 7371] = 1'b1;  addr_rom[ 7371]='h00003338;  wr_data_rom[ 7371]='h000013aa;
    rd_cycle[ 7372] = 1'b0;  wr_cycle[ 7372] = 1'b1;  addr_rom[ 7372]='h000004ac;  wr_data_rom[ 7372]='h000016f8;
    rd_cycle[ 7373] = 1'b1;  wr_cycle[ 7373] = 1'b0;  addr_rom[ 7373]='h000018a4;  wr_data_rom[ 7373]='h00000000;
    rd_cycle[ 7374] = 1'b0;  wr_cycle[ 7374] = 1'b1;  addr_rom[ 7374]='h00003610;  wr_data_rom[ 7374]='h000024e1;
    rd_cycle[ 7375] = 1'b1;  wr_cycle[ 7375] = 1'b0;  addr_rom[ 7375]='h00002e48;  wr_data_rom[ 7375]='h00000000;
    rd_cycle[ 7376] = 1'b0;  wr_cycle[ 7376] = 1'b1;  addr_rom[ 7376]='h000011a4;  wr_data_rom[ 7376]='h00002e5c;
    rd_cycle[ 7377] = 1'b1;  wr_cycle[ 7377] = 1'b0;  addr_rom[ 7377]='h00003530;  wr_data_rom[ 7377]='h00000000;
    rd_cycle[ 7378] = 1'b1;  wr_cycle[ 7378] = 1'b0;  addr_rom[ 7378]='h00003a7c;  wr_data_rom[ 7378]='h00000000;
    rd_cycle[ 7379] = 1'b1;  wr_cycle[ 7379] = 1'b0;  addr_rom[ 7379]='h000007e0;  wr_data_rom[ 7379]='h00000000;
    rd_cycle[ 7380] = 1'b1;  wr_cycle[ 7380] = 1'b0;  addr_rom[ 7380]='h00001118;  wr_data_rom[ 7380]='h00000000;
    rd_cycle[ 7381] = 1'b0;  wr_cycle[ 7381] = 1'b1;  addr_rom[ 7381]='h00001c68;  wr_data_rom[ 7381]='h00002b44;
    rd_cycle[ 7382] = 1'b0;  wr_cycle[ 7382] = 1'b1;  addr_rom[ 7382]='h00000cec;  wr_data_rom[ 7382]='h000008e7;
    rd_cycle[ 7383] = 1'b1;  wr_cycle[ 7383] = 1'b0;  addr_rom[ 7383]='h000030d0;  wr_data_rom[ 7383]='h00000000;
    rd_cycle[ 7384] = 1'b1;  wr_cycle[ 7384] = 1'b0;  addr_rom[ 7384]='h000030d4;  wr_data_rom[ 7384]='h00000000;
    rd_cycle[ 7385] = 1'b0;  wr_cycle[ 7385] = 1'b1;  addr_rom[ 7385]='h00003be0;  wr_data_rom[ 7385]='h000016b5;
    rd_cycle[ 7386] = 1'b1;  wr_cycle[ 7386] = 1'b0;  addr_rom[ 7386]='h00000094;  wr_data_rom[ 7386]='h00000000;
    rd_cycle[ 7387] = 1'b0;  wr_cycle[ 7387] = 1'b1;  addr_rom[ 7387]='h00003408;  wr_data_rom[ 7387]='h00002a00;
    rd_cycle[ 7388] = 1'b0;  wr_cycle[ 7388] = 1'b1;  addr_rom[ 7388]='h00003590;  wr_data_rom[ 7388]='h00000662;
    rd_cycle[ 7389] = 1'b0;  wr_cycle[ 7389] = 1'b1;  addr_rom[ 7389]='h00003614;  wr_data_rom[ 7389]='h0000033d;
    rd_cycle[ 7390] = 1'b0;  wr_cycle[ 7390] = 1'b1;  addr_rom[ 7390]='h000015f4;  wr_data_rom[ 7390]='h00002078;
    rd_cycle[ 7391] = 1'b1;  wr_cycle[ 7391] = 1'b0;  addr_rom[ 7391]='h00000318;  wr_data_rom[ 7391]='h00000000;
    rd_cycle[ 7392] = 1'b1;  wr_cycle[ 7392] = 1'b0;  addr_rom[ 7392]='h00003cfc;  wr_data_rom[ 7392]='h00000000;
    rd_cycle[ 7393] = 1'b1;  wr_cycle[ 7393] = 1'b0;  addr_rom[ 7393]='h000014bc;  wr_data_rom[ 7393]='h00000000;
    rd_cycle[ 7394] = 1'b0;  wr_cycle[ 7394] = 1'b1;  addr_rom[ 7394]='h0000399c;  wr_data_rom[ 7394]='h00002b03;
    rd_cycle[ 7395] = 1'b0;  wr_cycle[ 7395] = 1'b1;  addr_rom[ 7395]='h000024c8;  wr_data_rom[ 7395]='h00000394;
    rd_cycle[ 7396] = 1'b1;  wr_cycle[ 7396] = 1'b0;  addr_rom[ 7396]='h000037c8;  wr_data_rom[ 7396]='h00000000;
    rd_cycle[ 7397] = 1'b1;  wr_cycle[ 7397] = 1'b0;  addr_rom[ 7397]='h00000890;  wr_data_rom[ 7397]='h00000000;
    rd_cycle[ 7398] = 1'b1;  wr_cycle[ 7398] = 1'b0;  addr_rom[ 7398]='h00003d9c;  wr_data_rom[ 7398]='h00000000;
    rd_cycle[ 7399] = 1'b0;  wr_cycle[ 7399] = 1'b1;  addr_rom[ 7399]='h0000248c;  wr_data_rom[ 7399]='h000022d1;
    rd_cycle[ 7400] = 1'b0;  wr_cycle[ 7400] = 1'b1;  addr_rom[ 7400]='h000032a8;  wr_data_rom[ 7400]='h0000174a;
    rd_cycle[ 7401] = 1'b1;  wr_cycle[ 7401] = 1'b0;  addr_rom[ 7401]='h00001958;  wr_data_rom[ 7401]='h00000000;
    rd_cycle[ 7402] = 1'b1;  wr_cycle[ 7402] = 1'b0;  addr_rom[ 7402]='h00002974;  wr_data_rom[ 7402]='h00000000;
    rd_cycle[ 7403] = 1'b0;  wr_cycle[ 7403] = 1'b1;  addr_rom[ 7403]='h000004a8;  wr_data_rom[ 7403]='h00000063;
    rd_cycle[ 7404] = 1'b0;  wr_cycle[ 7404] = 1'b1;  addr_rom[ 7404]='h00002d30;  wr_data_rom[ 7404]='h00003b1b;
    rd_cycle[ 7405] = 1'b1;  wr_cycle[ 7405] = 1'b0;  addr_rom[ 7405]='h00000eb0;  wr_data_rom[ 7405]='h00000000;
    rd_cycle[ 7406] = 1'b1;  wr_cycle[ 7406] = 1'b0;  addr_rom[ 7406]='h00002a30;  wr_data_rom[ 7406]='h00000000;
    rd_cycle[ 7407] = 1'b1;  wr_cycle[ 7407] = 1'b0;  addr_rom[ 7407]='h00001eb4;  wr_data_rom[ 7407]='h00000000;
    rd_cycle[ 7408] = 1'b1;  wr_cycle[ 7408] = 1'b0;  addr_rom[ 7408]='h00003bec;  wr_data_rom[ 7408]='h00000000;
    rd_cycle[ 7409] = 1'b0;  wr_cycle[ 7409] = 1'b1;  addr_rom[ 7409]='h00001ec8;  wr_data_rom[ 7409]='h00003800;
    rd_cycle[ 7410] = 1'b1;  wr_cycle[ 7410] = 1'b0;  addr_rom[ 7410]='h00002470;  wr_data_rom[ 7410]='h00000000;
    rd_cycle[ 7411] = 1'b0;  wr_cycle[ 7411] = 1'b1;  addr_rom[ 7411]='h00002564;  wr_data_rom[ 7411]='h00002190;
    rd_cycle[ 7412] = 1'b1;  wr_cycle[ 7412] = 1'b0;  addr_rom[ 7412]='h00001804;  wr_data_rom[ 7412]='h00000000;
    rd_cycle[ 7413] = 1'b0;  wr_cycle[ 7413] = 1'b1;  addr_rom[ 7413]='h00003558;  wr_data_rom[ 7413]='h000013d1;
    rd_cycle[ 7414] = 1'b1;  wr_cycle[ 7414] = 1'b0;  addr_rom[ 7414]='h0000050c;  wr_data_rom[ 7414]='h00000000;
    rd_cycle[ 7415] = 1'b0;  wr_cycle[ 7415] = 1'b1;  addr_rom[ 7415]='h00000280;  wr_data_rom[ 7415]='h00002d8f;
    rd_cycle[ 7416] = 1'b1;  wr_cycle[ 7416] = 1'b0;  addr_rom[ 7416]='h00003768;  wr_data_rom[ 7416]='h00000000;
    rd_cycle[ 7417] = 1'b0;  wr_cycle[ 7417] = 1'b1;  addr_rom[ 7417]='h00001f0c;  wr_data_rom[ 7417]='h00003d02;
    rd_cycle[ 7418] = 1'b0;  wr_cycle[ 7418] = 1'b1;  addr_rom[ 7418]='h00001e54;  wr_data_rom[ 7418]='h000026b6;
    rd_cycle[ 7419] = 1'b0;  wr_cycle[ 7419] = 1'b1;  addr_rom[ 7419]='h000020b0;  wr_data_rom[ 7419]='h00002c28;
    rd_cycle[ 7420] = 1'b1;  wr_cycle[ 7420] = 1'b0;  addr_rom[ 7420]='h00003f40;  wr_data_rom[ 7420]='h00000000;
    rd_cycle[ 7421] = 1'b0;  wr_cycle[ 7421] = 1'b1;  addr_rom[ 7421]='h00001494;  wr_data_rom[ 7421]='h0000095f;
    rd_cycle[ 7422] = 1'b0;  wr_cycle[ 7422] = 1'b1;  addr_rom[ 7422]='h00002388;  wr_data_rom[ 7422]='h00001d8d;
    rd_cycle[ 7423] = 1'b1;  wr_cycle[ 7423] = 1'b0;  addr_rom[ 7423]='h00001c04;  wr_data_rom[ 7423]='h00000000;
    rd_cycle[ 7424] = 1'b1;  wr_cycle[ 7424] = 1'b0;  addr_rom[ 7424]='h00002204;  wr_data_rom[ 7424]='h00000000;
    rd_cycle[ 7425] = 1'b0;  wr_cycle[ 7425] = 1'b1;  addr_rom[ 7425]='h00002c0c;  wr_data_rom[ 7425]='h00002b07;
    rd_cycle[ 7426] = 1'b1;  wr_cycle[ 7426] = 1'b0;  addr_rom[ 7426]='h00001220;  wr_data_rom[ 7426]='h00000000;
    rd_cycle[ 7427] = 1'b1;  wr_cycle[ 7427] = 1'b0;  addr_rom[ 7427]='h00002fa8;  wr_data_rom[ 7427]='h00000000;
    rd_cycle[ 7428] = 1'b0;  wr_cycle[ 7428] = 1'b1;  addr_rom[ 7428]='h00000a50;  wr_data_rom[ 7428]='h00003434;
    rd_cycle[ 7429] = 1'b0;  wr_cycle[ 7429] = 1'b1;  addr_rom[ 7429]='h00001e64;  wr_data_rom[ 7429]='h00000453;
    rd_cycle[ 7430] = 1'b0;  wr_cycle[ 7430] = 1'b1;  addr_rom[ 7430]='h0000372c;  wr_data_rom[ 7430]='h0000340c;
    rd_cycle[ 7431] = 1'b0;  wr_cycle[ 7431] = 1'b1;  addr_rom[ 7431]='h00001d60;  wr_data_rom[ 7431]='h00003883;
    rd_cycle[ 7432] = 1'b0;  wr_cycle[ 7432] = 1'b1;  addr_rom[ 7432]='h00003140;  wr_data_rom[ 7432]='h000011ce;
    rd_cycle[ 7433] = 1'b1;  wr_cycle[ 7433] = 1'b0;  addr_rom[ 7433]='h00002064;  wr_data_rom[ 7433]='h00000000;
    rd_cycle[ 7434] = 1'b0;  wr_cycle[ 7434] = 1'b1;  addr_rom[ 7434]='h00001a14;  wr_data_rom[ 7434]='h00003f11;
    rd_cycle[ 7435] = 1'b1;  wr_cycle[ 7435] = 1'b0;  addr_rom[ 7435]='h00003514;  wr_data_rom[ 7435]='h00000000;
    rd_cycle[ 7436] = 1'b0;  wr_cycle[ 7436] = 1'b1;  addr_rom[ 7436]='h00001588;  wr_data_rom[ 7436]='h0000241b;
    rd_cycle[ 7437] = 1'b0;  wr_cycle[ 7437] = 1'b1;  addr_rom[ 7437]='h00001ef8;  wr_data_rom[ 7437]='h00001164;
    rd_cycle[ 7438] = 1'b0;  wr_cycle[ 7438] = 1'b1;  addr_rom[ 7438]='h000030f0;  wr_data_rom[ 7438]='h00002acb;
    rd_cycle[ 7439] = 1'b1;  wr_cycle[ 7439] = 1'b0;  addr_rom[ 7439]='h000024f8;  wr_data_rom[ 7439]='h00000000;
    rd_cycle[ 7440] = 1'b1;  wr_cycle[ 7440] = 1'b0;  addr_rom[ 7440]='h00002728;  wr_data_rom[ 7440]='h00000000;
    rd_cycle[ 7441] = 1'b1;  wr_cycle[ 7441] = 1'b0;  addr_rom[ 7441]='h00003b18;  wr_data_rom[ 7441]='h00000000;
    rd_cycle[ 7442] = 1'b0;  wr_cycle[ 7442] = 1'b1;  addr_rom[ 7442]='h00000500;  wr_data_rom[ 7442]='h000036b5;
    rd_cycle[ 7443] = 1'b0;  wr_cycle[ 7443] = 1'b1;  addr_rom[ 7443]='h00002a58;  wr_data_rom[ 7443]='h000017f6;
    rd_cycle[ 7444] = 1'b1;  wr_cycle[ 7444] = 1'b0;  addr_rom[ 7444]='h00002a98;  wr_data_rom[ 7444]='h00000000;
    rd_cycle[ 7445] = 1'b0;  wr_cycle[ 7445] = 1'b1;  addr_rom[ 7445]='h00000430;  wr_data_rom[ 7445]='h00003fbb;
    rd_cycle[ 7446] = 1'b0;  wr_cycle[ 7446] = 1'b1;  addr_rom[ 7446]='h00000580;  wr_data_rom[ 7446]='h000029b9;
    rd_cycle[ 7447] = 1'b1;  wr_cycle[ 7447] = 1'b0;  addr_rom[ 7447]='h00001c3c;  wr_data_rom[ 7447]='h00000000;
    rd_cycle[ 7448] = 1'b1;  wr_cycle[ 7448] = 1'b0;  addr_rom[ 7448]='h00001d84;  wr_data_rom[ 7448]='h00000000;
    rd_cycle[ 7449] = 1'b0;  wr_cycle[ 7449] = 1'b1;  addr_rom[ 7449]='h00001638;  wr_data_rom[ 7449]='h00002d2e;
    rd_cycle[ 7450] = 1'b0;  wr_cycle[ 7450] = 1'b1;  addr_rom[ 7450]='h0000357c;  wr_data_rom[ 7450]='h00001cb7;
    rd_cycle[ 7451] = 1'b1;  wr_cycle[ 7451] = 1'b0;  addr_rom[ 7451]='h00001038;  wr_data_rom[ 7451]='h00000000;
    rd_cycle[ 7452] = 1'b0;  wr_cycle[ 7452] = 1'b1;  addr_rom[ 7452]='h000038d0;  wr_data_rom[ 7452]='h000015fb;
    rd_cycle[ 7453] = 1'b0;  wr_cycle[ 7453] = 1'b1;  addr_rom[ 7453]='h000002a0;  wr_data_rom[ 7453]='h0000289c;
    rd_cycle[ 7454] = 1'b0;  wr_cycle[ 7454] = 1'b1;  addr_rom[ 7454]='h000022f4;  wr_data_rom[ 7454]='h00001b0b;
    rd_cycle[ 7455] = 1'b0;  wr_cycle[ 7455] = 1'b1;  addr_rom[ 7455]='h00001e34;  wr_data_rom[ 7455]='h00001a4b;
    rd_cycle[ 7456] = 1'b1;  wr_cycle[ 7456] = 1'b0;  addr_rom[ 7456]='h00001238;  wr_data_rom[ 7456]='h00000000;
    rd_cycle[ 7457] = 1'b0;  wr_cycle[ 7457] = 1'b1;  addr_rom[ 7457]='h00003dcc;  wr_data_rom[ 7457]='h00003c1c;
    rd_cycle[ 7458] = 1'b0;  wr_cycle[ 7458] = 1'b1;  addr_rom[ 7458]='h00002b48;  wr_data_rom[ 7458]='h0000085d;
    rd_cycle[ 7459] = 1'b1;  wr_cycle[ 7459] = 1'b0;  addr_rom[ 7459]='h000001a4;  wr_data_rom[ 7459]='h00000000;
    rd_cycle[ 7460] = 1'b0;  wr_cycle[ 7460] = 1'b1;  addr_rom[ 7460]='h00000328;  wr_data_rom[ 7460]='h0000125b;
    rd_cycle[ 7461] = 1'b1;  wr_cycle[ 7461] = 1'b0;  addr_rom[ 7461]='h00000244;  wr_data_rom[ 7461]='h00000000;
    rd_cycle[ 7462] = 1'b1;  wr_cycle[ 7462] = 1'b0;  addr_rom[ 7462]='h00003a78;  wr_data_rom[ 7462]='h00000000;
    rd_cycle[ 7463] = 1'b1;  wr_cycle[ 7463] = 1'b0;  addr_rom[ 7463]='h00001844;  wr_data_rom[ 7463]='h00000000;
    rd_cycle[ 7464] = 1'b1;  wr_cycle[ 7464] = 1'b0;  addr_rom[ 7464]='h00001928;  wr_data_rom[ 7464]='h00000000;
    rd_cycle[ 7465] = 1'b0;  wr_cycle[ 7465] = 1'b1;  addr_rom[ 7465]='h00003a38;  wr_data_rom[ 7465]='h000016dc;
    rd_cycle[ 7466] = 1'b0;  wr_cycle[ 7466] = 1'b1;  addr_rom[ 7466]='h00002458;  wr_data_rom[ 7466]='h000003ca;
    rd_cycle[ 7467] = 1'b1;  wr_cycle[ 7467] = 1'b0;  addr_rom[ 7467]='h00003638;  wr_data_rom[ 7467]='h00000000;
    rd_cycle[ 7468] = 1'b0;  wr_cycle[ 7468] = 1'b1;  addr_rom[ 7468]='h00001884;  wr_data_rom[ 7468]='h00000ec3;
    rd_cycle[ 7469] = 1'b1;  wr_cycle[ 7469] = 1'b0;  addr_rom[ 7469]='h00003234;  wr_data_rom[ 7469]='h00000000;
    rd_cycle[ 7470] = 1'b0;  wr_cycle[ 7470] = 1'b1;  addr_rom[ 7470]='h00003c6c;  wr_data_rom[ 7470]='h00000b8c;
    rd_cycle[ 7471] = 1'b1;  wr_cycle[ 7471] = 1'b0;  addr_rom[ 7471]='h00003bc4;  wr_data_rom[ 7471]='h00000000;
    rd_cycle[ 7472] = 1'b0;  wr_cycle[ 7472] = 1'b1;  addr_rom[ 7472]='h00002284;  wr_data_rom[ 7472]='h00003661;
    rd_cycle[ 7473] = 1'b1;  wr_cycle[ 7473] = 1'b0;  addr_rom[ 7473]='h00001438;  wr_data_rom[ 7473]='h00000000;
    rd_cycle[ 7474] = 1'b0;  wr_cycle[ 7474] = 1'b1;  addr_rom[ 7474]='h00002134;  wr_data_rom[ 7474]='h00000de7;
    rd_cycle[ 7475] = 1'b0;  wr_cycle[ 7475] = 1'b1;  addr_rom[ 7475]='h00001f34;  wr_data_rom[ 7475]='h00002aa0;
    rd_cycle[ 7476] = 1'b1;  wr_cycle[ 7476] = 1'b0;  addr_rom[ 7476]='h00002064;  wr_data_rom[ 7476]='h00000000;
    rd_cycle[ 7477] = 1'b0;  wr_cycle[ 7477] = 1'b1;  addr_rom[ 7477]='h00001d9c;  wr_data_rom[ 7477]='h00002c36;
    rd_cycle[ 7478] = 1'b0;  wr_cycle[ 7478] = 1'b1;  addr_rom[ 7478]='h00003804;  wr_data_rom[ 7478]='h000036e0;
    rd_cycle[ 7479] = 1'b1;  wr_cycle[ 7479] = 1'b0;  addr_rom[ 7479]='h00003008;  wr_data_rom[ 7479]='h00000000;
    rd_cycle[ 7480] = 1'b1;  wr_cycle[ 7480] = 1'b0;  addr_rom[ 7480]='h000010ac;  wr_data_rom[ 7480]='h00000000;
    rd_cycle[ 7481] = 1'b1;  wr_cycle[ 7481] = 1'b0;  addr_rom[ 7481]='h000014bc;  wr_data_rom[ 7481]='h00000000;
    rd_cycle[ 7482] = 1'b0;  wr_cycle[ 7482] = 1'b1;  addr_rom[ 7482]='h00002378;  wr_data_rom[ 7482]='h00000235;
    rd_cycle[ 7483] = 1'b1;  wr_cycle[ 7483] = 1'b0;  addr_rom[ 7483]='h000013ec;  wr_data_rom[ 7483]='h00000000;
    rd_cycle[ 7484] = 1'b1;  wr_cycle[ 7484] = 1'b0;  addr_rom[ 7484]='h00003384;  wr_data_rom[ 7484]='h00000000;
    rd_cycle[ 7485] = 1'b1;  wr_cycle[ 7485] = 1'b0;  addr_rom[ 7485]='h000030f4;  wr_data_rom[ 7485]='h00000000;
    rd_cycle[ 7486] = 1'b0;  wr_cycle[ 7486] = 1'b1;  addr_rom[ 7486]='h000012e8;  wr_data_rom[ 7486]='h000020ea;
    rd_cycle[ 7487] = 1'b1;  wr_cycle[ 7487] = 1'b0;  addr_rom[ 7487]='h00001d68;  wr_data_rom[ 7487]='h00000000;
    rd_cycle[ 7488] = 1'b0;  wr_cycle[ 7488] = 1'b1;  addr_rom[ 7488]='h000010c8;  wr_data_rom[ 7488]='h00001bce;
    rd_cycle[ 7489] = 1'b1;  wr_cycle[ 7489] = 1'b0;  addr_rom[ 7489]='h00000dd0;  wr_data_rom[ 7489]='h00000000;
    rd_cycle[ 7490] = 1'b0;  wr_cycle[ 7490] = 1'b1;  addr_rom[ 7490]='h00001610;  wr_data_rom[ 7490]='h000038aa;
    rd_cycle[ 7491] = 1'b1;  wr_cycle[ 7491] = 1'b0;  addr_rom[ 7491]='h00000a0c;  wr_data_rom[ 7491]='h00000000;
    rd_cycle[ 7492] = 1'b0;  wr_cycle[ 7492] = 1'b1;  addr_rom[ 7492]='h00000a14;  wr_data_rom[ 7492]='h00000f0c;
    rd_cycle[ 7493] = 1'b0;  wr_cycle[ 7493] = 1'b1;  addr_rom[ 7493]='h00000d00;  wr_data_rom[ 7493]='h00002448;
    rd_cycle[ 7494] = 1'b1;  wr_cycle[ 7494] = 1'b0;  addr_rom[ 7494]='h00000408;  wr_data_rom[ 7494]='h00000000;
    rd_cycle[ 7495] = 1'b1;  wr_cycle[ 7495] = 1'b0;  addr_rom[ 7495]='h00003408;  wr_data_rom[ 7495]='h00000000;
    rd_cycle[ 7496] = 1'b1;  wr_cycle[ 7496] = 1'b0;  addr_rom[ 7496]='h00000198;  wr_data_rom[ 7496]='h00000000;
    rd_cycle[ 7497] = 1'b0;  wr_cycle[ 7497] = 1'b1;  addr_rom[ 7497]='h00003660;  wr_data_rom[ 7497]='h00000763;
    rd_cycle[ 7498] = 1'b1;  wr_cycle[ 7498] = 1'b0;  addr_rom[ 7498]='h0000127c;  wr_data_rom[ 7498]='h00000000;
    rd_cycle[ 7499] = 1'b0;  wr_cycle[ 7499] = 1'b1;  addr_rom[ 7499]='h00001294;  wr_data_rom[ 7499]='h00002873;
    rd_cycle[ 7500] = 1'b0;  wr_cycle[ 7500] = 1'b1;  addr_rom[ 7500]='h000019b0;  wr_data_rom[ 7500]='h00002ad6;
    rd_cycle[ 7501] = 1'b0;  wr_cycle[ 7501] = 1'b1;  addr_rom[ 7501]='h000018e8;  wr_data_rom[ 7501]='h00001efc;
    rd_cycle[ 7502] = 1'b0;  wr_cycle[ 7502] = 1'b1;  addr_rom[ 7502]='h000009c8;  wr_data_rom[ 7502]='h00003df1;
    rd_cycle[ 7503] = 1'b1;  wr_cycle[ 7503] = 1'b0;  addr_rom[ 7503]='h00000504;  wr_data_rom[ 7503]='h00000000;
    rd_cycle[ 7504] = 1'b1;  wr_cycle[ 7504] = 1'b0;  addr_rom[ 7504]='h00000180;  wr_data_rom[ 7504]='h00000000;
    rd_cycle[ 7505] = 1'b1;  wr_cycle[ 7505] = 1'b0;  addr_rom[ 7505]='h0000080c;  wr_data_rom[ 7505]='h00000000;
    rd_cycle[ 7506] = 1'b1;  wr_cycle[ 7506] = 1'b0;  addr_rom[ 7506]='h0000126c;  wr_data_rom[ 7506]='h00000000;
    rd_cycle[ 7507] = 1'b1;  wr_cycle[ 7507] = 1'b0;  addr_rom[ 7507]='h000000c4;  wr_data_rom[ 7507]='h00000000;
    rd_cycle[ 7508] = 1'b1;  wr_cycle[ 7508] = 1'b0;  addr_rom[ 7508]='h00003fb8;  wr_data_rom[ 7508]='h00000000;
    rd_cycle[ 7509] = 1'b0;  wr_cycle[ 7509] = 1'b1;  addr_rom[ 7509]='h00002c6c;  wr_data_rom[ 7509]='h000003e8;
    rd_cycle[ 7510] = 1'b0;  wr_cycle[ 7510] = 1'b1;  addr_rom[ 7510]='h00000048;  wr_data_rom[ 7510]='h000029d8;
    rd_cycle[ 7511] = 1'b1;  wr_cycle[ 7511] = 1'b0;  addr_rom[ 7511]='h00001df8;  wr_data_rom[ 7511]='h00000000;
    rd_cycle[ 7512] = 1'b1;  wr_cycle[ 7512] = 1'b0;  addr_rom[ 7512]='h0000122c;  wr_data_rom[ 7512]='h00000000;
    rd_cycle[ 7513] = 1'b1;  wr_cycle[ 7513] = 1'b0;  addr_rom[ 7513]='h00001c7c;  wr_data_rom[ 7513]='h00000000;
    rd_cycle[ 7514] = 1'b1;  wr_cycle[ 7514] = 1'b0;  addr_rom[ 7514]='h0000123c;  wr_data_rom[ 7514]='h00000000;
    rd_cycle[ 7515] = 1'b0;  wr_cycle[ 7515] = 1'b1;  addr_rom[ 7515]='h00003208;  wr_data_rom[ 7515]='h00001c78;
    rd_cycle[ 7516] = 1'b1;  wr_cycle[ 7516] = 1'b0;  addr_rom[ 7516]='h000003b0;  wr_data_rom[ 7516]='h00000000;
    rd_cycle[ 7517] = 1'b0;  wr_cycle[ 7517] = 1'b1;  addr_rom[ 7517]='h00000fb4;  wr_data_rom[ 7517]='h00001134;
    rd_cycle[ 7518] = 1'b0;  wr_cycle[ 7518] = 1'b1;  addr_rom[ 7518]='h00003f1c;  wr_data_rom[ 7518]='h00000c3f;
    rd_cycle[ 7519] = 1'b0;  wr_cycle[ 7519] = 1'b1;  addr_rom[ 7519]='h000009bc;  wr_data_rom[ 7519]='h000024ce;
    rd_cycle[ 7520] = 1'b1;  wr_cycle[ 7520] = 1'b0;  addr_rom[ 7520]='h00003a30;  wr_data_rom[ 7520]='h00000000;
    rd_cycle[ 7521] = 1'b1;  wr_cycle[ 7521] = 1'b0;  addr_rom[ 7521]='h00000c24;  wr_data_rom[ 7521]='h00000000;
    rd_cycle[ 7522] = 1'b0;  wr_cycle[ 7522] = 1'b1;  addr_rom[ 7522]='h000000b4;  wr_data_rom[ 7522]='h00000f5b;
    rd_cycle[ 7523] = 1'b0;  wr_cycle[ 7523] = 1'b1;  addr_rom[ 7523]='h000015e4;  wr_data_rom[ 7523]='h00002a30;
    rd_cycle[ 7524] = 1'b0;  wr_cycle[ 7524] = 1'b1;  addr_rom[ 7524]='h00003424;  wr_data_rom[ 7524]='h000033fa;
    rd_cycle[ 7525] = 1'b0;  wr_cycle[ 7525] = 1'b1;  addr_rom[ 7525]='h00000674;  wr_data_rom[ 7525]='h00003e8f;
    rd_cycle[ 7526] = 1'b1;  wr_cycle[ 7526] = 1'b0;  addr_rom[ 7526]='h00002e40;  wr_data_rom[ 7526]='h00000000;
    rd_cycle[ 7527] = 1'b0;  wr_cycle[ 7527] = 1'b1;  addr_rom[ 7527]='h00003d14;  wr_data_rom[ 7527]='h000010e8;
    rd_cycle[ 7528] = 1'b0;  wr_cycle[ 7528] = 1'b1;  addr_rom[ 7528]='h00000724;  wr_data_rom[ 7528]='h00001d15;
    rd_cycle[ 7529] = 1'b0;  wr_cycle[ 7529] = 1'b1;  addr_rom[ 7529]='h00002910;  wr_data_rom[ 7529]='h000035fa;
    rd_cycle[ 7530] = 1'b1;  wr_cycle[ 7530] = 1'b0;  addr_rom[ 7530]='h00000d90;  wr_data_rom[ 7530]='h00000000;
    rd_cycle[ 7531] = 1'b1;  wr_cycle[ 7531] = 1'b0;  addr_rom[ 7531]='h00000f2c;  wr_data_rom[ 7531]='h00000000;
    rd_cycle[ 7532] = 1'b1;  wr_cycle[ 7532] = 1'b0;  addr_rom[ 7532]='h00002798;  wr_data_rom[ 7532]='h00000000;
    rd_cycle[ 7533] = 1'b0;  wr_cycle[ 7533] = 1'b1;  addr_rom[ 7533]='h00001c2c;  wr_data_rom[ 7533]='h00003f65;
    rd_cycle[ 7534] = 1'b0;  wr_cycle[ 7534] = 1'b1;  addr_rom[ 7534]='h00002ef8;  wr_data_rom[ 7534]='h00000674;
    rd_cycle[ 7535] = 1'b1;  wr_cycle[ 7535] = 1'b0;  addr_rom[ 7535]='h00001c4c;  wr_data_rom[ 7535]='h00000000;
    rd_cycle[ 7536] = 1'b1;  wr_cycle[ 7536] = 1'b0;  addr_rom[ 7536]='h00003034;  wr_data_rom[ 7536]='h00000000;
    rd_cycle[ 7537] = 1'b0;  wr_cycle[ 7537] = 1'b1;  addr_rom[ 7537]='h00002bbc;  wr_data_rom[ 7537]='h00001745;
    rd_cycle[ 7538] = 1'b1;  wr_cycle[ 7538] = 1'b0;  addr_rom[ 7538]='h00002f4c;  wr_data_rom[ 7538]='h00000000;
    rd_cycle[ 7539] = 1'b0;  wr_cycle[ 7539] = 1'b1;  addr_rom[ 7539]='h0000376c;  wr_data_rom[ 7539]='h00000362;
    rd_cycle[ 7540] = 1'b0;  wr_cycle[ 7540] = 1'b1;  addr_rom[ 7540]='h000027b4;  wr_data_rom[ 7540]='h000026ea;
    rd_cycle[ 7541] = 1'b1;  wr_cycle[ 7541] = 1'b0;  addr_rom[ 7541]='h0000178c;  wr_data_rom[ 7541]='h00000000;
    rd_cycle[ 7542] = 1'b0;  wr_cycle[ 7542] = 1'b1;  addr_rom[ 7542]='h00002870;  wr_data_rom[ 7542]='h000026e4;
    rd_cycle[ 7543] = 1'b0;  wr_cycle[ 7543] = 1'b1;  addr_rom[ 7543]='h0000231c;  wr_data_rom[ 7543]='h00002812;
    rd_cycle[ 7544] = 1'b1;  wr_cycle[ 7544] = 1'b0;  addr_rom[ 7544]='h00000958;  wr_data_rom[ 7544]='h00000000;
    rd_cycle[ 7545] = 1'b0;  wr_cycle[ 7545] = 1'b1;  addr_rom[ 7545]='h00001700;  wr_data_rom[ 7545]='h00002ccb;
    rd_cycle[ 7546] = 1'b1;  wr_cycle[ 7546] = 1'b0;  addr_rom[ 7546]='h00002fbc;  wr_data_rom[ 7546]='h00000000;
    rd_cycle[ 7547] = 1'b0;  wr_cycle[ 7547] = 1'b1;  addr_rom[ 7547]='h00002088;  wr_data_rom[ 7547]='h000020f4;
    rd_cycle[ 7548] = 1'b1;  wr_cycle[ 7548] = 1'b0;  addr_rom[ 7548]='h000020c4;  wr_data_rom[ 7548]='h00000000;
    rd_cycle[ 7549] = 1'b1;  wr_cycle[ 7549] = 1'b0;  addr_rom[ 7549]='h000014b8;  wr_data_rom[ 7549]='h00000000;
    rd_cycle[ 7550] = 1'b0;  wr_cycle[ 7550] = 1'b1;  addr_rom[ 7550]='h00001f4c;  wr_data_rom[ 7550]='h000034dc;
    rd_cycle[ 7551] = 1'b0;  wr_cycle[ 7551] = 1'b1;  addr_rom[ 7551]='h00000d30;  wr_data_rom[ 7551]='h0000245b;
    rd_cycle[ 7552] = 1'b0;  wr_cycle[ 7552] = 1'b1;  addr_rom[ 7552]='h00003330;  wr_data_rom[ 7552]='h00000768;
    rd_cycle[ 7553] = 1'b1;  wr_cycle[ 7553] = 1'b0;  addr_rom[ 7553]='h00000030;  wr_data_rom[ 7553]='h00000000;
    rd_cycle[ 7554] = 1'b1;  wr_cycle[ 7554] = 1'b0;  addr_rom[ 7554]='h00000a4c;  wr_data_rom[ 7554]='h00000000;
    rd_cycle[ 7555] = 1'b1;  wr_cycle[ 7555] = 1'b0;  addr_rom[ 7555]='h00001700;  wr_data_rom[ 7555]='h00000000;
    rd_cycle[ 7556] = 1'b0;  wr_cycle[ 7556] = 1'b1;  addr_rom[ 7556]='h00001068;  wr_data_rom[ 7556]='h0000021b;
    rd_cycle[ 7557] = 1'b1;  wr_cycle[ 7557] = 1'b0;  addr_rom[ 7557]='h000008c8;  wr_data_rom[ 7557]='h00000000;
    rd_cycle[ 7558] = 1'b1;  wr_cycle[ 7558] = 1'b0;  addr_rom[ 7558]='h00000b30;  wr_data_rom[ 7558]='h00000000;
    rd_cycle[ 7559] = 1'b1;  wr_cycle[ 7559] = 1'b0;  addr_rom[ 7559]='h000007b0;  wr_data_rom[ 7559]='h00000000;
    rd_cycle[ 7560] = 1'b1;  wr_cycle[ 7560] = 1'b0;  addr_rom[ 7560]='h00002588;  wr_data_rom[ 7560]='h00000000;
    rd_cycle[ 7561] = 1'b0;  wr_cycle[ 7561] = 1'b1;  addr_rom[ 7561]='h000000f4;  wr_data_rom[ 7561]='h00002a27;
    rd_cycle[ 7562] = 1'b1;  wr_cycle[ 7562] = 1'b0;  addr_rom[ 7562]='h0000066c;  wr_data_rom[ 7562]='h00000000;
    rd_cycle[ 7563] = 1'b0;  wr_cycle[ 7563] = 1'b1;  addr_rom[ 7563]='h000001fc;  wr_data_rom[ 7563]='h00003b0e;
    rd_cycle[ 7564] = 1'b1;  wr_cycle[ 7564] = 1'b0;  addr_rom[ 7564]='h000023f8;  wr_data_rom[ 7564]='h00000000;
    rd_cycle[ 7565] = 1'b0;  wr_cycle[ 7565] = 1'b1;  addr_rom[ 7565]='h0000168c;  wr_data_rom[ 7565]='h0000229d;
    rd_cycle[ 7566] = 1'b1;  wr_cycle[ 7566] = 1'b0;  addr_rom[ 7566]='h00003048;  wr_data_rom[ 7566]='h00000000;
    rd_cycle[ 7567] = 1'b1;  wr_cycle[ 7567] = 1'b0;  addr_rom[ 7567]='h00002c14;  wr_data_rom[ 7567]='h00000000;
    rd_cycle[ 7568] = 1'b0;  wr_cycle[ 7568] = 1'b1;  addr_rom[ 7568]='h000039b8;  wr_data_rom[ 7568]='h0000392e;
    rd_cycle[ 7569] = 1'b1;  wr_cycle[ 7569] = 1'b0;  addr_rom[ 7569]='h00001214;  wr_data_rom[ 7569]='h00000000;
    rd_cycle[ 7570] = 1'b0;  wr_cycle[ 7570] = 1'b1;  addr_rom[ 7570]='h00002264;  wr_data_rom[ 7570]='h00000b59;
    rd_cycle[ 7571] = 1'b0;  wr_cycle[ 7571] = 1'b1;  addr_rom[ 7571]='h00000e44;  wr_data_rom[ 7571]='h000004d9;
    rd_cycle[ 7572] = 1'b0;  wr_cycle[ 7572] = 1'b1;  addr_rom[ 7572]='h0000313c;  wr_data_rom[ 7572]='h00001d09;
    rd_cycle[ 7573] = 1'b0;  wr_cycle[ 7573] = 1'b1;  addr_rom[ 7573]='h00001724;  wr_data_rom[ 7573]='h00000b24;
    rd_cycle[ 7574] = 1'b1;  wr_cycle[ 7574] = 1'b0;  addr_rom[ 7574]='h000008b4;  wr_data_rom[ 7574]='h00000000;
    rd_cycle[ 7575] = 1'b0;  wr_cycle[ 7575] = 1'b1;  addr_rom[ 7575]='h000028cc;  wr_data_rom[ 7575]='h000004a5;
    rd_cycle[ 7576] = 1'b0;  wr_cycle[ 7576] = 1'b1;  addr_rom[ 7576]='h00003310;  wr_data_rom[ 7576]='h00001a05;
    rd_cycle[ 7577] = 1'b1;  wr_cycle[ 7577] = 1'b0;  addr_rom[ 7577]='h00002f94;  wr_data_rom[ 7577]='h00000000;
    rd_cycle[ 7578] = 1'b0;  wr_cycle[ 7578] = 1'b1;  addr_rom[ 7578]='h0000392c;  wr_data_rom[ 7578]='h00001064;
    rd_cycle[ 7579] = 1'b0;  wr_cycle[ 7579] = 1'b1;  addr_rom[ 7579]='h00000648;  wr_data_rom[ 7579]='h00001705;
    rd_cycle[ 7580] = 1'b1;  wr_cycle[ 7580] = 1'b0;  addr_rom[ 7580]='h000018e4;  wr_data_rom[ 7580]='h00000000;
    rd_cycle[ 7581] = 1'b0;  wr_cycle[ 7581] = 1'b1;  addr_rom[ 7581]='h000031a4;  wr_data_rom[ 7581]='h00002cae;
    rd_cycle[ 7582] = 1'b0;  wr_cycle[ 7582] = 1'b1;  addr_rom[ 7582]='h00001ee4;  wr_data_rom[ 7582]='h000011f5;
    rd_cycle[ 7583] = 1'b1;  wr_cycle[ 7583] = 1'b0;  addr_rom[ 7583]='h000016ec;  wr_data_rom[ 7583]='h00000000;
    rd_cycle[ 7584] = 1'b1;  wr_cycle[ 7584] = 1'b0;  addr_rom[ 7584]='h0000031c;  wr_data_rom[ 7584]='h00000000;
    rd_cycle[ 7585] = 1'b1;  wr_cycle[ 7585] = 1'b0;  addr_rom[ 7585]='h000008b8;  wr_data_rom[ 7585]='h00000000;
    rd_cycle[ 7586] = 1'b1;  wr_cycle[ 7586] = 1'b0;  addr_rom[ 7586]='h000019bc;  wr_data_rom[ 7586]='h00000000;
    rd_cycle[ 7587] = 1'b0;  wr_cycle[ 7587] = 1'b1;  addr_rom[ 7587]='h00001bd4;  wr_data_rom[ 7587]='h00003495;
    rd_cycle[ 7588] = 1'b1;  wr_cycle[ 7588] = 1'b0;  addr_rom[ 7588]='h000035e4;  wr_data_rom[ 7588]='h00000000;
    rd_cycle[ 7589] = 1'b1;  wr_cycle[ 7589] = 1'b0;  addr_rom[ 7589]='h00000590;  wr_data_rom[ 7589]='h00000000;
    rd_cycle[ 7590] = 1'b0;  wr_cycle[ 7590] = 1'b1;  addr_rom[ 7590]='h00003474;  wr_data_rom[ 7590]='h000031c7;
    rd_cycle[ 7591] = 1'b1;  wr_cycle[ 7591] = 1'b0;  addr_rom[ 7591]='h000022e0;  wr_data_rom[ 7591]='h00000000;
    rd_cycle[ 7592] = 1'b1;  wr_cycle[ 7592] = 1'b0;  addr_rom[ 7592]='h000015e0;  wr_data_rom[ 7592]='h00000000;
    rd_cycle[ 7593] = 1'b0;  wr_cycle[ 7593] = 1'b1;  addr_rom[ 7593]='h00000a04;  wr_data_rom[ 7593]='h00000f01;
    rd_cycle[ 7594] = 1'b1;  wr_cycle[ 7594] = 1'b0;  addr_rom[ 7594]='h0000354c;  wr_data_rom[ 7594]='h00000000;
    rd_cycle[ 7595] = 1'b0;  wr_cycle[ 7595] = 1'b1;  addr_rom[ 7595]='h00001354;  wr_data_rom[ 7595]='h0000316a;
    rd_cycle[ 7596] = 1'b0;  wr_cycle[ 7596] = 1'b1;  addr_rom[ 7596]='h000009b4;  wr_data_rom[ 7596]='h000039a4;
    rd_cycle[ 7597] = 1'b0;  wr_cycle[ 7597] = 1'b1;  addr_rom[ 7597]='h00003ee0;  wr_data_rom[ 7597]='h00000166;
    rd_cycle[ 7598] = 1'b1;  wr_cycle[ 7598] = 1'b0;  addr_rom[ 7598]='h00003468;  wr_data_rom[ 7598]='h00000000;
    rd_cycle[ 7599] = 1'b1;  wr_cycle[ 7599] = 1'b0;  addr_rom[ 7599]='h000010d4;  wr_data_rom[ 7599]='h00000000;
    rd_cycle[ 7600] = 1'b1;  wr_cycle[ 7600] = 1'b0;  addr_rom[ 7600]='h00003d08;  wr_data_rom[ 7600]='h00000000;
    rd_cycle[ 7601] = 1'b1;  wr_cycle[ 7601] = 1'b0;  addr_rom[ 7601]='h00000bfc;  wr_data_rom[ 7601]='h00000000;
    rd_cycle[ 7602] = 1'b0;  wr_cycle[ 7602] = 1'b1;  addr_rom[ 7602]='h00001d28;  wr_data_rom[ 7602]='h0000083f;
    rd_cycle[ 7603] = 1'b0;  wr_cycle[ 7603] = 1'b1;  addr_rom[ 7603]='h000007a0;  wr_data_rom[ 7603]='h000016b6;
    rd_cycle[ 7604] = 1'b1;  wr_cycle[ 7604] = 1'b0;  addr_rom[ 7604]='h00001854;  wr_data_rom[ 7604]='h00000000;
    rd_cycle[ 7605] = 1'b0;  wr_cycle[ 7605] = 1'b1;  addr_rom[ 7605]='h000038e4;  wr_data_rom[ 7605]='h0000247d;
    rd_cycle[ 7606] = 1'b1;  wr_cycle[ 7606] = 1'b0;  addr_rom[ 7606]='h00002c84;  wr_data_rom[ 7606]='h00000000;
    rd_cycle[ 7607] = 1'b1;  wr_cycle[ 7607] = 1'b0;  addr_rom[ 7607]='h00000794;  wr_data_rom[ 7607]='h00000000;
    rd_cycle[ 7608] = 1'b0;  wr_cycle[ 7608] = 1'b1;  addr_rom[ 7608]='h00000740;  wr_data_rom[ 7608]='h00000cf7;
    rd_cycle[ 7609] = 1'b0;  wr_cycle[ 7609] = 1'b1;  addr_rom[ 7609]='h000036bc;  wr_data_rom[ 7609]='h00003044;
    rd_cycle[ 7610] = 1'b0;  wr_cycle[ 7610] = 1'b1;  addr_rom[ 7610]='h000012fc;  wr_data_rom[ 7610]='h00000f28;
    rd_cycle[ 7611] = 1'b0;  wr_cycle[ 7611] = 1'b1;  addr_rom[ 7611]='h00002fa4;  wr_data_rom[ 7611]='h00002177;
    rd_cycle[ 7612] = 1'b1;  wr_cycle[ 7612] = 1'b0;  addr_rom[ 7612]='h00002d74;  wr_data_rom[ 7612]='h00000000;
    rd_cycle[ 7613] = 1'b0;  wr_cycle[ 7613] = 1'b1;  addr_rom[ 7613]='h00000c28;  wr_data_rom[ 7613]='h00000194;
    rd_cycle[ 7614] = 1'b0;  wr_cycle[ 7614] = 1'b1;  addr_rom[ 7614]='h00000f28;  wr_data_rom[ 7614]='h0000135b;
    rd_cycle[ 7615] = 1'b1;  wr_cycle[ 7615] = 1'b0;  addr_rom[ 7615]='h00002d88;  wr_data_rom[ 7615]='h00000000;
    rd_cycle[ 7616] = 1'b0;  wr_cycle[ 7616] = 1'b1;  addr_rom[ 7616]='h00003654;  wr_data_rom[ 7616]='h000031c7;
    rd_cycle[ 7617] = 1'b0;  wr_cycle[ 7617] = 1'b1;  addr_rom[ 7617]='h00001f2c;  wr_data_rom[ 7617]='h00001100;
    rd_cycle[ 7618] = 1'b1;  wr_cycle[ 7618] = 1'b0;  addr_rom[ 7618]='h000012a4;  wr_data_rom[ 7618]='h00000000;
    rd_cycle[ 7619] = 1'b0;  wr_cycle[ 7619] = 1'b1;  addr_rom[ 7619]='h00001e88;  wr_data_rom[ 7619]='h000022fa;
    rd_cycle[ 7620] = 1'b1;  wr_cycle[ 7620] = 1'b0;  addr_rom[ 7620]='h00002888;  wr_data_rom[ 7620]='h00000000;
    rd_cycle[ 7621] = 1'b1;  wr_cycle[ 7621] = 1'b0;  addr_rom[ 7621]='h00003a14;  wr_data_rom[ 7621]='h00000000;
    rd_cycle[ 7622] = 1'b0;  wr_cycle[ 7622] = 1'b1;  addr_rom[ 7622]='h0000344c;  wr_data_rom[ 7622]='h000006d5;
    rd_cycle[ 7623] = 1'b1;  wr_cycle[ 7623] = 1'b0;  addr_rom[ 7623]='h0000359c;  wr_data_rom[ 7623]='h00000000;
    rd_cycle[ 7624] = 1'b0;  wr_cycle[ 7624] = 1'b1;  addr_rom[ 7624]='h00001fcc;  wr_data_rom[ 7624]='h00002a4f;
    rd_cycle[ 7625] = 1'b0;  wr_cycle[ 7625] = 1'b1;  addr_rom[ 7625]='h00003278;  wr_data_rom[ 7625]='h00002a9d;
    rd_cycle[ 7626] = 1'b1;  wr_cycle[ 7626] = 1'b0;  addr_rom[ 7626]='h00001330;  wr_data_rom[ 7626]='h00000000;
    rd_cycle[ 7627] = 1'b0;  wr_cycle[ 7627] = 1'b1;  addr_rom[ 7627]='h00000b30;  wr_data_rom[ 7627]='h00002c6c;
    rd_cycle[ 7628] = 1'b0;  wr_cycle[ 7628] = 1'b1;  addr_rom[ 7628]='h000018c4;  wr_data_rom[ 7628]='h000022a4;
    rd_cycle[ 7629] = 1'b1;  wr_cycle[ 7629] = 1'b0;  addr_rom[ 7629]='h00001f90;  wr_data_rom[ 7629]='h00000000;
    rd_cycle[ 7630] = 1'b1;  wr_cycle[ 7630] = 1'b0;  addr_rom[ 7630]='h000025a8;  wr_data_rom[ 7630]='h00000000;
    rd_cycle[ 7631] = 1'b0;  wr_cycle[ 7631] = 1'b1;  addr_rom[ 7631]='h000033b4;  wr_data_rom[ 7631]='h0000392c;
    rd_cycle[ 7632] = 1'b1;  wr_cycle[ 7632] = 1'b0;  addr_rom[ 7632]='h000025b4;  wr_data_rom[ 7632]='h00000000;
    rd_cycle[ 7633] = 1'b0;  wr_cycle[ 7633] = 1'b1;  addr_rom[ 7633]='h00000588;  wr_data_rom[ 7633]='h00001095;
    rd_cycle[ 7634] = 1'b0;  wr_cycle[ 7634] = 1'b1;  addr_rom[ 7634]='h00002478;  wr_data_rom[ 7634]='h00001b83;
    rd_cycle[ 7635] = 1'b1;  wr_cycle[ 7635] = 1'b0;  addr_rom[ 7635]='h000026b8;  wr_data_rom[ 7635]='h00000000;
    rd_cycle[ 7636] = 1'b1;  wr_cycle[ 7636] = 1'b0;  addr_rom[ 7636]='h00000960;  wr_data_rom[ 7636]='h00000000;
    rd_cycle[ 7637] = 1'b0;  wr_cycle[ 7637] = 1'b1;  addr_rom[ 7637]='h00000898;  wr_data_rom[ 7637]='h000004cb;
    rd_cycle[ 7638] = 1'b0;  wr_cycle[ 7638] = 1'b1;  addr_rom[ 7638]='h000018d8;  wr_data_rom[ 7638]='h00002ddf;
    rd_cycle[ 7639] = 1'b0;  wr_cycle[ 7639] = 1'b1;  addr_rom[ 7639]='h000013e4;  wr_data_rom[ 7639]='h00001823;
    rd_cycle[ 7640] = 1'b0;  wr_cycle[ 7640] = 1'b1;  addr_rom[ 7640]='h00003d50;  wr_data_rom[ 7640]='h000003a4;
    rd_cycle[ 7641] = 1'b0;  wr_cycle[ 7641] = 1'b1;  addr_rom[ 7641]='h000019a4;  wr_data_rom[ 7641]='h00003e4d;
    rd_cycle[ 7642] = 1'b0;  wr_cycle[ 7642] = 1'b1;  addr_rom[ 7642]='h000007cc;  wr_data_rom[ 7642]='h000039b1;
    rd_cycle[ 7643] = 1'b1;  wr_cycle[ 7643] = 1'b0;  addr_rom[ 7643]='h00003760;  wr_data_rom[ 7643]='h00000000;
    rd_cycle[ 7644] = 1'b1;  wr_cycle[ 7644] = 1'b0;  addr_rom[ 7644]='h00002764;  wr_data_rom[ 7644]='h00000000;
    rd_cycle[ 7645] = 1'b1;  wr_cycle[ 7645] = 1'b0;  addr_rom[ 7645]='h00002e2c;  wr_data_rom[ 7645]='h00000000;
    rd_cycle[ 7646] = 1'b1;  wr_cycle[ 7646] = 1'b0;  addr_rom[ 7646]='h00000458;  wr_data_rom[ 7646]='h00000000;
    rd_cycle[ 7647] = 1'b1;  wr_cycle[ 7647] = 1'b0;  addr_rom[ 7647]='h00003c28;  wr_data_rom[ 7647]='h00000000;
    rd_cycle[ 7648] = 1'b1;  wr_cycle[ 7648] = 1'b0;  addr_rom[ 7648]='h00002a34;  wr_data_rom[ 7648]='h00000000;
    rd_cycle[ 7649] = 1'b1;  wr_cycle[ 7649] = 1'b0;  addr_rom[ 7649]='h00002a3c;  wr_data_rom[ 7649]='h00000000;
    rd_cycle[ 7650] = 1'b0;  wr_cycle[ 7650] = 1'b1;  addr_rom[ 7650]='h00002b30;  wr_data_rom[ 7650]='h0000329d;
    rd_cycle[ 7651] = 1'b0;  wr_cycle[ 7651] = 1'b1;  addr_rom[ 7651]='h00003564;  wr_data_rom[ 7651]='h00003af5;
    rd_cycle[ 7652] = 1'b0;  wr_cycle[ 7652] = 1'b1;  addr_rom[ 7652]='h000025f0;  wr_data_rom[ 7652]='h00002710;
    rd_cycle[ 7653] = 1'b1;  wr_cycle[ 7653] = 1'b0;  addr_rom[ 7653]='h00001fe8;  wr_data_rom[ 7653]='h00000000;
    rd_cycle[ 7654] = 1'b1;  wr_cycle[ 7654] = 1'b0;  addr_rom[ 7654]='h00001fe4;  wr_data_rom[ 7654]='h00000000;
    rd_cycle[ 7655] = 1'b1;  wr_cycle[ 7655] = 1'b0;  addr_rom[ 7655]='h000023e4;  wr_data_rom[ 7655]='h00000000;
    rd_cycle[ 7656] = 1'b1;  wr_cycle[ 7656] = 1'b0;  addr_rom[ 7656]='h00002588;  wr_data_rom[ 7656]='h00000000;
    rd_cycle[ 7657] = 1'b1;  wr_cycle[ 7657] = 1'b0;  addr_rom[ 7657]='h000000a0;  wr_data_rom[ 7657]='h00000000;
    rd_cycle[ 7658] = 1'b1;  wr_cycle[ 7658] = 1'b0;  addr_rom[ 7658]='h00000654;  wr_data_rom[ 7658]='h00000000;
    rd_cycle[ 7659] = 1'b0;  wr_cycle[ 7659] = 1'b1;  addr_rom[ 7659]='h00002950;  wr_data_rom[ 7659]='h000005e7;
    rd_cycle[ 7660] = 1'b0;  wr_cycle[ 7660] = 1'b1;  addr_rom[ 7660]='h0000224c;  wr_data_rom[ 7660]='h00002efe;
    rd_cycle[ 7661] = 1'b0;  wr_cycle[ 7661] = 1'b1;  addr_rom[ 7661]='h000029cc;  wr_data_rom[ 7661]='h00001c79;
    rd_cycle[ 7662] = 1'b1;  wr_cycle[ 7662] = 1'b0;  addr_rom[ 7662]='h00000bdc;  wr_data_rom[ 7662]='h00000000;
    rd_cycle[ 7663] = 1'b0;  wr_cycle[ 7663] = 1'b1;  addr_rom[ 7663]='h000006a4;  wr_data_rom[ 7663]='h0000010a;
    rd_cycle[ 7664] = 1'b1;  wr_cycle[ 7664] = 1'b0;  addr_rom[ 7664]='h00002640;  wr_data_rom[ 7664]='h00000000;
    rd_cycle[ 7665] = 1'b1;  wr_cycle[ 7665] = 1'b0;  addr_rom[ 7665]='h00002184;  wr_data_rom[ 7665]='h00000000;
    rd_cycle[ 7666] = 1'b0;  wr_cycle[ 7666] = 1'b1;  addr_rom[ 7666]='h00003e10;  wr_data_rom[ 7666]='h0000272f;
    rd_cycle[ 7667] = 1'b1;  wr_cycle[ 7667] = 1'b0;  addr_rom[ 7667]='h00002594;  wr_data_rom[ 7667]='h00000000;
    rd_cycle[ 7668] = 1'b1;  wr_cycle[ 7668] = 1'b0;  addr_rom[ 7668]='h00000a58;  wr_data_rom[ 7668]='h00000000;
    rd_cycle[ 7669] = 1'b0;  wr_cycle[ 7669] = 1'b1;  addr_rom[ 7669]='h000013cc;  wr_data_rom[ 7669]='h00001261;
    rd_cycle[ 7670] = 1'b1;  wr_cycle[ 7670] = 1'b0;  addr_rom[ 7670]='h00002500;  wr_data_rom[ 7670]='h00000000;
    rd_cycle[ 7671] = 1'b1;  wr_cycle[ 7671] = 1'b0;  addr_rom[ 7671]='h00002800;  wr_data_rom[ 7671]='h00000000;
    rd_cycle[ 7672] = 1'b1;  wr_cycle[ 7672] = 1'b0;  addr_rom[ 7672]='h00000c5c;  wr_data_rom[ 7672]='h00000000;
    rd_cycle[ 7673] = 1'b0;  wr_cycle[ 7673] = 1'b1;  addr_rom[ 7673]='h00000e38;  wr_data_rom[ 7673]='h00001dc7;
    rd_cycle[ 7674] = 1'b1;  wr_cycle[ 7674] = 1'b0;  addr_rom[ 7674]='h00003d8c;  wr_data_rom[ 7674]='h00000000;
    rd_cycle[ 7675] = 1'b0;  wr_cycle[ 7675] = 1'b1;  addr_rom[ 7675]='h00001b84;  wr_data_rom[ 7675]='h000018cb;
    rd_cycle[ 7676] = 1'b0;  wr_cycle[ 7676] = 1'b1;  addr_rom[ 7676]='h0000315c;  wr_data_rom[ 7676]='h00002c62;
    rd_cycle[ 7677] = 1'b0;  wr_cycle[ 7677] = 1'b1;  addr_rom[ 7677]='h0000213c;  wr_data_rom[ 7677]='h00002b67;
    rd_cycle[ 7678] = 1'b1;  wr_cycle[ 7678] = 1'b0;  addr_rom[ 7678]='h0000156c;  wr_data_rom[ 7678]='h00000000;
    rd_cycle[ 7679] = 1'b1;  wr_cycle[ 7679] = 1'b0;  addr_rom[ 7679]='h00003b30;  wr_data_rom[ 7679]='h00000000;
    rd_cycle[ 7680] = 1'b1;  wr_cycle[ 7680] = 1'b0;  addr_rom[ 7680]='h000022c0;  wr_data_rom[ 7680]='h00000000;
    rd_cycle[ 7681] = 1'b0;  wr_cycle[ 7681] = 1'b1;  addr_rom[ 7681]='h00002580;  wr_data_rom[ 7681]='h00002b1d;
    rd_cycle[ 7682] = 1'b1;  wr_cycle[ 7682] = 1'b0;  addr_rom[ 7682]='h0000184c;  wr_data_rom[ 7682]='h00000000;
    rd_cycle[ 7683] = 1'b1;  wr_cycle[ 7683] = 1'b0;  addr_rom[ 7683]='h00000d74;  wr_data_rom[ 7683]='h00000000;
    rd_cycle[ 7684] = 1'b0;  wr_cycle[ 7684] = 1'b1;  addr_rom[ 7684]='h00002e18;  wr_data_rom[ 7684]='h000001a7;
    rd_cycle[ 7685] = 1'b1;  wr_cycle[ 7685] = 1'b0;  addr_rom[ 7685]='h00003dcc;  wr_data_rom[ 7685]='h00000000;
    rd_cycle[ 7686] = 1'b1;  wr_cycle[ 7686] = 1'b0;  addr_rom[ 7686]='h00002008;  wr_data_rom[ 7686]='h00000000;
    rd_cycle[ 7687] = 1'b1;  wr_cycle[ 7687] = 1'b0;  addr_rom[ 7687]='h000006cc;  wr_data_rom[ 7687]='h00000000;
    rd_cycle[ 7688] = 1'b1;  wr_cycle[ 7688] = 1'b0;  addr_rom[ 7688]='h00002f90;  wr_data_rom[ 7688]='h00000000;
    rd_cycle[ 7689] = 1'b1;  wr_cycle[ 7689] = 1'b0;  addr_rom[ 7689]='h00002ed8;  wr_data_rom[ 7689]='h00000000;
    rd_cycle[ 7690] = 1'b0;  wr_cycle[ 7690] = 1'b1;  addr_rom[ 7690]='h0000042c;  wr_data_rom[ 7690]='h00003b3a;
    rd_cycle[ 7691] = 1'b1;  wr_cycle[ 7691] = 1'b0;  addr_rom[ 7691]='h000016b0;  wr_data_rom[ 7691]='h00000000;
    rd_cycle[ 7692] = 1'b1;  wr_cycle[ 7692] = 1'b0;  addr_rom[ 7692]='h00003690;  wr_data_rom[ 7692]='h00000000;
    rd_cycle[ 7693] = 1'b0;  wr_cycle[ 7693] = 1'b1;  addr_rom[ 7693]='h0000234c;  wr_data_rom[ 7693]='h00002569;
    rd_cycle[ 7694] = 1'b1;  wr_cycle[ 7694] = 1'b0;  addr_rom[ 7694]='h00003134;  wr_data_rom[ 7694]='h00000000;
    rd_cycle[ 7695] = 1'b1;  wr_cycle[ 7695] = 1'b0;  addr_rom[ 7695]='h00002004;  wr_data_rom[ 7695]='h00000000;
    rd_cycle[ 7696] = 1'b0;  wr_cycle[ 7696] = 1'b1;  addr_rom[ 7696]='h00001448;  wr_data_rom[ 7696]='h00001a18;
    rd_cycle[ 7697] = 1'b1;  wr_cycle[ 7697] = 1'b0;  addr_rom[ 7697]='h0000130c;  wr_data_rom[ 7697]='h00000000;
    rd_cycle[ 7698] = 1'b0;  wr_cycle[ 7698] = 1'b1;  addr_rom[ 7698]='h0000042c;  wr_data_rom[ 7698]='h00002afb;
    rd_cycle[ 7699] = 1'b1;  wr_cycle[ 7699] = 1'b0;  addr_rom[ 7699]='h000033bc;  wr_data_rom[ 7699]='h00000000;
    rd_cycle[ 7700] = 1'b1;  wr_cycle[ 7700] = 1'b0;  addr_rom[ 7700]='h00000928;  wr_data_rom[ 7700]='h00000000;
    rd_cycle[ 7701] = 1'b0;  wr_cycle[ 7701] = 1'b1;  addr_rom[ 7701]='h0000013c;  wr_data_rom[ 7701]='h00002478;
    rd_cycle[ 7702] = 1'b0;  wr_cycle[ 7702] = 1'b1;  addr_rom[ 7702]='h00001b1c;  wr_data_rom[ 7702]='h000014d5;
    rd_cycle[ 7703] = 1'b1;  wr_cycle[ 7703] = 1'b0;  addr_rom[ 7703]='h00000c3c;  wr_data_rom[ 7703]='h00000000;
    rd_cycle[ 7704] = 1'b1;  wr_cycle[ 7704] = 1'b0;  addr_rom[ 7704]='h00003364;  wr_data_rom[ 7704]='h00000000;
    rd_cycle[ 7705] = 1'b0;  wr_cycle[ 7705] = 1'b1;  addr_rom[ 7705]='h000022ac;  wr_data_rom[ 7705]='h0000106d;
    rd_cycle[ 7706] = 1'b0;  wr_cycle[ 7706] = 1'b1;  addr_rom[ 7706]='h000026f8;  wr_data_rom[ 7706]='h0000049e;
    rd_cycle[ 7707] = 1'b1;  wr_cycle[ 7707] = 1'b0;  addr_rom[ 7707]='h0000373c;  wr_data_rom[ 7707]='h00000000;
    rd_cycle[ 7708] = 1'b1;  wr_cycle[ 7708] = 1'b0;  addr_rom[ 7708]='h00002270;  wr_data_rom[ 7708]='h00000000;
    rd_cycle[ 7709] = 1'b0;  wr_cycle[ 7709] = 1'b1;  addr_rom[ 7709]='h000017f4;  wr_data_rom[ 7709]='h000012d3;
    rd_cycle[ 7710] = 1'b0;  wr_cycle[ 7710] = 1'b1;  addr_rom[ 7710]='h00002a90;  wr_data_rom[ 7710]='h00003a41;
    rd_cycle[ 7711] = 1'b0;  wr_cycle[ 7711] = 1'b1;  addr_rom[ 7711]='h00002534;  wr_data_rom[ 7711]='h000027df;
    rd_cycle[ 7712] = 1'b0;  wr_cycle[ 7712] = 1'b1;  addr_rom[ 7712]='h00001d44;  wr_data_rom[ 7712]='h00000829;
    rd_cycle[ 7713] = 1'b1;  wr_cycle[ 7713] = 1'b0;  addr_rom[ 7713]='h00003848;  wr_data_rom[ 7713]='h00000000;
    rd_cycle[ 7714] = 1'b1;  wr_cycle[ 7714] = 1'b0;  addr_rom[ 7714]='h00002cb4;  wr_data_rom[ 7714]='h00000000;
    rd_cycle[ 7715] = 1'b1;  wr_cycle[ 7715] = 1'b0;  addr_rom[ 7715]='h00001e54;  wr_data_rom[ 7715]='h00000000;
    rd_cycle[ 7716] = 1'b0;  wr_cycle[ 7716] = 1'b1;  addr_rom[ 7716]='h000033bc;  wr_data_rom[ 7716]='h00001d04;
    rd_cycle[ 7717] = 1'b0;  wr_cycle[ 7717] = 1'b1;  addr_rom[ 7717]='h00002f68;  wr_data_rom[ 7717]='h00002d2e;
    rd_cycle[ 7718] = 1'b1;  wr_cycle[ 7718] = 1'b0;  addr_rom[ 7718]='h00002530;  wr_data_rom[ 7718]='h00000000;
    rd_cycle[ 7719] = 1'b0;  wr_cycle[ 7719] = 1'b1;  addr_rom[ 7719]='h00001870;  wr_data_rom[ 7719]='h00003e6c;
    rd_cycle[ 7720] = 1'b0;  wr_cycle[ 7720] = 1'b1;  addr_rom[ 7720]='h000021fc;  wr_data_rom[ 7720]='h000032fb;
    rd_cycle[ 7721] = 1'b1;  wr_cycle[ 7721] = 1'b0;  addr_rom[ 7721]='h00002d24;  wr_data_rom[ 7721]='h00000000;
    rd_cycle[ 7722] = 1'b1;  wr_cycle[ 7722] = 1'b0;  addr_rom[ 7722]='h000029bc;  wr_data_rom[ 7722]='h00000000;
    rd_cycle[ 7723] = 1'b1;  wr_cycle[ 7723] = 1'b0;  addr_rom[ 7723]='h00002878;  wr_data_rom[ 7723]='h00000000;
    rd_cycle[ 7724] = 1'b1;  wr_cycle[ 7724] = 1'b0;  addr_rom[ 7724]='h00000cdc;  wr_data_rom[ 7724]='h00000000;
    rd_cycle[ 7725] = 1'b0;  wr_cycle[ 7725] = 1'b1;  addr_rom[ 7725]='h00001e24;  wr_data_rom[ 7725]='h000013ba;
    rd_cycle[ 7726] = 1'b1;  wr_cycle[ 7726] = 1'b0;  addr_rom[ 7726]='h00001ce4;  wr_data_rom[ 7726]='h00000000;
    rd_cycle[ 7727] = 1'b0;  wr_cycle[ 7727] = 1'b1;  addr_rom[ 7727]='h00001fd0;  wr_data_rom[ 7727]='h00001fd7;
    rd_cycle[ 7728] = 1'b0;  wr_cycle[ 7728] = 1'b1;  addr_rom[ 7728]='h00000c48;  wr_data_rom[ 7728]='h000030e3;
    rd_cycle[ 7729] = 1'b1;  wr_cycle[ 7729] = 1'b0;  addr_rom[ 7729]='h00001ad0;  wr_data_rom[ 7729]='h00000000;
    rd_cycle[ 7730] = 1'b1;  wr_cycle[ 7730] = 1'b0;  addr_rom[ 7730]='h00003820;  wr_data_rom[ 7730]='h00000000;
    rd_cycle[ 7731] = 1'b1;  wr_cycle[ 7731] = 1'b0;  addr_rom[ 7731]='h000001ac;  wr_data_rom[ 7731]='h00000000;
    rd_cycle[ 7732] = 1'b0;  wr_cycle[ 7732] = 1'b1;  addr_rom[ 7732]='h00003f44;  wr_data_rom[ 7732]='h00000f16;
    rd_cycle[ 7733] = 1'b0;  wr_cycle[ 7733] = 1'b1;  addr_rom[ 7733]='h00002ef4;  wr_data_rom[ 7733]='h0000094e;
    rd_cycle[ 7734] = 1'b1;  wr_cycle[ 7734] = 1'b0;  addr_rom[ 7734]='h00000dbc;  wr_data_rom[ 7734]='h00000000;
    rd_cycle[ 7735] = 1'b1;  wr_cycle[ 7735] = 1'b0;  addr_rom[ 7735]='h000012c4;  wr_data_rom[ 7735]='h00000000;
    rd_cycle[ 7736] = 1'b1;  wr_cycle[ 7736] = 1'b0;  addr_rom[ 7736]='h00001d2c;  wr_data_rom[ 7736]='h00000000;
    rd_cycle[ 7737] = 1'b1;  wr_cycle[ 7737] = 1'b0;  addr_rom[ 7737]='h000012dc;  wr_data_rom[ 7737]='h00000000;
    rd_cycle[ 7738] = 1'b0;  wr_cycle[ 7738] = 1'b1;  addr_rom[ 7738]='h00002f34;  wr_data_rom[ 7738]='h00000271;
    rd_cycle[ 7739] = 1'b1;  wr_cycle[ 7739] = 1'b0;  addr_rom[ 7739]='h00000a70;  wr_data_rom[ 7739]='h00000000;
    rd_cycle[ 7740] = 1'b0;  wr_cycle[ 7740] = 1'b1;  addr_rom[ 7740]='h00001978;  wr_data_rom[ 7740]='h00003d13;
    rd_cycle[ 7741] = 1'b0;  wr_cycle[ 7741] = 1'b1;  addr_rom[ 7741]='h00003fe4;  wr_data_rom[ 7741]='h00002938;
    rd_cycle[ 7742] = 1'b0;  wr_cycle[ 7742] = 1'b1;  addr_rom[ 7742]='h00001568;  wr_data_rom[ 7742]='h0000257b;
    rd_cycle[ 7743] = 1'b0;  wr_cycle[ 7743] = 1'b1;  addr_rom[ 7743]='h00000928;  wr_data_rom[ 7743]='h000022b4;
    rd_cycle[ 7744] = 1'b0;  wr_cycle[ 7744] = 1'b1;  addr_rom[ 7744]='h00002528;  wr_data_rom[ 7744]='h000032e6;
    rd_cycle[ 7745] = 1'b1;  wr_cycle[ 7745] = 1'b0;  addr_rom[ 7745]='h000020e4;  wr_data_rom[ 7745]='h00000000;
    rd_cycle[ 7746] = 1'b0;  wr_cycle[ 7746] = 1'b1;  addr_rom[ 7746]='h00002894;  wr_data_rom[ 7746]='h0000215b;
    rd_cycle[ 7747] = 1'b1;  wr_cycle[ 7747] = 1'b0;  addr_rom[ 7747]='h000001b4;  wr_data_rom[ 7747]='h00000000;
    rd_cycle[ 7748] = 1'b1;  wr_cycle[ 7748] = 1'b0;  addr_rom[ 7748]='h00003588;  wr_data_rom[ 7748]='h00000000;
    rd_cycle[ 7749] = 1'b1;  wr_cycle[ 7749] = 1'b0;  addr_rom[ 7749]='h00003c4c;  wr_data_rom[ 7749]='h00000000;
    rd_cycle[ 7750] = 1'b1;  wr_cycle[ 7750] = 1'b0;  addr_rom[ 7750]='h000015a8;  wr_data_rom[ 7750]='h00000000;
    rd_cycle[ 7751] = 1'b0;  wr_cycle[ 7751] = 1'b1;  addr_rom[ 7751]='h0000280c;  wr_data_rom[ 7751]='h00001811;
    rd_cycle[ 7752] = 1'b0;  wr_cycle[ 7752] = 1'b1;  addr_rom[ 7752]='h000018e4;  wr_data_rom[ 7752]='h00002104;
    rd_cycle[ 7753] = 1'b1;  wr_cycle[ 7753] = 1'b0;  addr_rom[ 7753]='h00000a24;  wr_data_rom[ 7753]='h00000000;
    rd_cycle[ 7754] = 1'b0;  wr_cycle[ 7754] = 1'b1;  addr_rom[ 7754]='h000023d0;  wr_data_rom[ 7754]='h00000a09;
    rd_cycle[ 7755] = 1'b1;  wr_cycle[ 7755] = 1'b0;  addr_rom[ 7755]='h00001dac;  wr_data_rom[ 7755]='h00000000;
    rd_cycle[ 7756] = 1'b0;  wr_cycle[ 7756] = 1'b1;  addr_rom[ 7756]='h00003460;  wr_data_rom[ 7756]='h000029a4;
    rd_cycle[ 7757] = 1'b1;  wr_cycle[ 7757] = 1'b0;  addr_rom[ 7757]='h0000000c;  wr_data_rom[ 7757]='h00000000;
    rd_cycle[ 7758] = 1'b1;  wr_cycle[ 7758] = 1'b0;  addr_rom[ 7758]='h00002b54;  wr_data_rom[ 7758]='h00000000;
    rd_cycle[ 7759] = 1'b1;  wr_cycle[ 7759] = 1'b0;  addr_rom[ 7759]='h00003484;  wr_data_rom[ 7759]='h00000000;
    rd_cycle[ 7760] = 1'b0;  wr_cycle[ 7760] = 1'b1;  addr_rom[ 7760]='h00001f64;  wr_data_rom[ 7760]='h00001dde;
    rd_cycle[ 7761] = 1'b0;  wr_cycle[ 7761] = 1'b1;  addr_rom[ 7761]='h00001d70;  wr_data_rom[ 7761]='h000008aa;
    rd_cycle[ 7762] = 1'b0;  wr_cycle[ 7762] = 1'b1;  addr_rom[ 7762]='h00002f9c;  wr_data_rom[ 7762]='h00001658;
    rd_cycle[ 7763] = 1'b0;  wr_cycle[ 7763] = 1'b1;  addr_rom[ 7763]='h00001778;  wr_data_rom[ 7763]='h000006f6;
    rd_cycle[ 7764] = 1'b1;  wr_cycle[ 7764] = 1'b0;  addr_rom[ 7764]='h00000460;  wr_data_rom[ 7764]='h00000000;
    rd_cycle[ 7765] = 1'b0;  wr_cycle[ 7765] = 1'b1;  addr_rom[ 7765]='h00003f0c;  wr_data_rom[ 7765]='h00001388;
    rd_cycle[ 7766] = 1'b1;  wr_cycle[ 7766] = 1'b0;  addr_rom[ 7766]='h00002d74;  wr_data_rom[ 7766]='h00000000;
    rd_cycle[ 7767] = 1'b1;  wr_cycle[ 7767] = 1'b0;  addr_rom[ 7767]='h000010b8;  wr_data_rom[ 7767]='h00000000;
    rd_cycle[ 7768] = 1'b0;  wr_cycle[ 7768] = 1'b1;  addr_rom[ 7768]='h00002a2c;  wr_data_rom[ 7768]='h00002307;
    rd_cycle[ 7769] = 1'b0;  wr_cycle[ 7769] = 1'b1;  addr_rom[ 7769]='h00000c1c;  wr_data_rom[ 7769]='h000036f6;
    rd_cycle[ 7770] = 1'b1;  wr_cycle[ 7770] = 1'b0;  addr_rom[ 7770]='h00000738;  wr_data_rom[ 7770]='h00000000;
    rd_cycle[ 7771] = 1'b1;  wr_cycle[ 7771] = 1'b0;  addr_rom[ 7771]='h000021d0;  wr_data_rom[ 7771]='h00000000;
    rd_cycle[ 7772] = 1'b0;  wr_cycle[ 7772] = 1'b1;  addr_rom[ 7772]='h00001954;  wr_data_rom[ 7772]='h00000ebc;
    rd_cycle[ 7773] = 1'b0;  wr_cycle[ 7773] = 1'b1;  addr_rom[ 7773]='h00003538;  wr_data_rom[ 7773]='h000007f9;
    rd_cycle[ 7774] = 1'b0;  wr_cycle[ 7774] = 1'b1;  addr_rom[ 7774]='h00001524;  wr_data_rom[ 7774]='h000038cd;
    rd_cycle[ 7775] = 1'b1;  wr_cycle[ 7775] = 1'b0;  addr_rom[ 7775]='h00003c24;  wr_data_rom[ 7775]='h00000000;
    rd_cycle[ 7776] = 1'b0;  wr_cycle[ 7776] = 1'b1;  addr_rom[ 7776]='h00001bd4;  wr_data_rom[ 7776]='h000020a6;
    rd_cycle[ 7777] = 1'b1;  wr_cycle[ 7777] = 1'b0;  addr_rom[ 7777]='h0000139c;  wr_data_rom[ 7777]='h00000000;
    rd_cycle[ 7778] = 1'b1;  wr_cycle[ 7778] = 1'b0;  addr_rom[ 7778]='h00000a04;  wr_data_rom[ 7778]='h00000000;
    rd_cycle[ 7779] = 1'b0;  wr_cycle[ 7779] = 1'b1;  addr_rom[ 7779]='h000020d8;  wr_data_rom[ 7779]='h00003496;
    rd_cycle[ 7780] = 1'b0;  wr_cycle[ 7780] = 1'b1;  addr_rom[ 7780]='h00001a08;  wr_data_rom[ 7780]='h00002bb5;
    rd_cycle[ 7781] = 1'b0;  wr_cycle[ 7781] = 1'b1;  addr_rom[ 7781]='h00002f8c;  wr_data_rom[ 7781]='h0000374e;
    rd_cycle[ 7782] = 1'b0;  wr_cycle[ 7782] = 1'b1;  addr_rom[ 7782]='h00002870;  wr_data_rom[ 7782]='h00002781;
    rd_cycle[ 7783] = 1'b0;  wr_cycle[ 7783] = 1'b1;  addr_rom[ 7783]='h00002308;  wr_data_rom[ 7783]='h00002bf9;
    rd_cycle[ 7784] = 1'b0;  wr_cycle[ 7784] = 1'b1;  addr_rom[ 7784]='h00003c30;  wr_data_rom[ 7784]='h00003459;
    rd_cycle[ 7785] = 1'b0;  wr_cycle[ 7785] = 1'b1;  addr_rom[ 7785]='h00001978;  wr_data_rom[ 7785]='h00002a38;
    rd_cycle[ 7786] = 1'b1;  wr_cycle[ 7786] = 1'b0;  addr_rom[ 7786]='h0000186c;  wr_data_rom[ 7786]='h00000000;
    rd_cycle[ 7787] = 1'b1;  wr_cycle[ 7787] = 1'b0;  addr_rom[ 7787]='h00003e34;  wr_data_rom[ 7787]='h00000000;
    rd_cycle[ 7788] = 1'b0;  wr_cycle[ 7788] = 1'b1;  addr_rom[ 7788]='h00000288;  wr_data_rom[ 7788]='h000035c5;
    rd_cycle[ 7789] = 1'b1;  wr_cycle[ 7789] = 1'b0;  addr_rom[ 7789]='h000015f4;  wr_data_rom[ 7789]='h00000000;
    rd_cycle[ 7790] = 1'b1;  wr_cycle[ 7790] = 1'b0;  addr_rom[ 7790]='h00002594;  wr_data_rom[ 7790]='h00000000;
    rd_cycle[ 7791] = 1'b0;  wr_cycle[ 7791] = 1'b1;  addr_rom[ 7791]='h000025fc;  wr_data_rom[ 7791]='h0000041c;
    rd_cycle[ 7792] = 1'b1;  wr_cycle[ 7792] = 1'b0;  addr_rom[ 7792]='h000018e4;  wr_data_rom[ 7792]='h00000000;
    rd_cycle[ 7793] = 1'b1;  wr_cycle[ 7793] = 1'b0;  addr_rom[ 7793]='h000020cc;  wr_data_rom[ 7793]='h00000000;
    rd_cycle[ 7794] = 1'b0;  wr_cycle[ 7794] = 1'b1;  addr_rom[ 7794]='h000032c4;  wr_data_rom[ 7794]='h00002040;
    rd_cycle[ 7795] = 1'b0;  wr_cycle[ 7795] = 1'b1;  addr_rom[ 7795]='h00000a3c;  wr_data_rom[ 7795]='h000008f4;
    rd_cycle[ 7796] = 1'b0;  wr_cycle[ 7796] = 1'b1;  addr_rom[ 7796]='h00003e94;  wr_data_rom[ 7796]='h000026c7;
    rd_cycle[ 7797] = 1'b0;  wr_cycle[ 7797] = 1'b1;  addr_rom[ 7797]='h0000293c;  wr_data_rom[ 7797]='h0000236f;
    rd_cycle[ 7798] = 1'b0;  wr_cycle[ 7798] = 1'b1;  addr_rom[ 7798]='h000007d4;  wr_data_rom[ 7798]='h0000032e;
    rd_cycle[ 7799] = 1'b1;  wr_cycle[ 7799] = 1'b0;  addr_rom[ 7799]='h00002e78;  wr_data_rom[ 7799]='h00000000;
    rd_cycle[ 7800] = 1'b1;  wr_cycle[ 7800] = 1'b0;  addr_rom[ 7800]='h00001bf8;  wr_data_rom[ 7800]='h00000000;
    rd_cycle[ 7801] = 1'b0;  wr_cycle[ 7801] = 1'b1;  addr_rom[ 7801]='h000018e8;  wr_data_rom[ 7801]='h0000320a;
    rd_cycle[ 7802] = 1'b0;  wr_cycle[ 7802] = 1'b1;  addr_rom[ 7802]='h00003690;  wr_data_rom[ 7802]='h00003db3;
    rd_cycle[ 7803] = 1'b0;  wr_cycle[ 7803] = 1'b1;  addr_rom[ 7803]='h00001d00;  wr_data_rom[ 7803]='h00002732;
    rd_cycle[ 7804] = 1'b0;  wr_cycle[ 7804] = 1'b1;  addr_rom[ 7804]='h000027a8;  wr_data_rom[ 7804]='h000032d2;
    rd_cycle[ 7805] = 1'b1;  wr_cycle[ 7805] = 1'b0;  addr_rom[ 7805]='h0000230c;  wr_data_rom[ 7805]='h00000000;
    rd_cycle[ 7806] = 1'b1;  wr_cycle[ 7806] = 1'b0;  addr_rom[ 7806]='h00003d9c;  wr_data_rom[ 7806]='h00000000;
    rd_cycle[ 7807] = 1'b0;  wr_cycle[ 7807] = 1'b1;  addr_rom[ 7807]='h00003810;  wr_data_rom[ 7807]='h00001c69;
    rd_cycle[ 7808] = 1'b0;  wr_cycle[ 7808] = 1'b1;  addr_rom[ 7808]='h000001f0;  wr_data_rom[ 7808]='h0000248f;
    rd_cycle[ 7809] = 1'b1;  wr_cycle[ 7809] = 1'b0;  addr_rom[ 7809]='h00001294;  wr_data_rom[ 7809]='h00000000;
    rd_cycle[ 7810] = 1'b1;  wr_cycle[ 7810] = 1'b0;  addr_rom[ 7810]='h000021ac;  wr_data_rom[ 7810]='h00000000;
    rd_cycle[ 7811] = 1'b0;  wr_cycle[ 7811] = 1'b1;  addr_rom[ 7811]='h00003890;  wr_data_rom[ 7811]='h00003110;
    rd_cycle[ 7812] = 1'b0;  wr_cycle[ 7812] = 1'b1;  addr_rom[ 7812]='h000034f4;  wr_data_rom[ 7812]='h000001cb;
    rd_cycle[ 7813] = 1'b1;  wr_cycle[ 7813] = 1'b0;  addr_rom[ 7813]='h000028f0;  wr_data_rom[ 7813]='h00000000;
    rd_cycle[ 7814] = 1'b1;  wr_cycle[ 7814] = 1'b0;  addr_rom[ 7814]='h00002448;  wr_data_rom[ 7814]='h00000000;
    rd_cycle[ 7815] = 1'b1;  wr_cycle[ 7815] = 1'b0;  addr_rom[ 7815]='h00000898;  wr_data_rom[ 7815]='h00000000;
    rd_cycle[ 7816] = 1'b0;  wr_cycle[ 7816] = 1'b1;  addr_rom[ 7816]='h00001ca4;  wr_data_rom[ 7816]='h000024e2;
    rd_cycle[ 7817] = 1'b1;  wr_cycle[ 7817] = 1'b0;  addr_rom[ 7817]='h00002cb4;  wr_data_rom[ 7817]='h00000000;
    rd_cycle[ 7818] = 1'b1;  wr_cycle[ 7818] = 1'b0;  addr_rom[ 7818]='h0000289c;  wr_data_rom[ 7818]='h00000000;
    rd_cycle[ 7819] = 1'b0;  wr_cycle[ 7819] = 1'b1;  addr_rom[ 7819]='h00000fc0;  wr_data_rom[ 7819]='h000011f2;
    rd_cycle[ 7820] = 1'b0;  wr_cycle[ 7820] = 1'b1;  addr_rom[ 7820]='h00002f64;  wr_data_rom[ 7820]='h00000003;
    rd_cycle[ 7821] = 1'b1;  wr_cycle[ 7821] = 1'b0;  addr_rom[ 7821]='h00000ed4;  wr_data_rom[ 7821]='h00000000;
    rd_cycle[ 7822] = 1'b0;  wr_cycle[ 7822] = 1'b1;  addr_rom[ 7822]='h00000338;  wr_data_rom[ 7822]='h000002ba;
    rd_cycle[ 7823] = 1'b0;  wr_cycle[ 7823] = 1'b1;  addr_rom[ 7823]='h00000cdc;  wr_data_rom[ 7823]='h00002955;
    rd_cycle[ 7824] = 1'b1;  wr_cycle[ 7824] = 1'b0;  addr_rom[ 7824]='h0000155c;  wr_data_rom[ 7824]='h00000000;
    rd_cycle[ 7825] = 1'b1;  wr_cycle[ 7825] = 1'b0;  addr_rom[ 7825]='h00001104;  wr_data_rom[ 7825]='h00000000;
    rd_cycle[ 7826] = 1'b0;  wr_cycle[ 7826] = 1'b1;  addr_rom[ 7826]='h000001a8;  wr_data_rom[ 7826]='h0000346e;
    rd_cycle[ 7827] = 1'b0;  wr_cycle[ 7827] = 1'b1;  addr_rom[ 7827]='h000022dc;  wr_data_rom[ 7827]='h0000258c;
    rd_cycle[ 7828] = 1'b1;  wr_cycle[ 7828] = 1'b0;  addr_rom[ 7828]='h0000124c;  wr_data_rom[ 7828]='h00000000;
    rd_cycle[ 7829] = 1'b1;  wr_cycle[ 7829] = 1'b0;  addr_rom[ 7829]='h00000794;  wr_data_rom[ 7829]='h00000000;
    rd_cycle[ 7830] = 1'b0;  wr_cycle[ 7830] = 1'b1;  addr_rom[ 7830]='h000020ac;  wr_data_rom[ 7830]='h00002632;
    rd_cycle[ 7831] = 1'b1;  wr_cycle[ 7831] = 1'b0;  addr_rom[ 7831]='h000028c4;  wr_data_rom[ 7831]='h00000000;
    rd_cycle[ 7832] = 1'b0;  wr_cycle[ 7832] = 1'b1;  addr_rom[ 7832]='h00000cc8;  wr_data_rom[ 7832]='h000021a3;
    rd_cycle[ 7833] = 1'b0;  wr_cycle[ 7833] = 1'b1;  addr_rom[ 7833]='h00001494;  wr_data_rom[ 7833]='h00000a66;
    rd_cycle[ 7834] = 1'b0;  wr_cycle[ 7834] = 1'b1;  addr_rom[ 7834]='h00000f9c;  wr_data_rom[ 7834]='h00003f73;
    rd_cycle[ 7835] = 1'b1;  wr_cycle[ 7835] = 1'b0;  addr_rom[ 7835]='h00003838;  wr_data_rom[ 7835]='h00000000;
    rd_cycle[ 7836] = 1'b1;  wr_cycle[ 7836] = 1'b0;  addr_rom[ 7836]='h00002fa8;  wr_data_rom[ 7836]='h00000000;
    rd_cycle[ 7837] = 1'b1;  wr_cycle[ 7837] = 1'b0;  addr_rom[ 7837]='h00000c44;  wr_data_rom[ 7837]='h00000000;
    rd_cycle[ 7838] = 1'b1;  wr_cycle[ 7838] = 1'b0;  addr_rom[ 7838]='h00003aa0;  wr_data_rom[ 7838]='h00000000;
    rd_cycle[ 7839] = 1'b0;  wr_cycle[ 7839] = 1'b1;  addr_rom[ 7839]='h00000e84;  wr_data_rom[ 7839]='h00000f2c;
    rd_cycle[ 7840] = 1'b0;  wr_cycle[ 7840] = 1'b1;  addr_rom[ 7840]='h00001620;  wr_data_rom[ 7840]='h00003178;
    rd_cycle[ 7841] = 1'b1;  wr_cycle[ 7841] = 1'b0;  addr_rom[ 7841]='h000019c4;  wr_data_rom[ 7841]='h00000000;
    rd_cycle[ 7842] = 1'b0;  wr_cycle[ 7842] = 1'b1;  addr_rom[ 7842]='h00001194;  wr_data_rom[ 7842]='h00001963;
    rd_cycle[ 7843] = 1'b0;  wr_cycle[ 7843] = 1'b1;  addr_rom[ 7843]='h00001fd4;  wr_data_rom[ 7843]='h000028bc;
    rd_cycle[ 7844] = 1'b0;  wr_cycle[ 7844] = 1'b1;  addr_rom[ 7844]='h00002b10;  wr_data_rom[ 7844]='h000023d9;
    rd_cycle[ 7845] = 1'b0;  wr_cycle[ 7845] = 1'b1;  addr_rom[ 7845]='h00002f20;  wr_data_rom[ 7845]='h00003c39;
    rd_cycle[ 7846] = 1'b0;  wr_cycle[ 7846] = 1'b1;  addr_rom[ 7846]='h00001984;  wr_data_rom[ 7846]='h00000032;
    rd_cycle[ 7847] = 1'b1;  wr_cycle[ 7847] = 1'b0;  addr_rom[ 7847]='h00003214;  wr_data_rom[ 7847]='h00000000;
    rd_cycle[ 7848] = 1'b0;  wr_cycle[ 7848] = 1'b1;  addr_rom[ 7848]='h00001ba0;  wr_data_rom[ 7848]='h00000547;
    rd_cycle[ 7849] = 1'b1;  wr_cycle[ 7849] = 1'b0;  addr_rom[ 7849]='h00002a8c;  wr_data_rom[ 7849]='h00000000;
    rd_cycle[ 7850] = 1'b1;  wr_cycle[ 7850] = 1'b0;  addr_rom[ 7850]='h0000091c;  wr_data_rom[ 7850]='h00000000;
    rd_cycle[ 7851] = 1'b1;  wr_cycle[ 7851] = 1'b0;  addr_rom[ 7851]='h00000c90;  wr_data_rom[ 7851]='h00000000;
    rd_cycle[ 7852] = 1'b1;  wr_cycle[ 7852] = 1'b0;  addr_rom[ 7852]='h00000628;  wr_data_rom[ 7852]='h00000000;
    rd_cycle[ 7853] = 1'b0;  wr_cycle[ 7853] = 1'b1;  addr_rom[ 7853]='h000037a8;  wr_data_rom[ 7853]='h0000265b;
    rd_cycle[ 7854] = 1'b1;  wr_cycle[ 7854] = 1'b0;  addr_rom[ 7854]='h000009c0;  wr_data_rom[ 7854]='h00000000;
    rd_cycle[ 7855] = 1'b0;  wr_cycle[ 7855] = 1'b1;  addr_rom[ 7855]='h00002458;  wr_data_rom[ 7855]='h00002420;
    rd_cycle[ 7856] = 1'b0;  wr_cycle[ 7856] = 1'b1;  addr_rom[ 7856]='h00003c38;  wr_data_rom[ 7856]='h00002a28;
    rd_cycle[ 7857] = 1'b0;  wr_cycle[ 7857] = 1'b1;  addr_rom[ 7857]='h00000c38;  wr_data_rom[ 7857]='h00002325;
    rd_cycle[ 7858] = 1'b0;  wr_cycle[ 7858] = 1'b1;  addr_rom[ 7858]='h00001fa0;  wr_data_rom[ 7858]='h00000507;
    rd_cycle[ 7859] = 1'b1;  wr_cycle[ 7859] = 1'b0;  addr_rom[ 7859]='h00000dd0;  wr_data_rom[ 7859]='h00000000;
    rd_cycle[ 7860] = 1'b0;  wr_cycle[ 7860] = 1'b1;  addr_rom[ 7860]='h00002274;  wr_data_rom[ 7860]='h00001b38;
    rd_cycle[ 7861] = 1'b1;  wr_cycle[ 7861] = 1'b0;  addr_rom[ 7861]='h00002568;  wr_data_rom[ 7861]='h00000000;
    rd_cycle[ 7862] = 1'b0;  wr_cycle[ 7862] = 1'b1;  addr_rom[ 7862]='h00001cc4;  wr_data_rom[ 7862]='h00001ca9;
    rd_cycle[ 7863] = 1'b0;  wr_cycle[ 7863] = 1'b1;  addr_rom[ 7863]='h00000e9c;  wr_data_rom[ 7863]='h000036fc;
    rd_cycle[ 7864] = 1'b0;  wr_cycle[ 7864] = 1'b1;  addr_rom[ 7864]='h00000f40;  wr_data_rom[ 7864]='h00001fa9;
    rd_cycle[ 7865] = 1'b0;  wr_cycle[ 7865] = 1'b1;  addr_rom[ 7865]='h00002abc;  wr_data_rom[ 7865]='h00001a80;
    rd_cycle[ 7866] = 1'b1;  wr_cycle[ 7866] = 1'b0;  addr_rom[ 7866]='h00002148;  wr_data_rom[ 7866]='h00000000;
    rd_cycle[ 7867] = 1'b1;  wr_cycle[ 7867] = 1'b0;  addr_rom[ 7867]='h000020e4;  wr_data_rom[ 7867]='h00000000;
    rd_cycle[ 7868] = 1'b0;  wr_cycle[ 7868] = 1'b1;  addr_rom[ 7868]='h00002d84;  wr_data_rom[ 7868]='h00001213;
    rd_cycle[ 7869] = 1'b0;  wr_cycle[ 7869] = 1'b1;  addr_rom[ 7869]='h00000080;  wr_data_rom[ 7869]='h00001948;
    rd_cycle[ 7870] = 1'b1;  wr_cycle[ 7870] = 1'b0;  addr_rom[ 7870]='h000020a8;  wr_data_rom[ 7870]='h00000000;
    rd_cycle[ 7871] = 1'b1;  wr_cycle[ 7871] = 1'b0;  addr_rom[ 7871]='h00001d48;  wr_data_rom[ 7871]='h00000000;
    rd_cycle[ 7872] = 1'b1;  wr_cycle[ 7872] = 1'b0;  addr_rom[ 7872]='h00002ecc;  wr_data_rom[ 7872]='h00000000;
    rd_cycle[ 7873] = 1'b1;  wr_cycle[ 7873] = 1'b0;  addr_rom[ 7873]='h00001a10;  wr_data_rom[ 7873]='h00000000;
    rd_cycle[ 7874] = 1'b1;  wr_cycle[ 7874] = 1'b0;  addr_rom[ 7874]='h000011f0;  wr_data_rom[ 7874]='h00000000;
    rd_cycle[ 7875] = 1'b0;  wr_cycle[ 7875] = 1'b1;  addr_rom[ 7875]='h0000357c;  wr_data_rom[ 7875]='h00000f8e;
    rd_cycle[ 7876] = 1'b0;  wr_cycle[ 7876] = 1'b1;  addr_rom[ 7876]='h00002048;  wr_data_rom[ 7876]='h00002f0a;
    rd_cycle[ 7877] = 1'b0;  wr_cycle[ 7877] = 1'b1;  addr_rom[ 7877]='h000002b0;  wr_data_rom[ 7877]='h000032be;
    rd_cycle[ 7878] = 1'b1;  wr_cycle[ 7878] = 1'b0;  addr_rom[ 7878]='h00001c7c;  wr_data_rom[ 7878]='h00000000;
    rd_cycle[ 7879] = 1'b0;  wr_cycle[ 7879] = 1'b1;  addr_rom[ 7879]='h000025f4;  wr_data_rom[ 7879]='h000007c1;
    rd_cycle[ 7880] = 1'b0;  wr_cycle[ 7880] = 1'b1;  addr_rom[ 7880]='h00003be0;  wr_data_rom[ 7880]='h000038fe;
    rd_cycle[ 7881] = 1'b1;  wr_cycle[ 7881] = 1'b0;  addr_rom[ 7881]='h000009b4;  wr_data_rom[ 7881]='h00000000;
    rd_cycle[ 7882] = 1'b0;  wr_cycle[ 7882] = 1'b1;  addr_rom[ 7882]='h000002f8;  wr_data_rom[ 7882]='h0000132d;
    rd_cycle[ 7883] = 1'b0;  wr_cycle[ 7883] = 1'b1;  addr_rom[ 7883]='h000010dc;  wr_data_rom[ 7883]='h0000379b;
    rd_cycle[ 7884] = 1'b0;  wr_cycle[ 7884] = 1'b1;  addr_rom[ 7884]='h00000b40;  wr_data_rom[ 7884]='h00002cb3;
    rd_cycle[ 7885] = 1'b1;  wr_cycle[ 7885] = 1'b0;  addr_rom[ 7885]='h00000b74;  wr_data_rom[ 7885]='h00000000;
    rd_cycle[ 7886] = 1'b0;  wr_cycle[ 7886] = 1'b1;  addr_rom[ 7886]='h00003f70;  wr_data_rom[ 7886]='h00001835;
    rd_cycle[ 7887] = 1'b1;  wr_cycle[ 7887] = 1'b0;  addr_rom[ 7887]='h00000dcc;  wr_data_rom[ 7887]='h00000000;
    rd_cycle[ 7888] = 1'b1;  wr_cycle[ 7888] = 1'b0;  addr_rom[ 7888]='h000004dc;  wr_data_rom[ 7888]='h00000000;
    rd_cycle[ 7889] = 1'b0;  wr_cycle[ 7889] = 1'b1;  addr_rom[ 7889]='h000026fc;  wr_data_rom[ 7889]='h00002c7e;
    rd_cycle[ 7890] = 1'b0;  wr_cycle[ 7890] = 1'b1;  addr_rom[ 7890]='h000016a8;  wr_data_rom[ 7890]='h00003f90;
    rd_cycle[ 7891] = 1'b0;  wr_cycle[ 7891] = 1'b1;  addr_rom[ 7891]='h000009e4;  wr_data_rom[ 7891]='h00003598;
    rd_cycle[ 7892] = 1'b0;  wr_cycle[ 7892] = 1'b1;  addr_rom[ 7892]='h00002d10;  wr_data_rom[ 7892]='h00003daf;
    rd_cycle[ 7893] = 1'b0;  wr_cycle[ 7893] = 1'b1;  addr_rom[ 7893]='h000008b8;  wr_data_rom[ 7893]='h000024ab;
    rd_cycle[ 7894] = 1'b1;  wr_cycle[ 7894] = 1'b0;  addr_rom[ 7894]='h00002cc4;  wr_data_rom[ 7894]='h00000000;
    rd_cycle[ 7895] = 1'b0;  wr_cycle[ 7895] = 1'b1;  addr_rom[ 7895]='h0000307c;  wr_data_rom[ 7895]='h00002cdf;
    rd_cycle[ 7896] = 1'b0;  wr_cycle[ 7896] = 1'b1;  addr_rom[ 7896]='h00000030;  wr_data_rom[ 7896]='h00003c66;
    rd_cycle[ 7897] = 1'b0;  wr_cycle[ 7897] = 1'b1;  addr_rom[ 7897]='h00001944;  wr_data_rom[ 7897]='h0000273b;
    rd_cycle[ 7898] = 1'b0;  wr_cycle[ 7898] = 1'b1;  addr_rom[ 7898]='h00001aa0;  wr_data_rom[ 7898]='h000003f5;
    rd_cycle[ 7899] = 1'b0;  wr_cycle[ 7899] = 1'b1;  addr_rom[ 7899]='h00003a08;  wr_data_rom[ 7899]='h00000b91;
    rd_cycle[ 7900] = 1'b1;  wr_cycle[ 7900] = 1'b0;  addr_rom[ 7900]='h00001320;  wr_data_rom[ 7900]='h00000000;
    rd_cycle[ 7901] = 1'b1;  wr_cycle[ 7901] = 1'b0;  addr_rom[ 7901]='h00000e3c;  wr_data_rom[ 7901]='h00000000;
    rd_cycle[ 7902] = 1'b0;  wr_cycle[ 7902] = 1'b1;  addr_rom[ 7902]='h00002ebc;  wr_data_rom[ 7902]='h000010db;
    rd_cycle[ 7903] = 1'b1;  wr_cycle[ 7903] = 1'b0;  addr_rom[ 7903]='h00003650;  wr_data_rom[ 7903]='h00000000;
    rd_cycle[ 7904] = 1'b1;  wr_cycle[ 7904] = 1'b0;  addr_rom[ 7904]='h00002548;  wr_data_rom[ 7904]='h00000000;
    rd_cycle[ 7905] = 1'b0;  wr_cycle[ 7905] = 1'b1;  addr_rom[ 7905]='h00002158;  wr_data_rom[ 7905]='h00000271;
    rd_cycle[ 7906] = 1'b1;  wr_cycle[ 7906] = 1'b0;  addr_rom[ 7906]='h00001ad4;  wr_data_rom[ 7906]='h00000000;
    rd_cycle[ 7907] = 1'b0;  wr_cycle[ 7907] = 1'b1;  addr_rom[ 7907]='h000026c4;  wr_data_rom[ 7907]='h00001f9c;
    rd_cycle[ 7908] = 1'b0;  wr_cycle[ 7908] = 1'b1;  addr_rom[ 7908]='h00000ea0;  wr_data_rom[ 7908]='h000019c6;
    rd_cycle[ 7909] = 1'b0;  wr_cycle[ 7909] = 1'b1;  addr_rom[ 7909]='h000018b8;  wr_data_rom[ 7909]='h00001d9b;
    rd_cycle[ 7910] = 1'b1;  wr_cycle[ 7910] = 1'b0;  addr_rom[ 7910]='h00001760;  wr_data_rom[ 7910]='h00000000;
    rd_cycle[ 7911] = 1'b1;  wr_cycle[ 7911] = 1'b0;  addr_rom[ 7911]='h0000083c;  wr_data_rom[ 7911]='h00000000;
    rd_cycle[ 7912] = 1'b0;  wr_cycle[ 7912] = 1'b1;  addr_rom[ 7912]='h00003a60;  wr_data_rom[ 7912]='h000030e4;
    rd_cycle[ 7913] = 1'b1;  wr_cycle[ 7913] = 1'b0;  addr_rom[ 7913]='h00003d14;  wr_data_rom[ 7913]='h00000000;
    rd_cycle[ 7914] = 1'b1;  wr_cycle[ 7914] = 1'b0;  addr_rom[ 7914]='h00002ab0;  wr_data_rom[ 7914]='h00000000;
    rd_cycle[ 7915] = 1'b0;  wr_cycle[ 7915] = 1'b1;  addr_rom[ 7915]='h000007f8;  wr_data_rom[ 7915]='h00002a73;
    rd_cycle[ 7916] = 1'b1;  wr_cycle[ 7916] = 1'b0;  addr_rom[ 7916]='h000025a4;  wr_data_rom[ 7916]='h00000000;
    rd_cycle[ 7917] = 1'b1;  wr_cycle[ 7917] = 1'b0;  addr_rom[ 7917]='h00002f68;  wr_data_rom[ 7917]='h00000000;
    rd_cycle[ 7918] = 1'b1;  wr_cycle[ 7918] = 1'b0;  addr_rom[ 7918]='h00002de8;  wr_data_rom[ 7918]='h00000000;
    rd_cycle[ 7919] = 1'b0;  wr_cycle[ 7919] = 1'b1;  addr_rom[ 7919]='h00002170;  wr_data_rom[ 7919]='h000016a2;
    rd_cycle[ 7920] = 1'b1;  wr_cycle[ 7920] = 1'b0;  addr_rom[ 7920]='h00002790;  wr_data_rom[ 7920]='h00000000;
    rd_cycle[ 7921] = 1'b1;  wr_cycle[ 7921] = 1'b0;  addr_rom[ 7921]='h000002ec;  wr_data_rom[ 7921]='h00000000;
    rd_cycle[ 7922] = 1'b0;  wr_cycle[ 7922] = 1'b1;  addr_rom[ 7922]='h00001610;  wr_data_rom[ 7922]='h00000c28;
    rd_cycle[ 7923] = 1'b0;  wr_cycle[ 7923] = 1'b1;  addr_rom[ 7923]='h00002860;  wr_data_rom[ 7923]='h000021ff;
    rd_cycle[ 7924] = 1'b1;  wr_cycle[ 7924] = 1'b0;  addr_rom[ 7924]='h00003098;  wr_data_rom[ 7924]='h00000000;
    rd_cycle[ 7925] = 1'b0;  wr_cycle[ 7925] = 1'b1;  addr_rom[ 7925]='h00003418;  wr_data_rom[ 7925]='h00001450;
    rd_cycle[ 7926] = 1'b1;  wr_cycle[ 7926] = 1'b0;  addr_rom[ 7926]='h00000390;  wr_data_rom[ 7926]='h00000000;
    rd_cycle[ 7927] = 1'b1;  wr_cycle[ 7927] = 1'b0;  addr_rom[ 7927]='h00000cdc;  wr_data_rom[ 7927]='h00000000;
    rd_cycle[ 7928] = 1'b1;  wr_cycle[ 7928] = 1'b0;  addr_rom[ 7928]='h00001574;  wr_data_rom[ 7928]='h00000000;
    rd_cycle[ 7929] = 1'b0;  wr_cycle[ 7929] = 1'b1;  addr_rom[ 7929]='h0000141c;  wr_data_rom[ 7929]='h00003fc3;
    rd_cycle[ 7930] = 1'b1;  wr_cycle[ 7930] = 1'b0;  addr_rom[ 7930]='h00002168;  wr_data_rom[ 7930]='h00000000;
    rd_cycle[ 7931] = 1'b0;  wr_cycle[ 7931] = 1'b1;  addr_rom[ 7931]='h00000e24;  wr_data_rom[ 7931]='h00002c3a;
    rd_cycle[ 7932] = 1'b0;  wr_cycle[ 7932] = 1'b1;  addr_rom[ 7932]='h00001c04;  wr_data_rom[ 7932]='h00002e75;
    rd_cycle[ 7933] = 1'b0;  wr_cycle[ 7933] = 1'b1;  addr_rom[ 7933]='h00002fd0;  wr_data_rom[ 7933]='h00000c92;
    rd_cycle[ 7934] = 1'b1;  wr_cycle[ 7934] = 1'b0;  addr_rom[ 7934]='h00000320;  wr_data_rom[ 7934]='h00000000;
    rd_cycle[ 7935] = 1'b0;  wr_cycle[ 7935] = 1'b1;  addr_rom[ 7935]='h00001818;  wr_data_rom[ 7935]='h00002984;
    rd_cycle[ 7936] = 1'b1;  wr_cycle[ 7936] = 1'b0;  addr_rom[ 7936]='h00001974;  wr_data_rom[ 7936]='h00000000;
    rd_cycle[ 7937] = 1'b1;  wr_cycle[ 7937] = 1'b0;  addr_rom[ 7937]='h000030d4;  wr_data_rom[ 7937]='h00000000;
    rd_cycle[ 7938] = 1'b1;  wr_cycle[ 7938] = 1'b0;  addr_rom[ 7938]='h000038d8;  wr_data_rom[ 7938]='h00000000;
    rd_cycle[ 7939] = 1'b0;  wr_cycle[ 7939] = 1'b1;  addr_rom[ 7939]='h00001bac;  wr_data_rom[ 7939]='h00002a08;
    rd_cycle[ 7940] = 1'b0;  wr_cycle[ 7940] = 1'b1;  addr_rom[ 7940]='h00003058;  wr_data_rom[ 7940]='h00003966;
    rd_cycle[ 7941] = 1'b1;  wr_cycle[ 7941] = 1'b0;  addr_rom[ 7941]='h00000670;  wr_data_rom[ 7941]='h00000000;
    rd_cycle[ 7942] = 1'b0;  wr_cycle[ 7942] = 1'b1;  addr_rom[ 7942]='h000011ec;  wr_data_rom[ 7942]='h00003ceb;
    rd_cycle[ 7943] = 1'b1;  wr_cycle[ 7943] = 1'b0;  addr_rom[ 7943]='h0000046c;  wr_data_rom[ 7943]='h00000000;
    rd_cycle[ 7944] = 1'b0;  wr_cycle[ 7944] = 1'b1;  addr_rom[ 7944]='h00001f88;  wr_data_rom[ 7944]='h00000441;
    rd_cycle[ 7945] = 1'b1;  wr_cycle[ 7945] = 1'b0;  addr_rom[ 7945]='h00003560;  wr_data_rom[ 7945]='h00000000;
    rd_cycle[ 7946] = 1'b0;  wr_cycle[ 7946] = 1'b1;  addr_rom[ 7946]='h00001f60;  wr_data_rom[ 7946]='h00003ef9;
    rd_cycle[ 7947] = 1'b0;  wr_cycle[ 7947] = 1'b1;  addr_rom[ 7947]='h00000110;  wr_data_rom[ 7947]='h000013a6;
    rd_cycle[ 7948] = 1'b1;  wr_cycle[ 7948] = 1'b0;  addr_rom[ 7948]='h00003d9c;  wr_data_rom[ 7948]='h00000000;
    rd_cycle[ 7949] = 1'b0;  wr_cycle[ 7949] = 1'b1;  addr_rom[ 7949]='h000030b0;  wr_data_rom[ 7949]='h000006a3;
    rd_cycle[ 7950] = 1'b0;  wr_cycle[ 7950] = 1'b1;  addr_rom[ 7950]='h000008f8;  wr_data_rom[ 7950]='h00001b21;
    rd_cycle[ 7951] = 1'b0;  wr_cycle[ 7951] = 1'b1;  addr_rom[ 7951]='h00001d34;  wr_data_rom[ 7951]='h000035a1;
    rd_cycle[ 7952] = 1'b0;  wr_cycle[ 7952] = 1'b1;  addr_rom[ 7952]='h00000e70;  wr_data_rom[ 7952]='h00003f08;
    rd_cycle[ 7953] = 1'b1;  wr_cycle[ 7953] = 1'b0;  addr_rom[ 7953]='h00003fd0;  wr_data_rom[ 7953]='h00000000;
    rd_cycle[ 7954] = 1'b0;  wr_cycle[ 7954] = 1'b1;  addr_rom[ 7954]='h00000d7c;  wr_data_rom[ 7954]='h00003d0a;
    rd_cycle[ 7955] = 1'b1;  wr_cycle[ 7955] = 1'b0;  addr_rom[ 7955]='h00001a48;  wr_data_rom[ 7955]='h00000000;
    rd_cycle[ 7956] = 1'b0;  wr_cycle[ 7956] = 1'b1;  addr_rom[ 7956]='h00000540;  wr_data_rom[ 7956]='h00002664;
    rd_cycle[ 7957] = 1'b0;  wr_cycle[ 7957] = 1'b1;  addr_rom[ 7957]='h000025a4;  wr_data_rom[ 7957]='h00001927;
    rd_cycle[ 7958] = 1'b0;  wr_cycle[ 7958] = 1'b1;  addr_rom[ 7958]='h00001250;  wr_data_rom[ 7958]='h0000226f;
    rd_cycle[ 7959] = 1'b1;  wr_cycle[ 7959] = 1'b0;  addr_rom[ 7959]='h00000398;  wr_data_rom[ 7959]='h00000000;
    rd_cycle[ 7960] = 1'b0;  wr_cycle[ 7960] = 1'b1;  addr_rom[ 7960]='h00001134;  wr_data_rom[ 7960]='h00003bfd;
    rd_cycle[ 7961] = 1'b0;  wr_cycle[ 7961] = 1'b1;  addr_rom[ 7961]='h0000019c;  wr_data_rom[ 7961]='h0000243b;
    rd_cycle[ 7962] = 1'b0;  wr_cycle[ 7962] = 1'b1;  addr_rom[ 7962]='h00003898;  wr_data_rom[ 7962]='h000018d0;
    rd_cycle[ 7963] = 1'b1;  wr_cycle[ 7963] = 1'b0;  addr_rom[ 7963]='h00000444;  wr_data_rom[ 7963]='h00000000;
    rd_cycle[ 7964] = 1'b0;  wr_cycle[ 7964] = 1'b1;  addr_rom[ 7964]='h00003820;  wr_data_rom[ 7964]='h000012c7;
    rd_cycle[ 7965] = 1'b0;  wr_cycle[ 7965] = 1'b1;  addr_rom[ 7965]='h00003a2c;  wr_data_rom[ 7965]='h00000469;
    rd_cycle[ 7966] = 1'b0;  wr_cycle[ 7966] = 1'b1;  addr_rom[ 7966]='h00001d1c;  wr_data_rom[ 7966]='h0000204f;
    rd_cycle[ 7967] = 1'b0;  wr_cycle[ 7967] = 1'b1;  addr_rom[ 7967]='h00003e40;  wr_data_rom[ 7967]='h00001a65;
    rd_cycle[ 7968] = 1'b0;  wr_cycle[ 7968] = 1'b1;  addr_rom[ 7968]='h000035a0;  wr_data_rom[ 7968]='h00000bb4;
    rd_cycle[ 7969] = 1'b1;  wr_cycle[ 7969] = 1'b0;  addr_rom[ 7969]='h000031b4;  wr_data_rom[ 7969]='h00000000;
    rd_cycle[ 7970] = 1'b0;  wr_cycle[ 7970] = 1'b1;  addr_rom[ 7970]='h00000108;  wr_data_rom[ 7970]='h00003428;
    rd_cycle[ 7971] = 1'b0;  wr_cycle[ 7971] = 1'b1;  addr_rom[ 7971]='h00000db4;  wr_data_rom[ 7971]='h000002a5;
    rd_cycle[ 7972] = 1'b1;  wr_cycle[ 7972] = 1'b0;  addr_rom[ 7972]='h000004c0;  wr_data_rom[ 7972]='h00000000;
    rd_cycle[ 7973] = 1'b1;  wr_cycle[ 7973] = 1'b0;  addr_rom[ 7973]='h00002f9c;  wr_data_rom[ 7973]='h00000000;
    rd_cycle[ 7974] = 1'b1;  wr_cycle[ 7974] = 1'b0;  addr_rom[ 7974]='h00000b1c;  wr_data_rom[ 7974]='h00000000;
    rd_cycle[ 7975] = 1'b1;  wr_cycle[ 7975] = 1'b0;  addr_rom[ 7975]='h000020d8;  wr_data_rom[ 7975]='h00000000;
    rd_cycle[ 7976] = 1'b0;  wr_cycle[ 7976] = 1'b1;  addr_rom[ 7976]='h00002a08;  wr_data_rom[ 7976]='h000023c8;
    rd_cycle[ 7977] = 1'b0;  wr_cycle[ 7977] = 1'b1;  addr_rom[ 7977]='h000008d0;  wr_data_rom[ 7977]='h00002512;
    rd_cycle[ 7978] = 1'b0;  wr_cycle[ 7978] = 1'b1;  addr_rom[ 7978]='h00003730;  wr_data_rom[ 7978]='h00000c77;
    rd_cycle[ 7979] = 1'b1;  wr_cycle[ 7979] = 1'b0;  addr_rom[ 7979]='h000002c4;  wr_data_rom[ 7979]='h00000000;
    rd_cycle[ 7980] = 1'b0;  wr_cycle[ 7980] = 1'b1;  addr_rom[ 7980]='h00001ef8;  wr_data_rom[ 7980]='h00002a7e;
    rd_cycle[ 7981] = 1'b1;  wr_cycle[ 7981] = 1'b0;  addr_rom[ 7981]='h00003220;  wr_data_rom[ 7981]='h00000000;
    rd_cycle[ 7982] = 1'b0;  wr_cycle[ 7982] = 1'b1;  addr_rom[ 7982]='h00002624;  wr_data_rom[ 7982]='h000033a8;
    rd_cycle[ 7983] = 1'b1;  wr_cycle[ 7983] = 1'b0;  addr_rom[ 7983]='h0000065c;  wr_data_rom[ 7983]='h00000000;
    rd_cycle[ 7984] = 1'b0;  wr_cycle[ 7984] = 1'b1;  addr_rom[ 7984]='h00000b3c;  wr_data_rom[ 7984]='h00003868;
    rd_cycle[ 7985] = 1'b1;  wr_cycle[ 7985] = 1'b0;  addr_rom[ 7985]='h00003228;  wr_data_rom[ 7985]='h00000000;
    rd_cycle[ 7986] = 1'b0;  wr_cycle[ 7986] = 1'b1;  addr_rom[ 7986]='h000019cc;  wr_data_rom[ 7986]='h00001b69;
    rd_cycle[ 7987] = 1'b1;  wr_cycle[ 7987] = 1'b0;  addr_rom[ 7987]='h00002330;  wr_data_rom[ 7987]='h00000000;
    rd_cycle[ 7988] = 1'b0;  wr_cycle[ 7988] = 1'b1;  addr_rom[ 7988]='h00000b44;  wr_data_rom[ 7988]='h00000f7d;
    rd_cycle[ 7989] = 1'b1;  wr_cycle[ 7989] = 1'b0;  addr_rom[ 7989]='h000015d8;  wr_data_rom[ 7989]='h00000000;
    rd_cycle[ 7990] = 1'b0;  wr_cycle[ 7990] = 1'b1;  addr_rom[ 7990]='h000007e4;  wr_data_rom[ 7990]='h00000339;
    rd_cycle[ 7991] = 1'b1;  wr_cycle[ 7991] = 1'b0;  addr_rom[ 7991]='h00000bf0;  wr_data_rom[ 7991]='h00000000;
    rd_cycle[ 7992] = 1'b1;  wr_cycle[ 7992] = 1'b0;  addr_rom[ 7992]='h00000634;  wr_data_rom[ 7992]='h00000000;
    rd_cycle[ 7993] = 1'b1;  wr_cycle[ 7993] = 1'b0;  addr_rom[ 7993]='h000023a4;  wr_data_rom[ 7993]='h00000000;
    rd_cycle[ 7994] = 1'b1;  wr_cycle[ 7994] = 1'b0;  addr_rom[ 7994]='h0000357c;  wr_data_rom[ 7994]='h00000000;
    rd_cycle[ 7995] = 1'b0;  wr_cycle[ 7995] = 1'b1;  addr_rom[ 7995]='h0000030c;  wr_data_rom[ 7995]='h000002aa;
    rd_cycle[ 7996] = 1'b1;  wr_cycle[ 7996] = 1'b0;  addr_rom[ 7996]='h00003178;  wr_data_rom[ 7996]='h00000000;
    rd_cycle[ 7997] = 1'b0;  wr_cycle[ 7997] = 1'b1;  addr_rom[ 7997]='h0000239c;  wr_data_rom[ 7997]='h0000030d;
    rd_cycle[ 7998] = 1'b0;  wr_cycle[ 7998] = 1'b1;  addr_rom[ 7998]='h000033a0;  wr_data_rom[ 7998]='h00001f1a;
    rd_cycle[ 7999] = 1'b0;  wr_cycle[ 7999] = 1'b1;  addr_rom[ 7999]='h000031b8;  wr_data_rom[ 7999]='h000005a5;
    rd_cycle[ 8000] = 1'b1;  wr_cycle[ 8000] = 1'b0;  addr_rom[ 8000]='h000031a4;  wr_data_rom[ 8000]='h00000000;
    rd_cycle[ 8001] = 1'b1;  wr_cycle[ 8001] = 1'b0;  addr_rom[ 8001]='h00001ae8;  wr_data_rom[ 8001]='h00000000;
    rd_cycle[ 8002] = 1'b1;  wr_cycle[ 8002] = 1'b0;  addr_rom[ 8002]='h00002e54;  wr_data_rom[ 8002]='h00000000;
    rd_cycle[ 8003] = 1'b0;  wr_cycle[ 8003] = 1'b1;  addr_rom[ 8003]='h00002228;  wr_data_rom[ 8003]='h00000b3a;
    rd_cycle[ 8004] = 1'b0;  wr_cycle[ 8004] = 1'b1;  addr_rom[ 8004]='h000034a0;  wr_data_rom[ 8004]='h00001f15;
    rd_cycle[ 8005] = 1'b1;  wr_cycle[ 8005] = 1'b0;  addr_rom[ 8005]='h000012f8;  wr_data_rom[ 8005]='h00000000;
    rd_cycle[ 8006] = 1'b0;  wr_cycle[ 8006] = 1'b1;  addr_rom[ 8006]='h00001d48;  wr_data_rom[ 8006]='h00002d39;
    rd_cycle[ 8007] = 1'b0;  wr_cycle[ 8007] = 1'b1;  addr_rom[ 8007]='h000009cc;  wr_data_rom[ 8007]='h00001c9c;
    rd_cycle[ 8008] = 1'b0;  wr_cycle[ 8008] = 1'b1;  addr_rom[ 8008]='h000029a4;  wr_data_rom[ 8008]='h0000084b;
    rd_cycle[ 8009] = 1'b0;  wr_cycle[ 8009] = 1'b1;  addr_rom[ 8009]='h000037ac;  wr_data_rom[ 8009]='h000014d7;
    rd_cycle[ 8010] = 1'b1;  wr_cycle[ 8010] = 1'b0;  addr_rom[ 8010]='h00002004;  wr_data_rom[ 8010]='h00000000;
    rd_cycle[ 8011] = 1'b0;  wr_cycle[ 8011] = 1'b1;  addr_rom[ 8011]='h000000a8;  wr_data_rom[ 8011]='h00000ee8;
    rd_cycle[ 8012] = 1'b1;  wr_cycle[ 8012] = 1'b0;  addr_rom[ 8012]='h00003e8c;  wr_data_rom[ 8012]='h00000000;
    rd_cycle[ 8013] = 1'b1;  wr_cycle[ 8013] = 1'b0;  addr_rom[ 8013]='h0000386c;  wr_data_rom[ 8013]='h00000000;
    rd_cycle[ 8014] = 1'b1;  wr_cycle[ 8014] = 1'b0;  addr_rom[ 8014]='h00000be0;  wr_data_rom[ 8014]='h00000000;
    rd_cycle[ 8015] = 1'b0;  wr_cycle[ 8015] = 1'b1;  addr_rom[ 8015]='h00002474;  wr_data_rom[ 8015]='h0000173a;
    rd_cycle[ 8016] = 1'b1;  wr_cycle[ 8016] = 1'b0;  addr_rom[ 8016]='h000009e0;  wr_data_rom[ 8016]='h00000000;
    rd_cycle[ 8017] = 1'b1;  wr_cycle[ 8017] = 1'b0;  addr_rom[ 8017]='h00003b30;  wr_data_rom[ 8017]='h00000000;
    rd_cycle[ 8018] = 1'b1;  wr_cycle[ 8018] = 1'b0;  addr_rom[ 8018]='h00000b08;  wr_data_rom[ 8018]='h00000000;
    rd_cycle[ 8019] = 1'b0;  wr_cycle[ 8019] = 1'b1;  addr_rom[ 8019]='h000021e8;  wr_data_rom[ 8019]='h00002328;
    rd_cycle[ 8020] = 1'b0;  wr_cycle[ 8020] = 1'b1;  addr_rom[ 8020]='h00001590;  wr_data_rom[ 8020]='h0000315b;
    rd_cycle[ 8021] = 1'b0;  wr_cycle[ 8021] = 1'b1;  addr_rom[ 8021]='h00000fa8;  wr_data_rom[ 8021]='h00000d97;
    rd_cycle[ 8022] = 1'b1;  wr_cycle[ 8022] = 1'b0;  addr_rom[ 8022]='h0000094c;  wr_data_rom[ 8022]='h00000000;
    rd_cycle[ 8023] = 1'b0;  wr_cycle[ 8023] = 1'b1;  addr_rom[ 8023]='h00000850;  wr_data_rom[ 8023]='h00002336;
    rd_cycle[ 8024] = 1'b1;  wr_cycle[ 8024] = 1'b0;  addr_rom[ 8024]='h000030b4;  wr_data_rom[ 8024]='h00000000;
    rd_cycle[ 8025] = 1'b0;  wr_cycle[ 8025] = 1'b1;  addr_rom[ 8025]='h00001410;  wr_data_rom[ 8025]='h00001e89;
    rd_cycle[ 8026] = 1'b1;  wr_cycle[ 8026] = 1'b0;  addr_rom[ 8026]='h00001298;  wr_data_rom[ 8026]='h00000000;
    rd_cycle[ 8027] = 1'b0;  wr_cycle[ 8027] = 1'b1;  addr_rom[ 8027]='h000019f0;  wr_data_rom[ 8027]='h0000338e;
    rd_cycle[ 8028] = 1'b0;  wr_cycle[ 8028] = 1'b1;  addr_rom[ 8028]='h00003d7c;  wr_data_rom[ 8028]='h00000599;
    rd_cycle[ 8029] = 1'b1;  wr_cycle[ 8029] = 1'b0;  addr_rom[ 8029]='h00002bf4;  wr_data_rom[ 8029]='h00000000;
    rd_cycle[ 8030] = 1'b1;  wr_cycle[ 8030] = 1'b0;  addr_rom[ 8030]='h0000002c;  wr_data_rom[ 8030]='h00000000;
    rd_cycle[ 8031] = 1'b0;  wr_cycle[ 8031] = 1'b1;  addr_rom[ 8031]='h000030a4;  wr_data_rom[ 8031]='h00000b27;
    rd_cycle[ 8032] = 1'b0;  wr_cycle[ 8032] = 1'b1;  addr_rom[ 8032]='h00000df0;  wr_data_rom[ 8032]='h000014d7;
    rd_cycle[ 8033] = 1'b0;  wr_cycle[ 8033] = 1'b1;  addr_rom[ 8033]='h00003580;  wr_data_rom[ 8033]='h0000199c;
    rd_cycle[ 8034] = 1'b0;  wr_cycle[ 8034] = 1'b1;  addr_rom[ 8034]='h00002390;  wr_data_rom[ 8034]='h000034aa;
    rd_cycle[ 8035] = 1'b1;  wr_cycle[ 8035] = 1'b0;  addr_rom[ 8035]='h000032b0;  wr_data_rom[ 8035]='h00000000;
    rd_cycle[ 8036] = 1'b0;  wr_cycle[ 8036] = 1'b1;  addr_rom[ 8036]='h00000604;  wr_data_rom[ 8036]='h0000177d;
    rd_cycle[ 8037] = 1'b1;  wr_cycle[ 8037] = 1'b0;  addr_rom[ 8037]='h000038f8;  wr_data_rom[ 8037]='h00000000;
    rd_cycle[ 8038] = 1'b0;  wr_cycle[ 8038] = 1'b1;  addr_rom[ 8038]='h00001158;  wr_data_rom[ 8038]='h0000280a;
    rd_cycle[ 8039] = 1'b1;  wr_cycle[ 8039] = 1'b0;  addr_rom[ 8039]='h0000109c;  wr_data_rom[ 8039]='h00000000;
    rd_cycle[ 8040] = 1'b1;  wr_cycle[ 8040] = 1'b0;  addr_rom[ 8040]='h000015a4;  wr_data_rom[ 8040]='h00000000;
    rd_cycle[ 8041] = 1'b1;  wr_cycle[ 8041] = 1'b0;  addr_rom[ 8041]='h00001cd4;  wr_data_rom[ 8041]='h00000000;
    rd_cycle[ 8042] = 1'b1;  wr_cycle[ 8042] = 1'b0;  addr_rom[ 8042]='h00003978;  wr_data_rom[ 8042]='h00000000;
    rd_cycle[ 8043] = 1'b0;  wr_cycle[ 8043] = 1'b1;  addr_rom[ 8043]='h0000369c;  wr_data_rom[ 8043]='h000025e9;
    rd_cycle[ 8044] = 1'b0;  wr_cycle[ 8044] = 1'b1;  addr_rom[ 8044]='h00001514;  wr_data_rom[ 8044]='h00002062;
    rd_cycle[ 8045] = 1'b0;  wr_cycle[ 8045] = 1'b1;  addr_rom[ 8045]='h00000544;  wr_data_rom[ 8045]='h00000d69;
    rd_cycle[ 8046] = 1'b0;  wr_cycle[ 8046] = 1'b1;  addr_rom[ 8046]='h000034a8;  wr_data_rom[ 8046]='h00003cdb;
    rd_cycle[ 8047] = 1'b1;  wr_cycle[ 8047] = 1'b0;  addr_rom[ 8047]='h00000e44;  wr_data_rom[ 8047]='h00000000;
    rd_cycle[ 8048] = 1'b1;  wr_cycle[ 8048] = 1'b0;  addr_rom[ 8048]='h000008e0;  wr_data_rom[ 8048]='h00000000;
    rd_cycle[ 8049] = 1'b0;  wr_cycle[ 8049] = 1'b1;  addr_rom[ 8049]='h00000c18;  wr_data_rom[ 8049]='h0000117e;
    rd_cycle[ 8050] = 1'b1;  wr_cycle[ 8050] = 1'b0;  addr_rom[ 8050]='h000036a4;  wr_data_rom[ 8050]='h00000000;
    rd_cycle[ 8051] = 1'b1;  wr_cycle[ 8051] = 1'b0;  addr_rom[ 8051]='h00002c34;  wr_data_rom[ 8051]='h00000000;
    rd_cycle[ 8052] = 1'b1;  wr_cycle[ 8052] = 1'b0;  addr_rom[ 8052]='h00003c48;  wr_data_rom[ 8052]='h00000000;
    rd_cycle[ 8053] = 1'b0;  wr_cycle[ 8053] = 1'b1;  addr_rom[ 8053]='h00001784;  wr_data_rom[ 8053]='h00002cb0;
    rd_cycle[ 8054] = 1'b0;  wr_cycle[ 8054] = 1'b1;  addr_rom[ 8054]='h00003940;  wr_data_rom[ 8054]='h000013e8;
    rd_cycle[ 8055] = 1'b1;  wr_cycle[ 8055] = 1'b0;  addr_rom[ 8055]='h0000306c;  wr_data_rom[ 8055]='h00000000;
    rd_cycle[ 8056] = 1'b1;  wr_cycle[ 8056] = 1'b0;  addr_rom[ 8056]='h00000258;  wr_data_rom[ 8056]='h00000000;
    rd_cycle[ 8057] = 1'b1;  wr_cycle[ 8057] = 1'b0;  addr_rom[ 8057]='h00002fcc;  wr_data_rom[ 8057]='h00000000;
    rd_cycle[ 8058] = 1'b0;  wr_cycle[ 8058] = 1'b1;  addr_rom[ 8058]='h00001d8c;  wr_data_rom[ 8058]='h000039c3;
    rd_cycle[ 8059] = 1'b1;  wr_cycle[ 8059] = 1'b0;  addr_rom[ 8059]='h00000288;  wr_data_rom[ 8059]='h00000000;
    rd_cycle[ 8060] = 1'b0;  wr_cycle[ 8060] = 1'b1;  addr_rom[ 8060]='h00001154;  wr_data_rom[ 8060]='h000003fb;
    rd_cycle[ 8061] = 1'b0;  wr_cycle[ 8061] = 1'b1;  addr_rom[ 8061]='h00002418;  wr_data_rom[ 8061]='h0000121b;
    rd_cycle[ 8062] = 1'b0;  wr_cycle[ 8062] = 1'b1;  addr_rom[ 8062]='h00001d4c;  wr_data_rom[ 8062]='h00001302;
    rd_cycle[ 8063] = 1'b1;  wr_cycle[ 8063] = 1'b0;  addr_rom[ 8063]='h00001e74;  wr_data_rom[ 8063]='h00000000;
    rd_cycle[ 8064] = 1'b0;  wr_cycle[ 8064] = 1'b1;  addr_rom[ 8064]='h0000025c;  wr_data_rom[ 8064]='h00003efa;
    rd_cycle[ 8065] = 1'b0;  wr_cycle[ 8065] = 1'b1;  addr_rom[ 8065]='h00001718;  wr_data_rom[ 8065]='h00002dd1;
    rd_cycle[ 8066] = 1'b1;  wr_cycle[ 8066] = 1'b0;  addr_rom[ 8066]='h0000024c;  wr_data_rom[ 8066]='h00000000;
    rd_cycle[ 8067] = 1'b0;  wr_cycle[ 8067] = 1'b1;  addr_rom[ 8067]='h0000140c;  wr_data_rom[ 8067]='h000009d2;
    rd_cycle[ 8068] = 1'b1;  wr_cycle[ 8068] = 1'b0;  addr_rom[ 8068]='h00002f74;  wr_data_rom[ 8068]='h00000000;
    rd_cycle[ 8069] = 1'b0;  wr_cycle[ 8069] = 1'b1;  addr_rom[ 8069]='h00002054;  wr_data_rom[ 8069]='h00001c3f;
    rd_cycle[ 8070] = 1'b1;  wr_cycle[ 8070] = 1'b0;  addr_rom[ 8070]='h00001524;  wr_data_rom[ 8070]='h00000000;
    rd_cycle[ 8071] = 1'b1;  wr_cycle[ 8071] = 1'b0;  addr_rom[ 8071]='h00002788;  wr_data_rom[ 8071]='h00000000;
    rd_cycle[ 8072] = 1'b1;  wr_cycle[ 8072] = 1'b0;  addr_rom[ 8072]='h000030e0;  wr_data_rom[ 8072]='h00000000;
    rd_cycle[ 8073] = 1'b0;  wr_cycle[ 8073] = 1'b1;  addr_rom[ 8073]='h0000304c;  wr_data_rom[ 8073]='h00000f9b;
    rd_cycle[ 8074] = 1'b1;  wr_cycle[ 8074] = 1'b0;  addr_rom[ 8074]='h00002e10;  wr_data_rom[ 8074]='h00000000;
    rd_cycle[ 8075] = 1'b1;  wr_cycle[ 8075] = 1'b0;  addr_rom[ 8075]='h00000f74;  wr_data_rom[ 8075]='h00000000;
    rd_cycle[ 8076] = 1'b0;  wr_cycle[ 8076] = 1'b1;  addr_rom[ 8076]='h0000073c;  wr_data_rom[ 8076]='h00000a53;
    rd_cycle[ 8077] = 1'b0;  wr_cycle[ 8077] = 1'b1;  addr_rom[ 8077]='h00002a9c;  wr_data_rom[ 8077]='h00002188;
    rd_cycle[ 8078] = 1'b1;  wr_cycle[ 8078] = 1'b0;  addr_rom[ 8078]='h000025c4;  wr_data_rom[ 8078]='h00000000;
    rd_cycle[ 8079] = 1'b0;  wr_cycle[ 8079] = 1'b1;  addr_rom[ 8079]='h0000018c;  wr_data_rom[ 8079]='h00000281;
    rd_cycle[ 8080] = 1'b0;  wr_cycle[ 8080] = 1'b1;  addr_rom[ 8080]='h000032fc;  wr_data_rom[ 8080]='h0000256b;
    rd_cycle[ 8081] = 1'b0;  wr_cycle[ 8081] = 1'b1;  addr_rom[ 8081]='h00003d6c;  wr_data_rom[ 8081]='h0000172d;
    rd_cycle[ 8082] = 1'b0;  wr_cycle[ 8082] = 1'b1;  addr_rom[ 8082]='h00001ae8;  wr_data_rom[ 8082]='h000002cd;
    rd_cycle[ 8083] = 1'b0;  wr_cycle[ 8083] = 1'b1;  addr_rom[ 8083]='h00001998;  wr_data_rom[ 8083]='h00000422;
    rd_cycle[ 8084] = 1'b1;  wr_cycle[ 8084] = 1'b0;  addr_rom[ 8084]='h00000810;  wr_data_rom[ 8084]='h00000000;
    rd_cycle[ 8085] = 1'b1;  wr_cycle[ 8085] = 1'b0;  addr_rom[ 8085]='h00001b78;  wr_data_rom[ 8085]='h00000000;
    rd_cycle[ 8086] = 1'b1;  wr_cycle[ 8086] = 1'b0;  addr_rom[ 8086]='h000015a4;  wr_data_rom[ 8086]='h00000000;
    rd_cycle[ 8087] = 1'b0;  wr_cycle[ 8087] = 1'b1;  addr_rom[ 8087]='h00001b80;  wr_data_rom[ 8087]='h0000080b;
    rd_cycle[ 8088] = 1'b0;  wr_cycle[ 8088] = 1'b1;  addr_rom[ 8088]='h000033b4;  wr_data_rom[ 8088]='h00000ed3;
    rd_cycle[ 8089] = 1'b0;  wr_cycle[ 8089] = 1'b1;  addr_rom[ 8089]='h00002264;  wr_data_rom[ 8089]='h000007da;
    rd_cycle[ 8090] = 1'b0;  wr_cycle[ 8090] = 1'b1;  addr_rom[ 8090]='h0000349c;  wr_data_rom[ 8090]='h00003c16;
    rd_cycle[ 8091] = 1'b1;  wr_cycle[ 8091] = 1'b0;  addr_rom[ 8091]='h0000217c;  wr_data_rom[ 8091]='h00000000;
    rd_cycle[ 8092] = 1'b1;  wr_cycle[ 8092] = 1'b0;  addr_rom[ 8092]='h00002aa0;  wr_data_rom[ 8092]='h00000000;
    rd_cycle[ 8093] = 1'b1;  wr_cycle[ 8093] = 1'b0;  addr_rom[ 8093]='h00000d2c;  wr_data_rom[ 8093]='h00000000;
    rd_cycle[ 8094] = 1'b0;  wr_cycle[ 8094] = 1'b1;  addr_rom[ 8094]='h000021cc;  wr_data_rom[ 8094]='h00002dd2;
    rd_cycle[ 8095] = 1'b0;  wr_cycle[ 8095] = 1'b1;  addr_rom[ 8095]='h00001be8;  wr_data_rom[ 8095]='h00002504;
    rd_cycle[ 8096] = 1'b1;  wr_cycle[ 8096] = 1'b0;  addr_rom[ 8096]='h00001ab8;  wr_data_rom[ 8096]='h00000000;
    rd_cycle[ 8097] = 1'b1;  wr_cycle[ 8097] = 1'b0;  addr_rom[ 8097]='h000008a8;  wr_data_rom[ 8097]='h00000000;
    rd_cycle[ 8098] = 1'b0;  wr_cycle[ 8098] = 1'b1;  addr_rom[ 8098]='h00002770;  wr_data_rom[ 8098]='h0000039c;
    rd_cycle[ 8099] = 1'b1;  wr_cycle[ 8099] = 1'b0;  addr_rom[ 8099]='h000016e4;  wr_data_rom[ 8099]='h00000000;
    rd_cycle[ 8100] = 1'b1;  wr_cycle[ 8100] = 1'b0;  addr_rom[ 8100]='h00000c20;  wr_data_rom[ 8100]='h00000000;
    rd_cycle[ 8101] = 1'b0;  wr_cycle[ 8101] = 1'b1;  addr_rom[ 8101]='h00003e80;  wr_data_rom[ 8101]='h0000145a;
    rd_cycle[ 8102] = 1'b0;  wr_cycle[ 8102] = 1'b1;  addr_rom[ 8102]='h00000a2c;  wr_data_rom[ 8102]='h00002809;
    rd_cycle[ 8103] = 1'b1;  wr_cycle[ 8103] = 1'b0;  addr_rom[ 8103]='h00002944;  wr_data_rom[ 8103]='h00000000;
    rd_cycle[ 8104] = 1'b0;  wr_cycle[ 8104] = 1'b1;  addr_rom[ 8104]='h00001f28;  wr_data_rom[ 8104]='h000039d7;
    rd_cycle[ 8105] = 1'b0;  wr_cycle[ 8105] = 1'b1;  addr_rom[ 8105]='h000013e4;  wr_data_rom[ 8105]='h00003a36;
    rd_cycle[ 8106] = 1'b1;  wr_cycle[ 8106] = 1'b0;  addr_rom[ 8106]='h0000010c;  wr_data_rom[ 8106]='h00000000;
    rd_cycle[ 8107] = 1'b1;  wr_cycle[ 8107] = 1'b0;  addr_rom[ 8107]='h00001fc8;  wr_data_rom[ 8107]='h00000000;
    rd_cycle[ 8108] = 1'b1;  wr_cycle[ 8108] = 1'b0;  addr_rom[ 8108]='h000037e4;  wr_data_rom[ 8108]='h00000000;
    rd_cycle[ 8109] = 1'b0;  wr_cycle[ 8109] = 1'b1;  addr_rom[ 8109]='h000031f8;  wr_data_rom[ 8109]='h000039ca;
    rd_cycle[ 8110] = 1'b0;  wr_cycle[ 8110] = 1'b1;  addr_rom[ 8110]='h00002510;  wr_data_rom[ 8110]='h00000ff4;
    rd_cycle[ 8111] = 1'b0;  wr_cycle[ 8111] = 1'b1;  addr_rom[ 8111]='h00002b98;  wr_data_rom[ 8111]='h0000100e;
    rd_cycle[ 8112] = 1'b0;  wr_cycle[ 8112] = 1'b1;  addr_rom[ 8112]='h00001908;  wr_data_rom[ 8112]='h000010b9;
    rd_cycle[ 8113] = 1'b1;  wr_cycle[ 8113] = 1'b0;  addr_rom[ 8113]='h00002650;  wr_data_rom[ 8113]='h00000000;
    rd_cycle[ 8114] = 1'b0;  wr_cycle[ 8114] = 1'b1;  addr_rom[ 8114]='h00000d34;  wr_data_rom[ 8114]='h000006fe;
    rd_cycle[ 8115] = 1'b0;  wr_cycle[ 8115] = 1'b1;  addr_rom[ 8115]='h00002f98;  wr_data_rom[ 8115]='h000027e7;
    rd_cycle[ 8116] = 1'b0;  wr_cycle[ 8116] = 1'b1;  addr_rom[ 8116]='h000007d4;  wr_data_rom[ 8116]='h000036a2;
    rd_cycle[ 8117] = 1'b1;  wr_cycle[ 8117] = 1'b0;  addr_rom[ 8117]='h0000310c;  wr_data_rom[ 8117]='h00000000;
    rd_cycle[ 8118] = 1'b0;  wr_cycle[ 8118] = 1'b1;  addr_rom[ 8118]='h000006e4;  wr_data_rom[ 8118]='h0000197d;
    rd_cycle[ 8119] = 1'b1;  wr_cycle[ 8119] = 1'b0;  addr_rom[ 8119]='h00000e8c;  wr_data_rom[ 8119]='h00000000;
    rd_cycle[ 8120] = 1'b0;  wr_cycle[ 8120] = 1'b1;  addr_rom[ 8120]='h000000f0;  wr_data_rom[ 8120]='h00000781;
    rd_cycle[ 8121] = 1'b1;  wr_cycle[ 8121] = 1'b0;  addr_rom[ 8121]='h00003384;  wr_data_rom[ 8121]='h00000000;
    rd_cycle[ 8122] = 1'b1;  wr_cycle[ 8122] = 1'b0;  addr_rom[ 8122]='h00002660;  wr_data_rom[ 8122]='h00000000;
    rd_cycle[ 8123] = 1'b0;  wr_cycle[ 8123] = 1'b1;  addr_rom[ 8123]='h00002fc8;  wr_data_rom[ 8123]='h00000f19;
    rd_cycle[ 8124] = 1'b0;  wr_cycle[ 8124] = 1'b1;  addr_rom[ 8124]='h00001a38;  wr_data_rom[ 8124]='h00003407;
    rd_cycle[ 8125] = 1'b1;  wr_cycle[ 8125] = 1'b0;  addr_rom[ 8125]='h00003a44;  wr_data_rom[ 8125]='h00000000;
    rd_cycle[ 8126] = 1'b1;  wr_cycle[ 8126] = 1'b0;  addr_rom[ 8126]='h00000850;  wr_data_rom[ 8126]='h00000000;
    rd_cycle[ 8127] = 1'b1;  wr_cycle[ 8127] = 1'b0;  addr_rom[ 8127]='h00003cf4;  wr_data_rom[ 8127]='h00000000;
    rd_cycle[ 8128] = 1'b1;  wr_cycle[ 8128] = 1'b0;  addr_rom[ 8128]='h000018d8;  wr_data_rom[ 8128]='h00000000;
    rd_cycle[ 8129] = 1'b1;  wr_cycle[ 8129] = 1'b0;  addr_rom[ 8129]='h000026d4;  wr_data_rom[ 8129]='h00000000;
    rd_cycle[ 8130] = 1'b0;  wr_cycle[ 8130] = 1'b1;  addr_rom[ 8130]='h00001bcc;  wr_data_rom[ 8130]='h00001fbf;
    rd_cycle[ 8131] = 1'b0;  wr_cycle[ 8131] = 1'b1;  addr_rom[ 8131]='h000029c0;  wr_data_rom[ 8131]='h00000648;
    rd_cycle[ 8132] = 1'b1;  wr_cycle[ 8132] = 1'b0;  addr_rom[ 8132]='h00003a00;  wr_data_rom[ 8132]='h00000000;
    rd_cycle[ 8133] = 1'b0;  wr_cycle[ 8133] = 1'b1;  addr_rom[ 8133]='h00001b4c;  wr_data_rom[ 8133]='h00003632;
    rd_cycle[ 8134] = 1'b1;  wr_cycle[ 8134] = 1'b0;  addr_rom[ 8134]='h000038a8;  wr_data_rom[ 8134]='h00000000;
    rd_cycle[ 8135] = 1'b0;  wr_cycle[ 8135] = 1'b1;  addr_rom[ 8135]='h00001cfc;  wr_data_rom[ 8135]='h00002ff2;
    rd_cycle[ 8136] = 1'b0;  wr_cycle[ 8136] = 1'b1;  addr_rom[ 8136]='h00003018;  wr_data_rom[ 8136]='h00000e6d;
    rd_cycle[ 8137] = 1'b0;  wr_cycle[ 8137] = 1'b1;  addr_rom[ 8137]='h000017b8;  wr_data_rom[ 8137]='h00003d6e;
    rd_cycle[ 8138] = 1'b1;  wr_cycle[ 8138] = 1'b0;  addr_rom[ 8138]='h00000b2c;  wr_data_rom[ 8138]='h00000000;
    rd_cycle[ 8139] = 1'b0;  wr_cycle[ 8139] = 1'b1;  addr_rom[ 8139]='h00002ce0;  wr_data_rom[ 8139]='h00000476;
    rd_cycle[ 8140] = 1'b0;  wr_cycle[ 8140] = 1'b1;  addr_rom[ 8140]='h00002418;  wr_data_rom[ 8140]='h00002991;
    rd_cycle[ 8141] = 1'b1;  wr_cycle[ 8141] = 1'b0;  addr_rom[ 8141]='h00001f94;  wr_data_rom[ 8141]='h00000000;
    rd_cycle[ 8142] = 1'b0;  wr_cycle[ 8142] = 1'b1;  addr_rom[ 8142]='h00000b7c;  wr_data_rom[ 8142]='h00003c1c;
    rd_cycle[ 8143] = 1'b0;  wr_cycle[ 8143] = 1'b1;  addr_rom[ 8143]='h00002ef4;  wr_data_rom[ 8143]='h000004ba;
    rd_cycle[ 8144] = 1'b1;  wr_cycle[ 8144] = 1'b0;  addr_rom[ 8144]='h000013d4;  wr_data_rom[ 8144]='h00000000;
    rd_cycle[ 8145] = 1'b1;  wr_cycle[ 8145] = 1'b0;  addr_rom[ 8145]='h0000198c;  wr_data_rom[ 8145]='h00000000;
    rd_cycle[ 8146] = 1'b0;  wr_cycle[ 8146] = 1'b1;  addr_rom[ 8146]='h00000be0;  wr_data_rom[ 8146]='h00002f26;
    rd_cycle[ 8147] = 1'b0;  wr_cycle[ 8147] = 1'b1;  addr_rom[ 8147]='h000033ac;  wr_data_rom[ 8147]='h00001914;
    rd_cycle[ 8148] = 1'b1;  wr_cycle[ 8148] = 1'b0;  addr_rom[ 8148]='h000024b8;  wr_data_rom[ 8148]='h00000000;
    rd_cycle[ 8149] = 1'b0;  wr_cycle[ 8149] = 1'b1;  addr_rom[ 8149]='h00003860;  wr_data_rom[ 8149]='h000010d2;
    rd_cycle[ 8150] = 1'b1;  wr_cycle[ 8150] = 1'b0;  addr_rom[ 8150]='h000005a4;  wr_data_rom[ 8150]='h00000000;
    rd_cycle[ 8151] = 1'b1;  wr_cycle[ 8151] = 1'b0;  addr_rom[ 8151]='h000008b0;  wr_data_rom[ 8151]='h00000000;
    rd_cycle[ 8152] = 1'b0;  wr_cycle[ 8152] = 1'b1;  addr_rom[ 8152]='h00001de0;  wr_data_rom[ 8152]='h00003f8a;
    rd_cycle[ 8153] = 1'b1;  wr_cycle[ 8153] = 1'b0;  addr_rom[ 8153]='h00003e70;  wr_data_rom[ 8153]='h00000000;
    rd_cycle[ 8154] = 1'b1;  wr_cycle[ 8154] = 1'b0;  addr_rom[ 8154]='h000009b0;  wr_data_rom[ 8154]='h00000000;
    rd_cycle[ 8155] = 1'b1;  wr_cycle[ 8155] = 1'b0;  addr_rom[ 8155]='h000039f0;  wr_data_rom[ 8155]='h00000000;
    rd_cycle[ 8156] = 1'b0;  wr_cycle[ 8156] = 1'b1;  addr_rom[ 8156]='h00002000;  wr_data_rom[ 8156]='h00001858;
    rd_cycle[ 8157] = 1'b0;  wr_cycle[ 8157] = 1'b1;  addr_rom[ 8157]='h00001208;  wr_data_rom[ 8157]='h00001f96;
    rd_cycle[ 8158] = 1'b1;  wr_cycle[ 8158] = 1'b0;  addr_rom[ 8158]='h000002d4;  wr_data_rom[ 8158]='h00000000;
    rd_cycle[ 8159] = 1'b1;  wr_cycle[ 8159] = 1'b0;  addr_rom[ 8159]='h00002390;  wr_data_rom[ 8159]='h00000000;
    rd_cycle[ 8160] = 1'b1;  wr_cycle[ 8160] = 1'b0;  addr_rom[ 8160]='h00000fd4;  wr_data_rom[ 8160]='h00000000;
    rd_cycle[ 8161] = 1'b1;  wr_cycle[ 8161] = 1'b0;  addr_rom[ 8161]='h000023ec;  wr_data_rom[ 8161]='h00000000;
    rd_cycle[ 8162] = 1'b0;  wr_cycle[ 8162] = 1'b1;  addr_rom[ 8162]='h000021d0;  wr_data_rom[ 8162]='h0000276a;
    rd_cycle[ 8163] = 1'b0;  wr_cycle[ 8163] = 1'b1;  addr_rom[ 8163]='h00002408;  wr_data_rom[ 8163]='h0000220a;
    rd_cycle[ 8164] = 1'b0;  wr_cycle[ 8164] = 1'b1;  addr_rom[ 8164]='h00000eb0;  wr_data_rom[ 8164]='h000022a3;
    rd_cycle[ 8165] = 1'b1;  wr_cycle[ 8165] = 1'b0;  addr_rom[ 8165]='h00003e84;  wr_data_rom[ 8165]='h00000000;
    rd_cycle[ 8166] = 1'b1;  wr_cycle[ 8166] = 1'b0;  addr_rom[ 8166]='h000005dc;  wr_data_rom[ 8166]='h00000000;
    rd_cycle[ 8167] = 1'b0;  wr_cycle[ 8167] = 1'b1;  addr_rom[ 8167]='h000000b0;  wr_data_rom[ 8167]='h00003434;
    rd_cycle[ 8168] = 1'b0;  wr_cycle[ 8168] = 1'b1;  addr_rom[ 8168]='h0000113c;  wr_data_rom[ 8168]='h00002b3f;
    rd_cycle[ 8169] = 1'b1;  wr_cycle[ 8169] = 1'b0;  addr_rom[ 8169]='h00000978;  wr_data_rom[ 8169]='h00000000;
    rd_cycle[ 8170] = 1'b0;  wr_cycle[ 8170] = 1'b1;  addr_rom[ 8170]='h00002e44;  wr_data_rom[ 8170]='h00003546;
    rd_cycle[ 8171] = 1'b1;  wr_cycle[ 8171] = 1'b0;  addr_rom[ 8171]='h00000160;  wr_data_rom[ 8171]='h00000000;
    rd_cycle[ 8172] = 1'b0;  wr_cycle[ 8172] = 1'b1;  addr_rom[ 8172]='h00001e5c;  wr_data_rom[ 8172]='h00002c66;
    rd_cycle[ 8173] = 1'b0;  wr_cycle[ 8173] = 1'b1;  addr_rom[ 8173]='h00000854;  wr_data_rom[ 8173]='h00003383;
    rd_cycle[ 8174] = 1'b1;  wr_cycle[ 8174] = 1'b0;  addr_rom[ 8174]='h00001a30;  wr_data_rom[ 8174]='h00000000;
    rd_cycle[ 8175] = 1'b1;  wr_cycle[ 8175] = 1'b0;  addr_rom[ 8175]='h000030b0;  wr_data_rom[ 8175]='h00000000;
    rd_cycle[ 8176] = 1'b1;  wr_cycle[ 8176] = 1'b0;  addr_rom[ 8176]='h000030bc;  wr_data_rom[ 8176]='h00000000;
    rd_cycle[ 8177] = 1'b0;  wr_cycle[ 8177] = 1'b1;  addr_rom[ 8177]='h00003044;  wr_data_rom[ 8177]='h00002a50;
    rd_cycle[ 8178] = 1'b1;  wr_cycle[ 8178] = 1'b0;  addr_rom[ 8178]='h000008f8;  wr_data_rom[ 8178]='h00000000;
    rd_cycle[ 8179] = 1'b0;  wr_cycle[ 8179] = 1'b1;  addr_rom[ 8179]='h00002a8c;  wr_data_rom[ 8179]='h000033af;
    rd_cycle[ 8180] = 1'b0;  wr_cycle[ 8180] = 1'b1;  addr_rom[ 8180]='h00000eb8;  wr_data_rom[ 8180]='h00003ec1;
    rd_cycle[ 8181] = 1'b0;  wr_cycle[ 8181] = 1'b1;  addr_rom[ 8181]='h0000076c;  wr_data_rom[ 8181]='h00001ea8;
    rd_cycle[ 8182] = 1'b0;  wr_cycle[ 8182] = 1'b1;  addr_rom[ 8182]='h00000a7c;  wr_data_rom[ 8182]='h00000117;
    rd_cycle[ 8183] = 1'b1;  wr_cycle[ 8183] = 1'b0;  addr_rom[ 8183]='h0000217c;  wr_data_rom[ 8183]='h00000000;
    rd_cycle[ 8184] = 1'b0;  wr_cycle[ 8184] = 1'b1;  addr_rom[ 8184]='h000025f0;  wr_data_rom[ 8184]='h0000324f;
    rd_cycle[ 8185] = 1'b0;  wr_cycle[ 8185] = 1'b1;  addr_rom[ 8185]='h00003418;  wr_data_rom[ 8185]='h00000799;
    rd_cycle[ 8186] = 1'b0;  wr_cycle[ 8186] = 1'b1;  addr_rom[ 8186]='h00000680;  wr_data_rom[ 8186]='h00001c47;
    rd_cycle[ 8187] = 1'b0;  wr_cycle[ 8187] = 1'b1;  addr_rom[ 8187]='h00002818;  wr_data_rom[ 8187]='h00000806;
    rd_cycle[ 8188] = 1'b1;  wr_cycle[ 8188] = 1'b0;  addr_rom[ 8188]='h0000058c;  wr_data_rom[ 8188]='h00000000;
    rd_cycle[ 8189] = 1'b0;  wr_cycle[ 8189] = 1'b1;  addr_rom[ 8189]='h000021e8;  wr_data_rom[ 8189]='h00003699;
    rd_cycle[ 8190] = 1'b0;  wr_cycle[ 8190] = 1'b1;  addr_rom[ 8190]='h0000118c;  wr_data_rom[ 8190]='h0000100a;
    rd_cycle[ 8191] = 1'b0;  wr_cycle[ 8191] = 1'b1;  addr_rom[ 8191]='h00000cb0;  wr_data_rom[ 8191]='h000000b6;
    rd_cycle[ 8192] = 1'b1;  wr_cycle[ 8192] = 1'b0;  addr_rom[ 8192]='h00001190;  wr_data_rom[ 8192]='h00000000;
    rd_cycle[ 8193] = 1'b1;  wr_cycle[ 8193] = 1'b0;  addr_rom[ 8193]='h000027e8;  wr_data_rom[ 8193]='h00000000;
    rd_cycle[ 8194] = 1'b1;  wr_cycle[ 8194] = 1'b0;  addr_rom[ 8194]='h000006ac;  wr_data_rom[ 8194]='h00000000;
    rd_cycle[ 8195] = 1'b1;  wr_cycle[ 8195] = 1'b0;  addr_rom[ 8195]='h00001910;  wr_data_rom[ 8195]='h00000000;
    rd_cycle[ 8196] = 1'b1;  wr_cycle[ 8196] = 1'b0;  addr_rom[ 8196]='h00000c40;  wr_data_rom[ 8196]='h00000000;
    rd_cycle[ 8197] = 1'b0;  wr_cycle[ 8197] = 1'b1;  addr_rom[ 8197]='h00002d00;  wr_data_rom[ 8197]='h00002488;
    rd_cycle[ 8198] = 1'b0;  wr_cycle[ 8198] = 1'b1;  addr_rom[ 8198]='h000005f0;  wr_data_rom[ 8198]='h00003f72;
    rd_cycle[ 8199] = 1'b0;  wr_cycle[ 8199] = 1'b1;  addr_rom[ 8199]='h000029a8;  wr_data_rom[ 8199]='h000000d4;
    rd_cycle[ 8200] = 1'b0;  wr_cycle[ 8200] = 1'b1;  addr_rom[ 8200]='h0000178c;  wr_data_rom[ 8200]='h000038d6;
    rd_cycle[ 8201] = 1'b0;  wr_cycle[ 8201] = 1'b1;  addr_rom[ 8201]='h00001e58;  wr_data_rom[ 8201]='h00003306;
    rd_cycle[ 8202] = 1'b0;  wr_cycle[ 8202] = 1'b1;  addr_rom[ 8202]='h00000220;  wr_data_rom[ 8202]='h000035f9;
    rd_cycle[ 8203] = 1'b1;  wr_cycle[ 8203] = 1'b0;  addr_rom[ 8203]='h00000478;  wr_data_rom[ 8203]='h00000000;
    rd_cycle[ 8204] = 1'b0;  wr_cycle[ 8204] = 1'b1;  addr_rom[ 8204]='h0000233c;  wr_data_rom[ 8204]='h000018ae;
    rd_cycle[ 8205] = 1'b1;  wr_cycle[ 8205] = 1'b0;  addr_rom[ 8205]='h0000249c;  wr_data_rom[ 8205]='h00000000;
    rd_cycle[ 8206] = 1'b0;  wr_cycle[ 8206] = 1'b1;  addr_rom[ 8206]='h0000391c;  wr_data_rom[ 8206]='h00002142;
    rd_cycle[ 8207] = 1'b1;  wr_cycle[ 8207] = 1'b0;  addr_rom[ 8207]='h00002920;  wr_data_rom[ 8207]='h00000000;
    rd_cycle[ 8208] = 1'b1;  wr_cycle[ 8208] = 1'b0;  addr_rom[ 8208]='h00000398;  wr_data_rom[ 8208]='h00000000;
    rd_cycle[ 8209] = 1'b0;  wr_cycle[ 8209] = 1'b1;  addr_rom[ 8209]='h00003328;  wr_data_rom[ 8209]='h00002a1e;
    rd_cycle[ 8210] = 1'b1;  wr_cycle[ 8210] = 1'b0;  addr_rom[ 8210]='h000027f8;  wr_data_rom[ 8210]='h00000000;
    rd_cycle[ 8211] = 1'b1;  wr_cycle[ 8211] = 1'b0;  addr_rom[ 8211]='h00002a70;  wr_data_rom[ 8211]='h00000000;
    rd_cycle[ 8212] = 1'b1;  wr_cycle[ 8212] = 1'b0;  addr_rom[ 8212]='h000003bc;  wr_data_rom[ 8212]='h00000000;
    rd_cycle[ 8213] = 1'b1;  wr_cycle[ 8213] = 1'b0;  addr_rom[ 8213]='h00000cf4;  wr_data_rom[ 8213]='h00000000;
    rd_cycle[ 8214] = 1'b1;  wr_cycle[ 8214] = 1'b0;  addr_rom[ 8214]='h000016a8;  wr_data_rom[ 8214]='h00000000;
    rd_cycle[ 8215] = 1'b0;  wr_cycle[ 8215] = 1'b1;  addr_rom[ 8215]='h000015b0;  wr_data_rom[ 8215]='h0000015f;
    rd_cycle[ 8216] = 1'b1;  wr_cycle[ 8216] = 1'b0;  addr_rom[ 8216]='h00003044;  wr_data_rom[ 8216]='h00000000;
    rd_cycle[ 8217] = 1'b0;  wr_cycle[ 8217] = 1'b1;  addr_rom[ 8217]='h000024bc;  wr_data_rom[ 8217]='h00000515;
    rd_cycle[ 8218] = 1'b0;  wr_cycle[ 8218] = 1'b1;  addr_rom[ 8218]='h00001cd0;  wr_data_rom[ 8218]='h000029c6;
    rd_cycle[ 8219] = 1'b1;  wr_cycle[ 8219] = 1'b0;  addr_rom[ 8219]='h00002b5c;  wr_data_rom[ 8219]='h00000000;
    rd_cycle[ 8220] = 1'b1;  wr_cycle[ 8220] = 1'b0;  addr_rom[ 8220]='h00000ab4;  wr_data_rom[ 8220]='h00000000;
    rd_cycle[ 8221] = 1'b0;  wr_cycle[ 8221] = 1'b1;  addr_rom[ 8221]='h00000864;  wr_data_rom[ 8221]='h00001b30;
    rd_cycle[ 8222] = 1'b0;  wr_cycle[ 8222] = 1'b1;  addr_rom[ 8222]='h00002300;  wr_data_rom[ 8222]='h00003bbc;
    rd_cycle[ 8223] = 1'b0;  wr_cycle[ 8223] = 1'b1;  addr_rom[ 8223]='h0000386c;  wr_data_rom[ 8223]='h00001786;
    rd_cycle[ 8224] = 1'b0;  wr_cycle[ 8224] = 1'b1;  addr_rom[ 8224]='h00000930;  wr_data_rom[ 8224]='h00003052;
    rd_cycle[ 8225] = 1'b0;  wr_cycle[ 8225] = 1'b1;  addr_rom[ 8225]='h00003c08;  wr_data_rom[ 8225]='h00001c3a;
    rd_cycle[ 8226] = 1'b1;  wr_cycle[ 8226] = 1'b0;  addr_rom[ 8226]='h0000179c;  wr_data_rom[ 8226]='h00000000;
    rd_cycle[ 8227] = 1'b1;  wr_cycle[ 8227] = 1'b0;  addr_rom[ 8227]='h00001380;  wr_data_rom[ 8227]='h00000000;
    rd_cycle[ 8228] = 1'b0;  wr_cycle[ 8228] = 1'b1;  addr_rom[ 8228]='h0000050c;  wr_data_rom[ 8228]='h0000092b;
    rd_cycle[ 8229] = 1'b0;  wr_cycle[ 8229] = 1'b1;  addr_rom[ 8229]='h0000253c;  wr_data_rom[ 8229]='h000011d2;
    rd_cycle[ 8230] = 1'b1;  wr_cycle[ 8230] = 1'b0;  addr_rom[ 8230]='h000006d0;  wr_data_rom[ 8230]='h00000000;
    rd_cycle[ 8231] = 1'b0;  wr_cycle[ 8231] = 1'b1;  addr_rom[ 8231]='h00002f18;  wr_data_rom[ 8231]='h00000891;
    rd_cycle[ 8232] = 1'b1;  wr_cycle[ 8232] = 1'b0;  addr_rom[ 8232]='h000034e0;  wr_data_rom[ 8232]='h00000000;
    rd_cycle[ 8233] = 1'b1;  wr_cycle[ 8233] = 1'b0;  addr_rom[ 8233]='h000003d0;  wr_data_rom[ 8233]='h00000000;
    rd_cycle[ 8234] = 1'b1;  wr_cycle[ 8234] = 1'b0;  addr_rom[ 8234]='h00002b24;  wr_data_rom[ 8234]='h00000000;
    rd_cycle[ 8235] = 1'b0;  wr_cycle[ 8235] = 1'b1;  addr_rom[ 8235]='h0000221c;  wr_data_rom[ 8235]='h00003a0a;
    rd_cycle[ 8236] = 1'b1;  wr_cycle[ 8236] = 1'b0;  addr_rom[ 8236]='h000023c4;  wr_data_rom[ 8236]='h00000000;
    rd_cycle[ 8237] = 1'b1;  wr_cycle[ 8237] = 1'b0;  addr_rom[ 8237]='h00001ee8;  wr_data_rom[ 8237]='h00000000;
    rd_cycle[ 8238] = 1'b1;  wr_cycle[ 8238] = 1'b0;  addr_rom[ 8238]='h00001514;  wr_data_rom[ 8238]='h00000000;
    rd_cycle[ 8239] = 1'b0;  wr_cycle[ 8239] = 1'b1;  addr_rom[ 8239]='h00001e1c;  wr_data_rom[ 8239]='h00003bd9;
    rd_cycle[ 8240] = 1'b1;  wr_cycle[ 8240] = 1'b0;  addr_rom[ 8240]='h00003274;  wr_data_rom[ 8240]='h00000000;
    rd_cycle[ 8241] = 1'b1;  wr_cycle[ 8241] = 1'b0;  addr_rom[ 8241]='h00003d5c;  wr_data_rom[ 8241]='h00000000;
    rd_cycle[ 8242] = 1'b0;  wr_cycle[ 8242] = 1'b1;  addr_rom[ 8242]='h00003518;  wr_data_rom[ 8242]='h000038b0;
    rd_cycle[ 8243] = 1'b1;  wr_cycle[ 8243] = 1'b0;  addr_rom[ 8243]='h00003dcc;  wr_data_rom[ 8243]='h00000000;
    rd_cycle[ 8244] = 1'b0;  wr_cycle[ 8244] = 1'b1;  addr_rom[ 8244]='h00003b7c;  wr_data_rom[ 8244]='h00003213;
    rd_cycle[ 8245] = 1'b1;  wr_cycle[ 8245] = 1'b0;  addr_rom[ 8245]='h00003bcc;  wr_data_rom[ 8245]='h00000000;
    rd_cycle[ 8246] = 1'b0;  wr_cycle[ 8246] = 1'b1;  addr_rom[ 8246]='h0000344c;  wr_data_rom[ 8246]='h00002751;
    rd_cycle[ 8247] = 1'b1;  wr_cycle[ 8247] = 1'b0;  addr_rom[ 8247]='h000012d8;  wr_data_rom[ 8247]='h00000000;
    rd_cycle[ 8248] = 1'b0;  wr_cycle[ 8248] = 1'b1;  addr_rom[ 8248]='h00002058;  wr_data_rom[ 8248]='h00000623;
    rd_cycle[ 8249] = 1'b0;  wr_cycle[ 8249] = 1'b1;  addr_rom[ 8249]='h0000182c;  wr_data_rom[ 8249]='h00003de8;
    rd_cycle[ 8250] = 1'b1;  wr_cycle[ 8250] = 1'b0;  addr_rom[ 8250]='h000013dc;  wr_data_rom[ 8250]='h00000000;
    rd_cycle[ 8251] = 1'b0;  wr_cycle[ 8251] = 1'b1;  addr_rom[ 8251]='h000005d8;  wr_data_rom[ 8251]='h00003bd6;
    rd_cycle[ 8252] = 1'b1;  wr_cycle[ 8252] = 1'b0;  addr_rom[ 8252]='h00001f40;  wr_data_rom[ 8252]='h00000000;
    rd_cycle[ 8253] = 1'b1;  wr_cycle[ 8253] = 1'b0;  addr_rom[ 8253]='h000032ac;  wr_data_rom[ 8253]='h00000000;
    rd_cycle[ 8254] = 1'b0;  wr_cycle[ 8254] = 1'b1;  addr_rom[ 8254]='h00001858;  wr_data_rom[ 8254]='h0000106a;
    rd_cycle[ 8255] = 1'b0;  wr_cycle[ 8255] = 1'b1;  addr_rom[ 8255]='h0000273c;  wr_data_rom[ 8255]='h00002d5a;
    rd_cycle[ 8256] = 1'b1;  wr_cycle[ 8256] = 1'b0;  addr_rom[ 8256]='h00002b84;  wr_data_rom[ 8256]='h00000000;
    rd_cycle[ 8257] = 1'b0;  wr_cycle[ 8257] = 1'b1;  addr_rom[ 8257]='h0000028c;  wr_data_rom[ 8257]='h00001855;
    rd_cycle[ 8258] = 1'b0;  wr_cycle[ 8258] = 1'b1;  addr_rom[ 8258]='h00001aa8;  wr_data_rom[ 8258]='h00002878;
    rd_cycle[ 8259] = 1'b1;  wr_cycle[ 8259] = 1'b0;  addr_rom[ 8259]='h000037b8;  wr_data_rom[ 8259]='h00000000;
    rd_cycle[ 8260] = 1'b0;  wr_cycle[ 8260] = 1'b1;  addr_rom[ 8260]='h000013f0;  wr_data_rom[ 8260]='h0000082b;
    rd_cycle[ 8261] = 1'b1;  wr_cycle[ 8261] = 1'b0;  addr_rom[ 8261]='h00003c28;  wr_data_rom[ 8261]='h00000000;
    rd_cycle[ 8262] = 1'b0;  wr_cycle[ 8262] = 1'b1;  addr_rom[ 8262]='h0000059c;  wr_data_rom[ 8262]='h00002562;
    rd_cycle[ 8263] = 1'b0;  wr_cycle[ 8263] = 1'b1;  addr_rom[ 8263]='h00002ef4;  wr_data_rom[ 8263]='h000013cf;
    rd_cycle[ 8264] = 1'b0;  wr_cycle[ 8264] = 1'b1;  addr_rom[ 8264]='h00001058;  wr_data_rom[ 8264]='h00002a5a;
    rd_cycle[ 8265] = 1'b0;  wr_cycle[ 8265] = 1'b1;  addr_rom[ 8265]='h00001aa0;  wr_data_rom[ 8265]='h00003227;
    rd_cycle[ 8266] = 1'b1;  wr_cycle[ 8266] = 1'b0;  addr_rom[ 8266]='h00003d84;  wr_data_rom[ 8266]='h00000000;
    rd_cycle[ 8267] = 1'b0;  wr_cycle[ 8267] = 1'b1;  addr_rom[ 8267]='h00001c24;  wr_data_rom[ 8267]='h00003455;
    rd_cycle[ 8268] = 1'b1;  wr_cycle[ 8268] = 1'b0;  addr_rom[ 8268]='h00003be0;  wr_data_rom[ 8268]='h00000000;
    rd_cycle[ 8269] = 1'b1;  wr_cycle[ 8269] = 1'b0;  addr_rom[ 8269]='h00001ec4;  wr_data_rom[ 8269]='h00000000;
    rd_cycle[ 8270] = 1'b0;  wr_cycle[ 8270] = 1'b1;  addr_rom[ 8270]='h00000238;  wr_data_rom[ 8270]='h00003bdb;
    rd_cycle[ 8271] = 1'b1;  wr_cycle[ 8271] = 1'b0;  addr_rom[ 8271]='h00002ee4;  wr_data_rom[ 8271]='h00000000;
    rd_cycle[ 8272] = 1'b1;  wr_cycle[ 8272] = 1'b0;  addr_rom[ 8272]='h000002b8;  wr_data_rom[ 8272]='h00000000;
    rd_cycle[ 8273] = 1'b0;  wr_cycle[ 8273] = 1'b1;  addr_rom[ 8273]='h00002604;  wr_data_rom[ 8273]='h00001e6f;
    rd_cycle[ 8274] = 1'b0;  wr_cycle[ 8274] = 1'b1;  addr_rom[ 8274]='h00001d18;  wr_data_rom[ 8274]='h00002df1;
    rd_cycle[ 8275] = 1'b0;  wr_cycle[ 8275] = 1'b1;  addr_rom[ 8275]='h000004dc;  wr_data_rom[ 8275]='h00002e86;
    rd_cycle[ 8276] = 1'b0;  wr_cycle[ 8276] = 1'b1;  addr_rom[ 8276]='h00001588;  wr_data_rom[ 8276]='h0000168a;
    rd_cycle[ 8277] = 1'b1;  wr_cycle[ 8277] = 1'b0;  addr_rom[ 8277]='h00001344;  wr_data_rom[ 8277]='h00000000;
    rd_cycle[ 8278] = 1'b0;  wr_cycle[ 8278] = 1'b1;  addr_rom[ 8278]='h0000164c;  wr_data_rom[ 8278]='h000014c9;
    rd_cycle[ 8279] = 1'b0;  wr_cycle[ 8279] = 1'b1;  addr_rom[ 8279]='h00002cac;  wr_data_rom[ 8279]='h00002478;
    rd_cycle[ 8280] = 1'b0;  wr_cycle[ 8280] = 1'b1;  addr_rom[ 8280]='h000004d4;  wr_data_rom[ 8280]='h000035cf;
    rd_cycle[ 8281] = 1'b0;  wr_cycle[ 8281] = 1'b1;  addr_rom[ 8281]='h00002384;  wr_data_rom[ 8281]='h00000991;
    rd_cycle[ 8282] = 1'b1;  wr_cycle[ 8282] = 1'b0;  addr_rom[ 8282]='h00000268;  wr_data_rom[ 8282]='h00000000;
    rd_cycle[ 8283] = 1'b0;  wr_cycle[ 8283] = 1'b1;  addr_rom[ 8283]='h00002810;  wr_data_rom[ 8283]='h00003384;
    rd_cycle[ 8284] = 1'b0;  wr_cycle[ 8284] = 1'b1;  addr_rom[ 8284]='h00003a70;  wr_data_rom[ 8284]='h000033d8;
    rd_cycle[ 8285] = 1'b0;  wr_cycle[ 8285] = 1'b1;  addr_rom[ 8285]='h00000328;  wr_data_rom[ 8285]='h000017c2;
    rd_cycle[ 8286] = 1'b1;  wr_cycle[ 8286] = 1'b0;  addr_rom[ 8286]='h000030f8;  wr_data_rom[ 8286]='h00000000;
    rd_cycle[ 8287] = 1'b0;  wr_cycle[ 8287] = 1'b1;  addr_rom[ 8287]='h0000037c;  wr_data_rom[ 8287]='h000017cf;
    rd_cycle[ 8288] = 1'b0;  wr_cycle[ 8288] = 1'b1;  addr_rom[ 8288]='h0000138c;  wr_data_rom[ 8288]='h00002d2d;
    rd_cycle[ 8289] = 1'b1;  wr_cycle[ 8289] = 1'b0;  addr_rom[ 8289]='h00002c38;  wr_data_rom[ 8289]='h00000000;
    rd_cycle[ 8290] = 1'b1;  wr_cycle[ 8290] = 1'b0;  addr_rom[ 8290]='h000019e0;  wr_data_rom[ 8290]='h00000000;
    rd_cycle[ 8291] = 1'b1;  wr_cycle[ 8291] = 1'b0;  addr_rom[ 8291]='h000024c4;  wr_data_rom[ 8291]='h00000000;
    rd_cycle[ 8292] = 1'b1;  wr_cycle[ 8292] = 1'b0;  addr_rom[ 8292]='h00001a1c;  wr_data_rom[ 8292]='h00000000;
    rd_cycle[ 8293] = 1'b0;  wr_cycle[ 8293] = 1'b1;  addr_rom[ 8293]='h00002bb4;  wr_data_rom[ 8293]='h00002667;
    rd_cycle[ 8294] = 1'b0;  wr_cycle[ 8294] = 1'b1;  addr_rom[ 8294]='h00002ac8;  wr_data_rom[ 8294]='h0000397b;
    rd_cycle[ 8295] = 1'b0;  wr_cycle[ 8295] = 1'b1;  addr_rom[ 8295]='h00001cac;  wr_data_rom[ 8295]='h00001dd1;
    rd_cycle[ 8296] = 1'b1;  wr_cycle[ 8296] = 1'b0;  addr_rom[ 8296]='h00002bd8;  wr_data_rom[ 8296]='h00000000;
    rd_cycle[ 8297] = 1'b0;  wr_cycle[ 8297] = 1'b1;  addr_rom[ 8297]='h00003cd0;  wr_data_rom[ 8297]='h000019cf;
    rd_cycle[ 8298] = 1'b1;  wr_cycle[ 8298] = 1'b0;  addr_rom[ 8298]='h000037d0;  wr_data_rom[ 8298]='h00000000;
    rd_cycle[ 8299] = 1'b0;  wr_cycle[ 8299] = 1'b1;  addr_rom[ 8299]='h00000ed4;  wr_data_rom[ 8299]='h000026ef;
    rd_cycle[ 8300] = 1'b1;  wr_cycle[ 8300] = 1'b0;  addr_rom[ 8300]='h00001390;  wr_data_rom[ 8300]='h00000000;
    rd_cycle[ 8301] = 1'b0;  wr_cycle[ 8301] = 1'b1;  addr_rom[ 8301]='h000022c4;  wr_data_rom[ 8301]='h000034e1;
    rd_cycle[ 8302] = 1'b1;  wr_cycle[ 8302] = 1'b0;  addr_rom[ 8302]='h000009b4;  wr_data_rom[ 8302]='h00000000;
    rd_cycle[ 8303] = 1'b0;  wr_cycle[ 8303] = 1'b1;  addr_rom[ 8303]='h00003f20;  wr_data_rom[ 8303]='h00003659;
    rd_cycle[ 8304] = 1'b1;  wr_cycle[ 8304] = 1'b0;  addr_rom[ 8304]='h000032f0;  wr_data_rom[ 8304]='h00000000;
    rd_cycle[ 8305] = 1'b1;  wr_cycle[ 8305] = 1'b0;  addr_rom[ 8305]='h00001254;  wr_data_rom[ 8305]='h00000000;
    rd_cycle[ 8306] = 1'b1;  wr_cycle[ 8306] = 1'b0;  addr_rom[ 8306]='h000013ec;  wr_data_rom[ 8306]='h00000000;
    rd_cycle[ 8307] = 1'b0;  wr_cycle[ 8307] = 1'b1;  addr_rom[ 8307]='h000032f4;  wr_data_rom[ 8307]='h00000bba;
    rd_cycle[ 8308] = 1'b1;  wr_cycle[ 8308] = 1'b0;  addr_rom[ 8308]='h000011ac;  wr_data_rom[ 8308]='h00000000;
    rd_cycle[ 8309] = 1'b1;  wr_cycle[ 8309] = 1'b0;  addr_rom[ 8309]='h00003d9c;  wr_data_rom[ 8309]='h00000000;
    rd_cycle[ 8310] = 1'b1;  wr_cycle[ 8310] = 1'b0;  addr_rom[ 8310]='h000006cc;  wr_data_rom[ 8310]='h00000000;
    rd_cycle[ 8311] = 1'b0;  wr_cycle[ 8311] = 1'b1;  addr_rom[ 8311]='h00002cc4;  wr_data_rom[ 8311]='h00001da6;
    rd_cycle[ 8312] = 1'b0;  wr_cycle[ 8312] = 1'b1;  addr_rom[ 8312]='h00002e84;  wr_data_rom[ 8312]='h000027aa;
    rd_cycle[ 8313] = 1'b0;  wr_cycle[ 8313] = 1'b1;  addr_rom[ 8313]='h00003778;  wr_data_rom[ 8313]='h00002b00;
    rd_cycle[ 8314] = 1'b1;  wr_cycle[ 8314] = 1'b0;  addr_rom[ 8314]='h000038ec;  wr_data_rom[ 8314]='h00000000;
    rd_cycle[ 8315] = 1'b0;  wr_cycle[ 8315] = 1'b1;  addr_rom[ 8315]='h000009c8;  wr_data_rom[ 8315]='h00003243;
    rd_cycle[ 8316] = 1'b0;  wr_cycle[ 8316] = 1'b1;  addr_rom[ 8316]='h00002cdc;  wr_data_rom[ 8316]='h0000362c;
    rd_cycle[ 8317] = 1'b1;  wr_cycle[ 8317] = 1'b0;  addr_rom[ 8317]='h00003834;  wr_data_rom[ 8317]='h00000000;
    rd_cycle[ 8318] = 1'b1;  wr_cycle[ 8318] = 1'b0;  addr_rom[ 8318]='h00002ba8;  wr_data_rom[ 8318]='h00000000;
    rd_cycle[ 8319] = 1'b0;  wr_cycle[ 8319] = 1'b1;  addr_rom[ 8319]='h000035f8;  wr_data_rom[ 8319]='h00000e5b;
    rd_cycle[ 8320] = 1'b1;  wr_cycle[ 8320] = 1'b0;  addr_rom[ 8320]='h00003524;  wr_data_rom[ 8320]='h00000000;
    rd_cycle[ 8321] = 1'b1;  wr_cycle[ 8321] = 1'b0;  addr_rom[ 8321]='h000011b8;  wr_data_rom[ 8321]='h00000000;
    rd_cycle[ 8322] = 1'b0;  wr_cycle[ 8322] = 1'b1;  addr_rom[ 8322]='h000037f0;  wr_data_rom[ 8322]='h00000c4e;
    rd_cycle[ 8323] = 1'b0;  wr_cycle[ 8323] = 1'b1;  addr_rom[ 8323]='h000036e0;  wr_data_rom[ 8323]='h00003ee5;
    rd_cycle[ 8324] = 1'b1;  wr_cycle[ 8324] = 1'b0;  addr_rom[ 8324]='h00003aa4;  wr_data_rom[ 8324]='h00000000;
    rd_cycle[ 8325] = 1'b0;  wr_cycle[ 8325] = 1'b1;  addr_rom[ 8325]='h00003264;  wr_data_rom[ 8325]='h000014ff;
    rd_cycle[ 8326] = 1'b0;  wr_cycle[ 8326] = 1'b1;  addr_rom[ 8326]='h000022f0;  wr_data_rom[ 8326]='h0000238f;
    rd_cycle[ 8327] = 1'b0;  wr_cycle[ 8327] = 1'b1;  addr_rom[ 8327]='h00000c78;  wr_data_rom[ 8327]='h00002a7b;
    rd_cycle[ 8328] = 1'b0;  wr_cycle[ 8328] = 1'b1;  addr_rom[ 8328]='h00003890;  wr_data_rom[ 8328]='h000001ca;
    rd_cycle[ 8329] = 1'b1;  wr_cycle[ 8329] = 1'b0;  addr_rom[ 8329]='h00001310;  wr_data_rom[ 8329]='h00000000;
    rd_cycle[ 8330] = 1'b1;  wr_cycle[ 8330] = 1'b0;  addr_rom[ 8330]='h00002128;  wr_data_rom[ 8330]='h00000000;
    rd_cycle[ 8331] = 1'b1;  wr_cycle[ 8331] = 1'b0;  addr_rom[ 8331]='h00002f68;  wr_data_rom[ 8331]='h00000000;
    rd_cycle[ 8332] = 1'b0;  wr_cycle[ 8332] = 1'b1;  addr_rom[ 8332]='h00003f08;  wr_data_rom[ 8332]='h000028c7;
    rd_cycle[ 8333] = 1'b1;  wr_cycle[ 8333] = 1'b0;  addr_rom[ 8333]='h00002b14;  wr_data_rom[ 8333]='h00000000;
    rd_cycle[ 8334] = 1'b0;  wr_cycle[ 8334] = 1'b1;  addr_rom[ 8334]='h00001d7c;  wr_data_rom[ 8334]='h00002b8a;
    rd_cycle[ 8335] = 1'b1;  wr_cycle[ 8335] = 1'b0;  addr_rom[ 8335]='h000023e4;  wr_data_rom[ 8335]='h00000000;
    rd_cycle[ 8336] = 1'b1;  wr_cycle[ 8336] = 1'b0;  addr_rom[ 8336]='h00002c28;  wr_data_rom[ 8336]='h00000000;
    rd_cycle[ 8337] = 1'b0;  wr_cycle[ 8337] = 1'b1;  addr_rom[ 8337]='h00001d84;  wr_data_rom[ 8337]='h00001677;
    rd_cycle[ 8338] = 1'b1;  wr_cycle[ 8338] = 1'b0;  addr_rom[ 8338]='h00000708;  wr_data_rom[ 8338]='h00000000;
    rd_cycle[ 8339] = 1'b0;  wr_cycle[ 8339] = 1'b1;  addr_rom[ 8339]='h000030a0;  wr_data_rom[ 8339]='h00001548;
    rd_cycle[ 8340] = 1'b0;  wr_cycle[ 8340] = 1'b1;  addr_rom[ 8340]='h00000834;  wr_data_rom[ 8340]='h000030a1;
    rd_cycle[ 8341] = 1'b1;  wr_cycle[ 8341] = 1'b0;  addr_rom[ 8341]='h00000fb4;  wr_data_rom[ 8341]='h00000000;
    rd_cycle[ 8342] = 1'b0;  wr_cycle[ 8342] = 1'b1;  addr_rom[ 8342]='h000031f8;  wr_data_rom[ 8342]='h00003f60;
    rd_cycle[ 8343] = 1'b0;  wr_cycle[ 8343] = 1'b1;  addr_rom[ 8343]='h000035a4;  wr_data_rom[ 8343]='h00000cdc;
    rd_cycle[ 8344] = 1'b0;  wr_cycle[ 8344] = 1'b1;  addr_rom[ 8344]='h000031a8;  wr_data_rom[ 8344]='h00000442;
    rd_cycle[ 8345] = 1'b1;  wr_cycle[ 8345] = 1'b0;  addr_rom[ 8345]='h00002820;  wr_data_rom[ 8345]='h00000000;
    rd_cycle[ 8346] = 1'b1;  wr_cycle[ 8346] = 1'b0;  addr_rom[ 8346]='h00000820;  wr_data_rom[ 8346]='h00000000;
    rd_cycle[ 8347] = 1'b1;  wr_cycle[ 8347] = 1'b0;  addr_rom[ 8347]='h00001608;  wr_data_rom[ 8347]='h00000000;
    rd_cycle[ 8348] = 1'b0;  wr_cycle[ 8348] = 1'b1;  addr_rom[ 8348]='h00001dd0;  wr_data_rom[ 8348]='h00003fe8;
    rd_cycle[ 8349] = 1'b0;  wr_cycle[ 8349] = 1'b1;  addr_rom[ 8349]='h0000161c;  wr_data_rom[ 8349]='h00000bfe;
    rd_cycle[ 8350] = 1'b1;  wr_cycle[ 8350] = 1'b0;  addr_rom[ 8350]='h000002a8;  wr_data_rom[ 8350]='h00000000;
    rd_cycle[ 8351] = 1'b0;  wr_cycle[ 8351] = 1'b1;  addr_rom[ 8351]='h00003ea8;  wr_data_rom[ 8351]='h00001866;
    rd_cycle[ 8352] = 1'b1;  wr_cycle[ 8352] = 1'b0;  addr_rom[ 8352]='h00002cb8;  wr_data_rom[ 8352]='h00000000;
    rd_cycle[ 8353] = 1'b1;  wr_cycle[ 8353] = 1'b0;  addr_rom[ 8353]='h000023f4;  wr_data_rom[ 8353]='h00000000;
    rd_cycle[ 8354] = 1'b1;  wr_cycle[ 8354] = 1'b0;  addr_rom[ 8354]='h00002578;  wr_data_rom[ 8354]='h00000000;
    rd_cycle[ 8355] = 1'b0;  wr_cycle[ 8355] = 1'b1;  addr_rom[ 8355]='h00003858;  wr_data_rom[ 8355]='h00001951;
    rd_cycle[ 8356] = 1'b0;  wr_cycle[ 8356] = 1'b1;  addr_rom[ 8356]='h000028ac;  wr_data_rom[ 8356]='h0000311c;
    rd_cycle[ 8357] = 1'b0;  wr_cycle[ 8357] = 1'b1;  addr_rom[ 8357]='h000031ec;  wr_data_rom[ 8357]='h00000c9e;
    rd_cycle[ 8358] = 1'b0;  wr_cycle[ 8358] = 1'b1;  addr_rom[ 8358]='h00001488;  wr_data_rom[ 8358]='h00000efe;
    rd_cycle[ 8359] = 1'b1;  wr_cycle[ 8359] = 1'b0;  addr_rom[ 8359]='h000028ac;  wr_data_rom[ 8359]='h00000000;
    rd_cycle[ 8360] = 1'b1;  wr_cycle[ 8360] = 1'b0;  addr_rom[ 8360]='h000026b8;  wr_data_rom[ 8360]='h00000000;
    rd_cycle[ 8361] = 1'b0;  wr_cycle[ 8361] = 1'b1;  addr_rom[ 8361]='h000017b0;  wr_data_rom[ 8361]='h00003ae9;
    rd_cycle[ 8362] = 1'b1;  wr_cycle[ 8362] = 1'b0;  addr_rom[ 8362]='h0000318c;  wr_data_rom[ 8362]='h00000000;
    rd_cycle[ 8363] = 1'b1;  wr_cycle[ 8363] = 1'b0;  addr_rom[ 8363]='h00002c00;  wr_data_rom[ 8363]='h00000000;
    rd_cycle[ 8364] = 1'b1;  wr_cycle[ 8364] = 1'b0;  addr_rom[ 8364]='h00002478;  wr_data_rom[ 8364]='h00000000;
    rd_cycle[ 8365] = 1'b0;  wr_cycle[ 8365] = 1'b1;  addr_rom[ 8365]='h0000051c;  wr_data_rom[ 8365]='h00001bdc;
    rd_cycle[ 8366] = 1'b0;  wr_cycle[ 8366] = 1'b1;  addr_rom[ 8366]='h00000874;  wr_data_rom[ 8366]='h000038f7;
    rd_cycle[ 8367] = 1'b0;  wr_cycle[ 8367] = 1'b1;  addr_rom[ 8367]='h00001aa4;  wr_data_rom[ 8367]='h00000ae5;
    rd_cycle[ 8368] = 1'b1;  wr_cycle[ 8368] = 1'b0;  addr_rom[ 8368]='h000023fc;  wr_data_rom[ 8368]='h00000000;
    rd_cycle[ 8369] = 1'b1;  wr_cycle[ 8369] = 1'b0;  addr_rom[ 8369]='h00000f14;  wr_data_rom[ 8369]='h00000000;
    rd_cycle[ 8370] = 1'b0;  wr_cycle[ 8370] = 1'b1;  addr_rom[ 8370]='h00003e50;  wr_data_rom[ 8370]='h00001860;
    rd_cycle[ 8371] = 1'b1;  wr_cycle[ 8371] = 1'b0;  addr_rom[ 8371]='h00001664;  wr_data_rom[ 8371]='h00000000;
    rd_cycle[ 8372] = 1'b1;  wr_cycle[ 8372] = 1'b0;  addr_rom[ 8372]='h00001a00;  wr_data_rom[ 8372]='h00000000;
    rd_cycle[ 8373] = 1'b1;  wr_cycle[ 8373] = 1'b0;  addr_rom[ 8373]='h0000214c;  wr_data_rom[ 8373]='h00000000;
    rd_cycle[ 8374] = 1'b0;  wr_cycle[ 8374] = 1'b1;  addr_rom[ 8374]='h000022c4;  wr_data_rom[ 8374]='h00003375;
    rd_cycle[ 8375] = 1'b0;  wr_cycle[ 8375] = 1'b1;  addr_rom[ 8375]='h00003eec;  wr_data_rom[ 8375]='h00002d39;
    rd_cycle[ 8376] = 1'b0;  wr_cycle[ 8376] = 1'b1;  addr_rom[ 8376]='h000027a0;  wr_data_rom[ 8376]='h0000260e;
    rd_cycle[ 8377] = 1'b0;  wr_cycle[ 8377] = 1'b1;  addr_rom[ 8377]='h000006ac;  wr_data_rom[ 8377]='h00001269;
    rd_cycle[ 8378] = 1'b1;  wr_cycle[ 8378] = 1'b0;  addr_rom[ 8378]='h00001284;  wr_data_rom[ 8378]='h00000000;
    rd_cycle[ 8379] = 1'b0;  wr_cycle[ 8379] = 1'b1;  addr_rom[ 8379]='h00002f74;  wr_data_rom[ 8379]='h00000823;
    rd_cycle[ 8380] = 1'b0;  wr_cycle[ 8380] = 1'b1;  addr_rom[ 8380]='h00002738;  wr_data_rom[ 8380]='h000023b6;
    rd_cycle[ 8381] = 1'b0;  wr_cycle[ 8381] = 1'b1;  addr_rom[ 8381]='h0000343c;  wr_data_rom[ 8381]='h00002326;
    rd_cycle[ 8382] = 1'b1;  wr_cycle[ 8382] = 1'b0;  addr_rom[ 8382]='h00000c1c;  wr_data_rom[ 8382]='h00000000;
    rd_cycle[ 8383] = 1'b1;  wr_cycle[ 8383] = 1'b0;  addr_rom[ 8383]='h00000460;  wr_data_rom[ 8383]='h00000000;
    rd_cycle[ 8384] = 1'b0;  wr_cycle[ 8384] = 1'b1;  addr_rom[ 8384]='h00001fdc;  wr_data_rom[ 8384]='h00000f05;
    rd_cycle[ 8385] = 1'b1;  wr_cycle[ 8385] = 1'b0;  addr_rom[ 8385]='h000015c8;  wr_data_rom[ 8385]='h00000000;
    rd_cycle[ 8386] = 1'b0;  wr_cycle[ 8386] = 1'b1;  addr_rom[ 8386]='h00000dbc;  wr_data_rom[ 8386]='h000031ec;
    rd_cycle[ 8387] = 1'b0;  wr_cycle[ 8387] = 1'b1;  addr_rom[ 8387]='h00000bc0;  wr_data_rom[ 8387]='h000020c2;
    rd_cycle[ 8388] = 1'b0;  wr_cycle[ 8388] = 1'b1;  addr_rom[ 8388]='h00001920;  wr_data_rom[ 8388]='h0000050c;
    rd_cycle[ 8389] = 1'b1;  wr_cycle[ 8389] = 1'b0;  addr_rom[ 8389]='h00001b40;  wr_data_rom[ 8389]='h00000000;
    rd_cycle[ 8390] = 1'b1;  wr_cycle[ 8390] = 1'b0;  addr_rom[ 8390]='h00002308;  wr_data_rom[ 8390]='h00000000;
    rd_cycle[ 8391] = 1'b1;  wr_cycle[ 8391] = 1'b0;  addr_rom[ 8391]='h00002158;  wr_data_rom[ 8391]='h00000000;
    rd_cycle[ 8392] = 1'b1;  wr_cycle[ 8392] = 1'b0;  addr_rom[ 8392]='h00000b0c;  wr_data_rom[ 8392]='h00000000;
    rd_cycle[ 8393] = 1'b1;  wr_cycle[ 8393] = 1'b0;  addr_rom[ 8393]='h000019d0;  wr_data_rom[ 8393]='h00000000;
    rd_cycle[ 8394] = 1'b1;  wr_cycle[ 8394] = 1'b0;  addr_rom[ 8394]='h00003260;  wr_data_rom[ 8394]='h00000000;
    rd_cycle[ 8395] = 1'b1;  wr_cycle[ 8395] = 1'b0;  addr_rom[ 8395]='h00003824;  wr_data_rom[ 8395]='h00000000;
    rd_cycle[ 8396] = 1'b1;  wr_cycle[ 8396] = 1'b0;  addr_rom[ 8396]='h00003540;  wr_data_rom[ 8396]='h00000000;
    rd_cycle[ 8397] = 1'b1;  wr_cycle[ 8397] = 1'b0;  addr_rom[ 8397]='h00000df0;  wr_data_rom[ 8397]='h00000000;
    rd_cycle[ 8398] = 1'b1;  wr_cycle[ 8398] = 1'b0;  addr_rom[ 8398]='h00002e40;  wr_data_rom[ 8398]='h00000000;
    rd_cycle[ 8399] = 1'b1;  wr_cycle[ 8399] = 1'b0;  addr_rom[ 8399]='h0000389c;  wr_data_rom[ 8399]='h00000000;
    rd_cycle[ 8400] = 1'b0;  wr_cycle[ 8400] = 1'b1;  addr_rom[ 8400]='h0000306c;  wr_data_rom[ 8400]='h00000611;
    rd_cycle[ 8401] = 1'b1;  wr_cycle[ 8401] = 1'b0;  addr_rom[ 8401]='h000013b4;  wr_data_rom[ 8401]='h00000000;
    rd_cycle[ 8402] = 1'b1;  wr_cycle[ 8402] = 1'b0;  addr_rom[ 8402]='h00002670;  wr_data_rom[ 8402]='h00000000;
    rd_cycle[ 8403] = 1'b1;  wr_cycle[ 8403] = 1'b0;  addr_rom[ 8403]='h000009a8;  wr_data_rom[ 8403]='h00000000;
    rd_cycle[ 8404] = 1'b0;  wr_cycle[ 8404] = 1'b1;  addr_rom[ 8404]='h00002088;  wr_data_rom[ 8404]='h0000007d;
    rd_cycle[ 8405] = 1'b1;  wr_cycle[ 8405] = 1'b0;  addr_rom[ 8405]='h00001ce4;  wr_data_rom[ 8405]='h00000000;
    rd_cycle[ 8406] = 1'b1;  wr_cycle[ 8406] = 1'b0;  addr_rom[ 8406]='h00001b54;  wr_data_rom[ 8406]='h00000000;
    rd_cycle[ 8407] = 1'b1;  wr_cycle[ 8407] = 1'b0;  addr_rom[ 8407]='h000036d8;  wr_data_rom[ 8407]='h00000000;
    rd_cycle[ 8408] = 1'b1;  wr_cycle[ 8408] = 1'b0;  addr_rom[ 8408]='h00000794;  wr_data_rom[ 8408]='h00000000;
    rd_cycle[ 8409] = 1'b0;  wr_cycle[ 8409] = 1'b1;  addr_rom[ 8409]='h00002c0c;  wr_data_rom[ 8409]='h00003d63;
    rd_cycle[ 8410] = 1'b1;  wr_cycle[ 8410] = 1'b0;  addr_rom[ 8410]='h000010e8;  wr_data_rom[ 8410]='h00000000;
    rd_cycle[ 8411] = 1'b0;  wr_cycle[ 8411] = 1'b1;  addr_rom[ 8411]='h00001fe0;  wr_data_rom[ 8411]='h00000746;
    rd_cycle[ 8412] = 1'b0;  wr_cycle[ 8412] = 1'b1;  addr_rom[ 8412]='h00001988;  wr_data_rom[ 8412]='h00001ad3;
    rd_cycle[ 8413] = 1'b0;  wr_cycle[ 8413] = 1'b1;  addr_rom[ 8413]='h00001614;  wr_data_rom[ 8413]='h00000fbd;
    rd_cycle[ 8414] = 1'b0;  wr_cycle[ 8414] = 1'b1;  addr_rom[ 8414]='h000005a0;  wr_data_rom[ 8414]='h0000026b;
    rd_cycle[ 8415] = 1'b0;  wr_cycle[ 8415] = 1'b1;  addr_rom[ 8415]='h00003ab4;  wr_data_rom[ 8415]='h00003e74;
    rd_cycle[ 8416] = 1'b1;  wr_cycle[ 8416] = 1'b0;  addr_rom[ 8416]='h00000c90;  wr_data_rom[ 8416]='h00000000;
    rd_cycle[ 8417] = 1'b0;  wr_cycle[ 8417] = 1'b1;  addr_rom[ 8417]='h00003d78;  wr_data_rom[ 8417]='h00003ca5;
    rd_cycle[ 8418] = 1'b1;  wr_cycle[ 8418] = 1'b0;  addr_rom[ 8418]='h00000860;  wr_data_rom[ 8418]='h00000000;
    rd_cycle[ 8419] = 1'b1;  wr_cycle[ 8419] = 1'b0;  addr_rom[ 8419]='h00002714;  wr_data_rom[ 8419]='h00000000;
    rd_cycle[ 8420] = 1'b0;  wr_cycle[ 8420] = 1'b1;  addr_rom[ 8420]='h000039c4;  wr_data_rom[ 8420]='h00003ae1;
    rd_cycle[ 8421] = 1'b1;  wr_cycle[ 8421] = 1'b0;  addr_rom[ 8421]='h000029c4;  wr_data_rom[ 8421]='h00000000;
    rd_cycle[ 8422] = 1'b1;  wr_cycle[ 8422] = 1'b0;  addr_rom[ 8422]='h000035a0;  wr_data_rom[ 8422]='h00000000;
    rd_cycle[ 8423] = 1'b0;  wr_cycle[ 8423] = 1'b1;  addr_rom[ 8423]='h000031ac;  wr_data_rom[ 8423]='h00000ad7;
    rd_cycle[ 8424] = 1'b0;  wr_cycle[ 8424] = 1'b1;  addr_rom[ 8424]='h00000f68;  wr_data_rom[ 8424]='h00001e72;
    rd_cycle[ 8425] = 1'b1;  wr_cycle[ 8425] = 1'b0;  addr_rom[ 8425]='h000035c0;  wr_data_rom[ 8425]='h00000000;
    rd_cycle[ 8426] = 1'b0;  wr_cycle[ 8426] = 1'b1;  addr_rom[ 8426]='h00000220;  wr_data_rom[ 8426]='h000023f3;
    rd_cycle[ 8427] = 1'b1;  wr_cycle[ 8427] = 1'b0;  addr_rom[ 8427]='h00003d50;  wr_data_rom[ 8427]='h00000000;
    rd_cycle[ 8428] = 1'b1;  wr_cycle[ 8428] = 1'b0;  addr_rom[ 8428]='h00002ebc;  wr_data_rom[ 8428]='h00000000;
    rd_cycle[ 8429] = 1'b0;  wr_cycle[ 8429] = 1'b1;  addr_rom[ 8429]='h00003820;  wr_data_rom[ 8429]='h00003caf;
    rd_cycle[ 8430] = 1'b0;  wr_cycle[ 8430] = 1'b1;  addr_rom[ 8430]='h000027e8;  wr_data_rom[ 8430]='h0000228f;
    rd_cycle[ 8431] = 1'b1;  wr_cycle[ 8431] = 1'b0;  addr_rom[ 8431]='h00003d48;  wr_data_rom[ 8431]='h00000000;
    rd_cycle[ 8432] = 1'b1;  wr_cycle[ 8432] = 1'b0;  addr_rom[ 8432]='h000026f8;  wr_data_rom[ 8432]='h00000000;
    rd_cycle[ 8433] = 1'b1;  wr_cycle[ 8433] = 1'b0;  addr_rom[ 8433]='h00002300;  wr_data_rom[ 8433]='h00000000;
    rd_cycle[ 8434] = 1'b0;  wr_cycle[ 8434] = 1'b1;  addr_rom[ 8434]='h000011fc;  wr_data_rom[ 8434]='h00001e7d;
    rd_cycle[ 8435] = 1'b1;  wr_cycle[ 8435] = 1'b0;  addr_rom[ 8435]='h000021a8;  wr_data_rom[ 8435]='h00000000;
    rd_cycle[ 8436] = 1'b0;  wr_cycle[ 8436] = 1'b1;  addr_rom[ 8436]='h00001cf0;  wr_data_rom[ 8436]='h00003a79;
    rd_cycle[ 8437] = 1'b0;  wr_cycle[ 8437] = 1'b1;  addr_rom[ 8437]='h000010d8;  wr_data_rom[ 8437]='h000034c7;
    rd_cycle[ 8438] = 1'b0;  wr_cycle[ 8438] = 1'b1;  addr_rom[ 8438]='h00001744;  wr_data_rom[ 8438]='h00000b15;
    rd_cycle[ 8439] = 1'b1;  wr_cycle[ 8439] = 1'b0;  addr_rom[ 8439]='h000037b8;  wr_data_rom[ 8439]='h00000000;
    rd_cycle[ 8440] = 1'b0;  wr_cycle[ 8440] = 1'b1;  addr_rom[ 8440]='h00002f40;  wr_data_rom[ 8440]='h000013db;
    rd_cycle[ 8441] = 1'b1;  wr_cycle[ 8441] = 1'b0;  addr_rom[ 8441]='h0000007c;  wr_data_rom[ 8441]='h00000000;
    rd_cycle[ 8442] = 1'b0;  wr_cycle[ 8442] = 1'b1;  addr_rom[ 8442]='h00002a04;  wr_data_rom[ 8442]='h00003802;
    rd_cycle[ 8443] = 1'b1;  wr_cycle[ 8443] = 1'b0;  addr_rom[ 8443]='h0000371c;  wr_data_rom[ 8443]='h00000000;
    rd_cycle[ 8444] = 1'b1;  wr_cycle[ 8444] = 1'b0;  addr_rom[ 8444]='h00002054;  wr_data_rom[ 8444]='h00000000;
    rd_cycle[ 8445] = 1'b1;  wr_cycle[ 8445] = 1'b0;  addr_rom[ 8445]='h00002194;  wr_data_rom[ 8445]='h00000000;
    rd_cycle[ 8446] = 1'b0;  wr_cycle[ 8446] = 1'b1;  addr_rom[ 8446]='h00000b54;  wr_data_rom[ 8446]='h000001cb;
    rd_cycle[ 8447] = 1'b1;  wr_cycle[ 8447] = 1'b0;  addr_rom[ 8447]='h00000a14;  wr_data_rom[ 8447]='h00000000;
    rd_cycle[ 8448] = 1'b1;  wr_cycle[ 8448] = 1'b0;  addr_rom[ 8448]='h00000d1c;  wr_data_rom[ 8448]='h00000000;
    rd_cycle[ 8449] = 1'b1;  wr_cycle[ 8449] = 1'b0;  addr_rom[ 8449]='h00000f58;  wr_data_rom[ 8449]='h00000000;
    rd_cycle[ 8450] = 1'b0;  wr_cycle[ 8450] = 1'b1;  addr_rom[ 8450]='h00000038;  wr_data_rom[ 8450]='h0000149e;
    rd_cycle[ 8451] = 1'b1;  wr_cycle[ 8451] = 1'b0;  addr_rom[ 8451]='h00000fc4;  wr_data_rom[ 8451]='h00000000;
    rd_cycle[ 8452] = 1'b0;  wr_cycle[ 8452] = 1'b1;  addr_rom[ 8452]='h00001930;  wr_data_rom[ 8452]='h00001c71;
    rd_cycle[ 8453] = 1'b1;  wr_cycle[ 8453] = 1'b0;  addr_rom[ 8453]='h00001ea4;  wr_data_rom[ 8453]='h00000000;
    rd_cycle[ 8454] = 1'b1;  wr_cycle[ 8454] = 1'b0;  addr_rom[ 8454]='h00001f74;  wr_data_rom[ 8454]='h00000000;
    rd_cycle[ 8455] = 1'b1;  wr_cycle[ 8455] = 1'b0;  addr_rom[ 8455]='h00000260;  wr_data_rom[ 8455]='h00000000;
    rd_cycle[ 8456] = 1'b0;  wr_cycle[ 8456] = 1'b1;  addr_rom[ 8456]='h00003854;  wr_data_rom[ 8456]='h000039dd;
    rd_cycle[ 8457] = 1'b0;  wr_cycle[ 8457] = 1'b1;  addr_rom[ 8457]='h000022d0;  wr_data_rom[ 8457]='h0000332c;
    rd_cycle[ 8458] = 1'b1;  wr_cycle[ 8458] = 1'b0;  addr_rom[ 8458]='h00001aa0;  wr_data_rom[ 8458]='h00000000;
    rd_cycle[ 8459] = 1'b0;  wr_cycle[ 8459] = 1'b1;  addr_rom[ 8459]='h00000b5c;  wr_data_rom[ 8459]='h0000319b;
    rd_cycle[ 8460] = 1'b1;  wr_cycle[ 8460] = 1'b0;  addr_rom[ 8460]='h00002f84;  wr_data_rom[ 8460]='h00000000;
    rd_cycle[ 8461] = 1'b1;  wr_cycle[ 8461] = 1'b0;  addr_rom[ 8461]='h00000b88;  wr_data_rom[ 8461]='h00000000;
    rd_cycle[ 8462] = 1'b0;  wr_cycle[ 8462] = 1'b1;  addr_rom[ 8462]='h00001d44;  wr_data_rom[ 8462]='h00002109;
    rd_cycle[ 8463] = 1'b1;  wr_cycle[ 8463] = 1'b0;  addr_rom[ 8463]='h000008e4;  wr_data_rom[ 8463]='h00000000;
    rd_cycle[ 8464] = 1'b1;  wr_cycle[ 8464] = 1'b0;  addr_rom[ 8464]='h00001528;  wr_data_rom[ 8464]='h00000000;
    rd_cycle[ 8465] = 1'b0;  wr_cycle[ 8465] = 1'b1;  addr_rom[ 8465]='h00003cc0;  wr_data_rom[ 8465]='h00002fb8;
    rd_cycle[ 8466] = 1'b0;  wr_cycle[ 8466] = 1'b1;  addr_rom[ 8466]='h00003020;  wr_data_rom[ 8466]='h000015dc;
    rd_cycle[ 8467] = 1'b1;  wr_cycle[ 8467] = 1'b0;  addr_rom[ 8467]='h000013dc;  wr_data_rom[ 8467]='h00000000;
    rd_cycle[ 8468] = 1'b0;  wr_cycle[ 8468] = 1'b1;  addr_rom[ 8468]='h00003aac;  wr_data_rom[ 8468]='h00001d2e;
    rd_cycle[ 8469] = 1'b1;  wr_cycle[ 8469] = 1'b0;  addr_rom[ 8469]='h00002530;  wr_data_rom[ 8469]='h00000000;
    rd_cycle[ 8470] = 1'b1;  wr_cycle[ 8470] = 1'b0;  addr_rom[ 8470]='h000033f0;  wr_data_rom[ 8470]='h00000000;
    rd_cycle[ 8471] = 1'b1;  wr_cycle[ 8471] = 1'b0;  addr_rom[ 8471]='h00000954;  wr_data_rom[ 8471]='h00000000;
    rd_cycle[ 8472] = 1'b1;  wr_cycle[ 8472] = 1'b0;  addr_rom[ 8472]='h0000198c;  wr_data_rom[ 8472]='h00000000;
    rd_cycle[ 8473] = 1'b1;  wr_cycle[ 8473] = 1'b0;  addr_rom[ 8473]='h00000590;  wr_data_rom[ 8473]='h00000000;
    rd_cycle[ 8474] = 1'b1;  wr_cycle[ 8474] = 1'b0;  addr_rom[ 8474]='h000021f0;  wr_data_rom[ 8474]='h00000000;
    rd_cycle[ 8475] = 1'b0;  wr_cycle[ 8475] = 1'b1;  addr_rom[ 8475]='h000005e4;  wr_data_rom[ 8475]='h00001785;
    rd_cycle[ 8476] = 1'b1;  wr_cycle[ 8476] = 1'b0;  addr_rom[ 8476]='h00001038;  wr_data_rom[ 8476]='h00000000;
    rd_cycle[ 8477] = 1'b1;  wr_cycle[ 8477] = 1'b0;  addr_rom[ 8477]='h000021c8;  wr_data_rom[ 8477]='h00000000;
    rd_cycle[ 8478] = 1'b0;  wr_cycle[ 8478] = 1'b1;  addr_rom[ 8478]='h00001d3c;  wr_data_rom[ 8478]='h000005f7;
    rd_cycle[ 8479] = 1'b0;  wr_cycle[ 8479] = 1'b1;  addr_rom[ 8479]='h00000b24;  wr_data_rom[ 8479]='h00002d15;
    rd_cycle[ 8480] = 1'b0;  wr_cycle[ 8480] = 1'b1;  addr_rom[ 8480]='h00000cec;  wr_data_rom[ 8480]='h00002059;
    rd_cycle[ 8481] = 1'b1;  wr_cycle[ 8481] = 1'b0;  addr_rom[ 8481]='h00002e80;  wr_data_rom[ 8481]='h00000000;
    rd_cycle[ 8482] = 1'b1;  wr_cycle[ 8482] = 1'b0;  addr_rom[ 8482]='h00003650;  wr_data_rom[ 8482]='h00000000;
    rd_cycle[ 8483] = 1'b0;  wr_cycle[ 8483] = 1'b1;  addr_rom[ 8483]='h000036f4;  wr_data_rom[ 8483]='h00003a81;
    rd_cycle[ 8484] = 1'b1;  wr_cycle[ 8484] = 1'b0;  addr_rom[ 8484]='h00003e7c;  wr_data_rom[ 8484]='h00000000;
    rd_cycle[ 8485] = 1'b1;  wr_cycle[ 8485] = 1'b0;  addr_rom[ 8485]='h00001f24;  wr_data_rom[ 8485]='h00000000;
    rd_cycle[ 8486] = 1'b0;  wr_cycle[ 8486] = 1'b1;  addr_rom[ 8486]='h00002d4c;  wr_data_rom[ 8486]='h000005e6;
    rd_cycle[ 8487] = 1'b0;  wr_cycle[ 8487] = 1'b1;  addr_rom[ 8487]='h00001bbc;  wr_data_rom[ 8487]='h00001c67;
    rd_cycle[ 8488] = 1'b0;  wr_cycle[ 8488] = 1'b1;  addr_rom[ 8488]='h00003864;  wr_data_rom[ 8488]='h00002ddd;
    rd_cycle[ 8489] = 1'b0;  wr_cycle[ 8489] = 1'b1;  addr_rom[ 8489]='h000000f4;  wr_data_rom[ 8489]='h0000089c;
    rd_cycle[ 8490] = 1'b0;  wr_cycle[ 8490] = 1'b1;  addr_rom[ 8490]='h00001028;  wr_data_rom[ 8490]='h00000cca;
    rd_cycle[ 8491] = 1'b0;  wr_cycle[ 8491] = 1'b1;  addr_rom[ 8491]='h00001b3c;  wr_data_rom[ 8491]='h00002af1;
    rd_cycle[ 8492] = 1'b0;  wr_cycle[ 8492] = 1'b1;  addr_rom[ 8492]='h00003b54;  wr_data_rom[ 8492]='h00002ff3;
    rd_cycle[ 8493] = 1'b1;  wr_cycle[ 8493] = 1'b0;  addr_rom[ 8493]='h00001eb0;  wr_data_rom[ 8493]='h00000000;
    rd_cycle[ 8494] = 1'b1;  wr_cycle[ 8494] = 1'b0;  addr_rom[ 8494]='h0000217c;  wr_data_rom[ 8494]='h00000000;
    rd_cycle[ 8495] = 1'b1;  wr_cycle[ 8495] = 1'b0;  addr_rom[ 8495]='h00003eac;  wr_data_rom[ 8495]='h00000000;
    rd_cycle[ 8496] = 1'b0;  wr_cycle[ 8496] = 1'b1;  addr_rom[ 8496]='h00001f20;  wr_data_rom[ 8496]='h000032a4;
    rd_cycle[ 8497] = 1'b0;  wr_cycle[ 8497] = 1'b1;  addr_rom[ 8497]='h0000244c;  wr_data_rom[ 8497]='h00003e98;
    rd_cycle[ 8498] = 1'b1;  wr_cycle[ 8498] = 1'b0;  addr_rom[ 8498]='h00002424;  wr_data_rom[ 8498]='h00000000;
    rd_cycle[ 8499] = 1'b0;  wr_cycle[ 8499] = 1'b1;  addr_rom[ 8499]='h000021cc;  wr_data_rom[ 8499]='h00001379;
    rd_cycle[ 8500] = 1'b0;  wr_cycle[ 8500] = 1'b1;  addr_rom[ 8500]='h0000367c;  wr_data_rom[ 8500]='h00001980;
    rd_cycle[ 8501] = 1'b0;  wr_cycle[ 8501] = 1'b1;  addr_rom[ 8501]='h0000348c;  wr_data_rom[ 8501]='h000027d1;
    rd_cycle[ 8502] = 1'b0;  wr_cycle[ 8502] = 1'b1;  addr_rom[ 8502]='h00001810;  wr_data_rom[ 8502]='h00001fbd;
    rd_cycle[ 8503] = 1'b0;  wr_cycle[ 8503] = 1'b1;  addr_rom[ 8503]='h000009a8;  wr_data_rom[ 8503]='h0000319a;
    rd_cycle[ 8504] = 1'b1;  wr_cycle[ 8504] = 1'b0;  addr_rom[ 8504]='h00001c6c;  wr_data_rom[ 8504]='h00000000;
    rd_cycle[ 8505] = 1'b1;  wr_cycle[ 8505] = 1'b0;  addr_rom[ 8505]='h00002b58;  wr_data_rom[ 8505]='h00000000;
    rd_cycle[ 8506] = 1'b0;  wr_cycle[ 8506] = 1'b1;  addr_rom[ 8506]='h000007e0;  wr_data_rom[ 8506]='h000033f7;
    rd_cycle[ 8507] = 1'b1;  wr_cycle[ 8507] = 1'b0;  addr_rom[ 8507]='h00002870;  wr_data_rom[ 8507]='h00000000;
    rd_cycle[ 8508] = 1'b0;  wr_cycle[ 8508] = 1'b1;  addr_rom[ 8508]='h00002884;  wr_data_rom[ 8508]='h0000035a;
    rd_cycle[ 8509] = 1'b0;  wr_cycle[ 8509] = 1'b1;  addr_rom[ 8509]='h00003e88;  wr_data_rom[ 8509]='h00000cbf;
    rd_cycle[ 8510] = 1'b0;  wr_cycle[ 8510] = 1'b1;  addr_rom[ 8510]='h00000744;  wr_data_rom[ 8510]='h0000070a;
    rd_cycle[ 8511] = 1'b0;  wr_cycle[ 8511] = 1'b1;  addr_rom[ 8511]='h00001cbc;  wr_data_rom[ 8511]='h00002113;
    rd_cycle[ 8512] = 1'b0;  wr_cycle[ 8512] = 1'b1;  addr_rom[ 8512]='h00003064;  wr_data_rom[ 8512]='h000012ed;
    rd_cycle[ 8513] = 1'b0;  wr_cycle[ 8513] = 1'b1;  addr_rom[ 8513]='h00003b68;  wr_data_rom[ 8513]='h000035f6;
    rd_cycle[ 8514] = 1'b1;  wr_cycle[ 8514] = 1'b0;  addr_rom[ 8514]='h000009ec;  wr_data_rom[ 8514]='h00000000;
    rd_cycle[ 8515] = 1'b1;  wr_cycle[ 8515] = 1'b0;  addr_rom[ 8515]='h00003360;  wr_data_rom[ 8515]='h00000000;
    rd_cycle[ 8516] = 1'b0;  wr_cycle[ 8516] = 1'b1;  addr_rom[ 8516]='h00003ab4;  wr_data_rom[ 8516]='h0000212c;
    rd_cycle[ 8517] = 1'b0;  wr_cycle[ 8517] = 1'b1;  addr_rom[ 8517]='h00003af0;  wr_data_rom[ 8517]='h0000064b;
    rd_cycle[ 8518] = 1'b0;  wr_cycle[ 8518] = 1'b1;  addr_rom[ 8518]='h00002230;  wr_data_rom[ 8518]='h00001816;
    rd_cycle[ 8519] = 1'b1;  wr_cycle[ 8519] = 1'b0;  addr_rom[ 8519]='h00000090;  wr_data_rom[ 8519]='h00000000;
    rd_cycle[ 8520] = 1'b0;  wr_cycle[ 8520] = 1'b1;  addr_rom[ 8520]='h00003564;  wr_data_rom[ 8520]='h00000f99;
    rd_cycle[ 8521] = 1'b1;  wr_cycle[ 8521] = 1'b0;  addr_rom[ 8521]='h000007a8;  wr_data_rom[ 8521]='h00000000;
    rd_cycle[ 8522] = 1'b1;  wr_cycle[ 8522] = 1'b0;  addr_rom[ 8522]='h00003c24;  wr_data_rom[ 8522]='h00000000;
    rd_cycle[ 8523] = 1'b0;  wr_cycle[ 8523] = 1'b1;  addr_rom[ 8523]='h0000048c;  wr_data_rom[ 8523]='h00001f64;
    rd_cycle[ 8524] = 1'b0;  wr_cycle[ 8524] = 1'b1;  addr_rom[ 8524]='h00001310;  wr_data_rom[ 8524]='h00003217;
    rd_cycle[ 8525] = 1'b1;  wr_cycle[ 8525] = 1'b0;  addr_rom[ 8525]='h00001ea8;  wr_data_rom[ 8525]='h00000000;
    rd_cycle[ 8526] = 1'b1;  wr_cycle[ 8526] = 1'b0;  addr_rom[ 8526]='h00002ebc;  wr_data_rom[ 8526]='h00000000;
    rd_cycle[ 8527] = 1'b1;  wr_cycle[ 8527] = 1'b0;  addr_rom[ 8527]='h0000323c;  wr_data_rom[ 8527]='h00000000;
    rd_cycle[ 8528] = 1'b1;  wr_cycle[ 8528] = 1'b0;  addr_rom[ 8528]='h00002b28;  wr_data_rom[ 8528]='h00000000;
    rd_cycle[ 8529] = 1'b0;  wr_cycle[ 8529] = 1'b1;  addr_rom[ 8529]='h00003060;  wr_data_rom[ 8529]='h00003718;
    rd_cycle[ 8530] = 1'b1;  wr_cycle[ 8530] = 1'b0;  addr_rom[ 8530]='h00000208;  wr_data_rom[ 8530]='h00000000;
    rd_cycle[ 8531] = 1'b1;  wr_cycle[ 8531] = 1'b0;  addr_rom[ 8531]='h00000b90;  wr_data_rom[ 8531]='h00000000;
    rd_cycle[ 8532] = 1'b1;  wr_cycle[ 8532] = 1'b0;  addr_rom[ 8532]='h0000024c;  wr_data_rom[ 8532]='h00000000;
    rd_cycle[ 8533] = 1'b1;  wr_cycle[ 8533] = 1'b0;  addr_rom[ 8533]='h00002c24;  wr_data_rom[ 8533]='h00000000;
    rd_cycle[ 8534] = 1'b1;  wr_cycle[ 8534] = 1'b0;  addr_rom[ 8534]='h000006d0;  wr_data_rom[ 8534]='h00000000;
    rd_cycle[ 8535] = 1'b1;  wr_cycle[ 8535] = 1'b0;  addr_rom[ 8535]='h00001e6c;  wr_data_rom[ 8535]='h00000000;
    rd_cycle[ 8536] = 1'b0;  wr_cycle[ 8536] = 1'b1;  addr_rom[ 8536]='h0000339c;  wr_data_rom[ 8536]='h0000316b;
    rd_cycle[ 8537] = 1'b1;  wr_cycle[ 8537] = 1'b0;  addr_rom[ 8537]='h00002574;  wr_data_rom[ 8537]='h00000000;
    rd_cycle[ 8538] = 1'b0;  wr_cycle[ 8538] = 1'b1;  addr_rom[ 8538]='h00003844;  wr_data_rom[ 8538]='h00001c7c;
    rd_cycle[ 8539] = 1'b1;  wr_cycle[ 8539] = 1'b0;  addr_rom[ 8539]='h000019b4;  wr_data_rom[ 8539]='h00000000;
    rd_cycle[ 8540] = 1'b1;  wr_cycle[ 8540] = 1'b0;  addr_rom[ 8540]='h00003180;  wr_data_rom[ 8540]='h00000000;
    rd_cycle[ 8541] = 1'b0;  wr_cycle[ 8541] = 1'b1;  addr_rom[ 8541]='h00000698;  wr_data_rom[ 8541]='h00001685;
    rd_cycle[ 8542] = 1'b0;  wr_cycle[ 8542] = 1'b1;  addr_rom[ 8542]='h00003018;  wr_data_rom[ 8542]='h00003e71;
    rd_cycle[ 8543] = 1'b1;  wr_cycle[ 8543] = 1'b0;  addr_rom[ 8543]='h00001590;  wr_data_rom[ 8543]='h00000000;
    rd_cycle[ 8544] = 1'b1;  wr_cycle[ 8544] = 1'b0;  addr_rom[ 8544]='h000009f8;  wr_data_rom[ 8544]='h00000000;
    rd_cycle[ 8545] = 1'b1;  wr_cycle[ 8545] = 1'b0;  addr_rom[ 8545]='h00000420;  wr_data_rom[ 8545]='h00000000;
    rd_cycle[ 8546] = 1'b1;  wr_cycle[ 8546] = 1'b0;  addr_rom[ 8546]='h000022a0;  wr_data_rom[ 8546]='h00000000;
    rd_cycle[ 8547] = 1'b1;  wr_cycle[ 8547] = 1'b0;  addr_rom[ 8547]='h000006bc;  wr_data_rom[ 8547]='h00000000;
    rd_cycle[ 8548] = 1'b0;  wr_cycle[ 8548] = 1'b1;  addr_rom[ 8548]='h000038ac;  wr_data_rom[ 8548]='h00001515;
    rd_cycle[ 8549] = 1'b0;  wr_cycle[ 8549] = 1'b1;  addr_rom[ 8549]='h00003788;  wr_data_rom[ 8549]='h00002c10;
    rd_cycle[ 8550] = 1'b0;  wr_cycle[ 8550] = 1'b1;  addr_rom[ 8550]='h0000164c;  wr_data_rom[ 8550]='h00002f02;
    rd_cycle[ 8551] = 1'b0;  wr_cycle[ 8551] = 1'b1;  addr_rom[ 8551]='h00001560;  wr_data_rom[ 8551]='h00003396;
    rd_cycle[ 8552] = 1'b1;  wr_cycle[ 8552] = 1'b0;  addr_rom[ 8552]='h000005d4;  wr_data_rom[ 8552]='h00000000;
    rd_cycle[ 8553] = 1'b1;  wr_cycle[ 8553] = 1'b0;  addr_rom[ 8553]='h00002f38;  wr_data_rom[ 8553]='h00000000;
    rd_cycle[ 8554] = 1'b1;  wr_cycle[ 8554] = 1'b0;  addr_rom[ 8554]='h00000230;  wr_data_rom[ 8554]='h00000000;
    rd_cycle[ 8555] = 1'b1;  wr_cycle[ 8555] = 1'b0;  addr_rom[ 8555]='h00001230;  wr_data_rom[ 8555]='h00000000;
    rd_cycle[ 8556] = 1'b1;  wr_cycle[ 8556] = 1'b0;  addr_rom[ 8556]='h000011f4;  wr_data_rom[ 8556]='h00000000;
    rd_cycle[ 8557] = 1'b1;  wr_cycle[ 8557] = 1'b0;  addr_rom[ 8557]='h00002568;  wr_data_rom[ 8557]='h00000000;
    rd_cycle[ 8558] = 1'b1;  wr_cycle[ 8558] = 1'b0;  addr_rom[ 8558]='h00000004;  wr_data_rom[ 8558]='h00000000;
    rd_cycle[ 8559] = 1'b1;  wr_cycle[ 8559] = 1'b0;  addr_rom[ 8559]='h00002488;  wr_data_rom[ 8559]='h00000000;
    rd_cycle[ 8560] = 1'b0;  wr_cycle[ 8560] = 1'b1;  addr_rom[ 8560]='h00000a9c;  wr_data_rom[ 8560]='h000006b2;
    rd_cycle[ 8561] = 1'b0;  wr_cycle[ 8561] = 1'b1;  addr_rom[ 8561]='h00002a34;  wr_data_rom[ 8561]='h00002276;
    rd_cycle[ 8562] = 1'b1;  wr_cycle[ 8562] = 1'b0;  addr_rom[ 8562]='h00001d90;  wr_data_rom[ 8562]='h00000000;
    rd_cycle[ 8563] = 1'b1;  wr_cycle[ 8563] = 1'b0;  addr_rom[ 8563]='h00002e98;  wr_data_rom[ 8563]='h00000000;
    rd_cycle[ 8564] = 1'b1;  wr_cycle[ 8564] = 1'b0;  addr_rom[ 8564]='h00000f80;  wr_data_rom[ 8564]='h00000000;
    rd_cycle[ 8565] = 1'b0;  wr_cycle[ 8565] = 1'b1;  addr_rom[ 8565]='h000019a4;  wr_data_rom[ 8565]='h0000001c;
    rd_cycle[ 8566] = 1'b1;  wr_cycle[ 8566] = 1'b0;  addr_rom[ 8566]='h00003dcc;  wr_data_rom[ 8566]='h00000000;
    rd_cycle[ 8567] = 1'b1;  wr_cycle[ 8567] = 1'b0;  addr_rom[ 8567]='h000014fc;  wr_data_rom[ 8567]='h00000000;
    rd_cycle[ 8568] = 1'b0;  wr_cycle[ 8568] = 1'b1;  addr_rom[ 8568]='h00000184;  wr_data_rom[ 8568]='h00000471;
    rd_cycle[ 8569] = 1'b0;  wr_cycle[ 8569] = 1'b1;  addr_rom[ 8569]='h000009d4;  wr_data_rom[ 8569]='h00001eaf;
    rd_cycle[ 8570] = 1'b1;  wr_cycle[ 8570] = 1'b0;  addr_rom[ 8570]='h000027ac;  wr_data_rom[ 8570]='h00000000;
    rd_cycle[ 8571] = 1'b1;  wr_cycle[ 8571] = 1'b0;  addr_rom[ 8571]='h00002a84;  wr_data_rom[ 8571]='h00000000;
    rd_cycle[ 8572] = 1'b0;  wr_cycle[ 8572] = 1'b1;  addr_rom[ 8572]='h000009b8;  wr_data_rom[ 8572]='h00003aab;
    rd_cycle[ 8573] = 1'b0;  wr_cycle[ 8573] = 1'b1;  addr_rom[ 8573]='h00000b80;  wr_data_rom[ 8573]='h000011cd;
    rd_cycle[ 8574] = 1'b1;  wr_cycle[ 8574] = 1'b0;  addr_rom[ 8574]='h00000908;  wr_data_rom[ 8574]='h00000000;
    rd_cycle[ 8575] = 1'b0;  wr_cycle[ 8575] = 1'b1;  addr_rom[ 8575]='h00003ca8;  wr_data_rom[ 8575]='h00003e01;
    rd_cycle[ 8576] = 1'b0;  wr_cycle[ 8576] = 1'b1;  addr_rom[ 8576]='h00003268;  wr_data_rom[ 8576]='h00003b0f;
    rd_cycle[ 8577] = 1'b1;  wr_cycle[ 8577] = 1'b0;  addr_rom[ 8577]='h000021a0;  wr_data_rom[ 8577]='h00000000;
    rd_cycle[ 8578] = 1'b0;  wr_cycle[ 8578] = 1'b1;  addr_rom[ 8578]='h00000a3c;  wr_data_rom[ 8578]='h000039b4;
    rd_cycle[ 8579] = 1'b1;  wr_cycle[ 8579] = 1'b0;  addr_rom[ 8579]='h00003e4c;  wr_data_rom[ 8579]='h00000000;
    rd_cycle[ 8580] = 1'b1;  wr_cycle[ 8580] = 1'b0;  addr_rom[ 8580]='h00000338;  wr_data_rom[ 8580]='h00000000;
    rd_cycle[ 8581] = 1'b1;  wr_cycle[ 8581] = 1'b0;  addr_rom[ 8581]='h000009fc;  wr_data_rom[ 8581]='h00000000;
    rd_cycle[ 8582] = 1'b0;  wr_cycle[ 8582] = 1'b1;  addr_rom[ 8582]='h000020f0;  wr_data_rom[ 8582]='h00000fe5;
    rd_cycle[ 8583] = 1'b1;  wr_cycle[ 8583] = 1'b0;  addr_rom[ 8583]='h0000233c;  wr_data_rom[ 8583]='h00000000;
    rd_cycle[ 8584] = 1'b1;  wr_cycle[ 8584] = 1'b0;  addr_rom[ 8584]='h00003b00;  wr_data_rom[ 8584]='h00000000;
    rd_cycle[ 8585] = 1'b1;  wr_cycle[ 8585] = 1'b0;  addr_rom[ 8585]='h00000c24;  wr_data_rom[ 8585]='h00000000;
    rd_cycle[ 8586] = 1'b0;  wr_cycle[ 8586] = 1'b1;  addr_rom[ 8586]='h00002b80;  wr_data_rom[ 8586]='h00003336;
    rd_cycle[ 8587] = 1'b1;  wr_cycle[ 8587] = 1'b0;  addr_rom[ 8587]='h0000166c;  wr_data_rom[ 8587]='h00000000;
    rd_cycle[ 8588] = 1'b0;  wr_cycle[ 8588] = 1'b1;  addr_rom[ 8588]='h000014a0;  wr_data_rom[ 8588]='h00001186;
    rd_cycle[ 8589] = 1'b0;  wr_cycle[ 8589] = 1'b1;  addr_rom[ 8589]='h00002f18;  wr_data_rom[ 8589]='h00002346;
    rd_cycle[ 8590] = 1'b0;  wr_cycle[ 8590] = 1'b1;  addr_rom[ 8590]='h000038bc;  wr_data_rom[ 8590]='h0000202e;
    rd_cycle[ 8591] = 1'b0;  wr_cycle[ 8591] = 1'b1;  addr_rom[ 8591]='h000031d0;  wr_data_rom[ 8591]='h00000249;
    rd_cycle[ 8592] = 1'b1;  wr_cycle[ 8592] = 1'b0;  addr_rom[ 8592]='h00002dc8;  wr_data_rom[ 8592]='h00000000;
    rd_cycle[ 8593] = 1'b1;  wr_cycle[ 8593] = 1'b0;  addr_rom[ 8593]='h0000113c;  wr_data_rom[ 8593]='h00000000;
    rd_cycle[ 8594] = 1'b1;  wr_cycle[ 8594] = 1'b0;  addr_rom[ 8594]='h0000340c;  wr_data_rom[ 8594]='h00000000;
    rd_cycle[ 8595] = 1'b1;  wr_cycle[ 8595] = 1'b0;  addr_rom[ 8595]='h000029d8;  wr_data_rom[ 8595]='h00000000;
    rd_cycle[ 8596] = 1'b1;  wr_cycle[ 8596] = 1'b0;  addr_rom[ 8596]='h00002aa8;  wr_data_rom[ 8596]='h00000000;
    rd_cycle[ 8597] = 1'b1;  wr_cycle[ 8597] = 1'b0;  addr_rom[ 8597]='h000028bc;  wr_data_rom[ 8597]='h00000000;
    rd_cycle[ 8598] = 1'b0;  wr_cycle[ 8598] = 1'b1;  addr_rom[ 8598]='h00001f6c;  wr_data_rom[ 8598]='h000017c1;
    rd_cycle[ 8599] = 1'b0;  wr_cycle[ 8599] = 1'b1;  addr_rom[ 8599]='h000011a0;  wr_data_rom[ 8599]='h00003af0;
    rd_cycle[ 8600] = 1'b0;  wr_cycle[ 8600] = 1'b1;  addr_rom[ 8600]='h00001efc;  wr_data_rom[ 8600]='h00000a2c;
    rd_cycle[ 8601] = 1'b0;  wr_cycle[ 8601] = 1'b1;  addr_rom[ 8601]='h00000a28;  wr_data_rom[ 8601]='h00003a3c;
    rd_cycle[ 8602] = 1'b1;  wr_cycle[ 8602] = 1'b0;  addr_rom[ 8602]='h000021cc;  wr_data_rom[ 8602]='h00000000;
    rd_cycle[ 8603] = 1'b0;  wr_cycle[ 8603] = 1'b1;  addr_rom[ 8603]='h00003790;  wr_data_rom[ 8603]='h000013b9;
    rd_cycle[ 8604] = 1'b0;  wr_cycle[ 8604] = 1'b1;  addr_rom[ 8604]='h000016b8;  wr_data_rom[ 8604]='h00001eba;
    rd_cycle[ 8605] = 1'b0;  wr_cycle[ 8605] = 1'b1;  addr_rom[ 8605]='h00002724;  wr_data_rom[ 8605]='h00002928;
    rd_cycle[ 8606] = 1'b0;  wr_cycle[ 8606] = 1'b1;  addr_rom[ 8606]='h00001508;  wr_data_rom[ 8606]='h00001ca7;
    rd_cycle[ 8607] = 1'b1;  wr_cycle[ 8607] = 1'b0;  addr_rom[ 8607]='h00002720;  wr_data_rom[ 8607]='h00000000;
    rd_cycle[ 8608] = 1'b1;  wr_cycle[ 8608] = 1'b0;  addr_rom[ 8608]='h00002778;  wr_data_rom[ 8608]='h00000000;
    rd_cycle[ 8609] = 1'b0;  wr_cycle[ 8609] = 1'b1;  addr_rom[ 8609]='h0000372c;  wr_data_rom[ 8609]='h0000132e;
    rd_cycle[ 8610] = 1'b0;  wr_cycle[ 8610] = 1'b1;  addr_rom[ 8610]='h00003934;  wr_data_rom[ 8610]='h00003717;
    rd_cycle[ 8611] = 1'b0;  wr_cycle[ 8611] = 1'b1;  addr_rom[ 8611]='h000023a4;  wr_data_rom[ 8611]='h00003156;
    rd_cycle[ 8612] = 1'b0;  wr_cycle[ 8612] = 1'b1;  addr_rom[ 8612]='h00001ee0;  wr_data_rom[ 8612]='h000030ef;
    rd_cycle[ 8613] = 1'b0;  wr_cycle[ 8613] = 1'b1;  addr_rom[ 8613]='h000007d4;  wr_data_rom[ 8613]='h00002e28;
    rd_cycle[ 8614] = 1'b1;  wr_cycle[ 8614] = 1'b0;  addr_rom[ 8614]='h00003afc;  wr_data_rom[ 8614]='h00000000;
    rd_cycle[ 8615] = 1'b0;  wr_cycle[ 8615] = 1'b1;  addr_rom[ 8615]='h00003774;  wr_data_rom[ 8615]='h0000076a;
    rd_cycle[ 8616] = 1'b0;  wr_cycle[ 8616] = 1'b1;  addr_rom[ 8616]='h00003c58;  wr_data_rom[ 8616]='h0000094f;
    rd_cycle[ 8617] = 1'b1;  wr_cycle[ 8617] = 1'b0;  addr_rom[ 8617]='h00003d74;  wr_data_rom[ 8617]='h00000000;
    rd_cycle[ 8618] = 1'b0;  wr_cycle[ 8618] = 1'b1;  addr_rom[ 8618]='h00003130;  wr_data_rom[ 8618]='h0000038f;
    rd_cycle[ 8619] = 1'b1;  wr_cycle[ 8619] = 1'b0;  addr_rom[ 8619]='h000011e0;  wr_data_rom[ 8619]='h00000000;
    rd_cycle[ 8620] = 1'b1;  wr_cycle[ 8620] = 1'b0;  addr_rom[ 8620]='h00002474;  wr_data_rom[ 8620]='h00000000;
    rd_cycle[ 8621] = 1'b1;  wr_cycle[ 8621] = 1'b0;  addr_rom[ 8621]='h000027c8;  wr_data_rom[ 8621]='h00000000;
    rd_cycle[ 8622] = 1'b0;  wr_cycle[ 8622] = 1'b1;  addr_rom[ 8622]='h00002a3c;  wr_data_rom[ 8622]='h00000698;
    rd_cycle[ 8623] = 1'b1;  wr_cycle[ 8623] = 1'b0;  addr_rom[ 8623]='h00000748;  wr_data_rom[ 8623]='h00000000;
    rd_cycle[ 8624] = 1'b1;  wr_cycle[ 8624] = 1'b0;  addr_rom[ 8624]='h00001dd0;  wr_data_rom[ 8624]='h00000000;
    rd_cycle[ 8625] = 1'b0;  wr_cycle[ 8625] = 1'b1;  addr_rom[ 8625]='h00003470;  wr_data_rom[ 8625]='h00003639;
    rd_cycle[ 8626] = 1'b0;  wr_cycle[ 8626] = 1'b1;  addr_rom[ 8626]='h00002af0;  wr_data_rom[ 8626]='h00001877;
    rd_cycle[ 8627] = 1'b0;  wr_cycle[ 8627] = 1'b1;  addr_rom[ 8627]='h00000d00;  wr_data_rom[ 8627]='h00003b27;
    rd_cycle[ 8628] = 1'b0;  wr_cycle[ 8628] = 1'b1;  addr_rom[ 8628]='h000011f4;  wr_data_rom[ 8628]='h00003414;
    rd_cycle[ 8629] = 1'b1;  wr_cycle[ 8629] = 1'b0;  addr_rom[ 8629]='h00000090;  wr_data_rom[ 8629]='h00000000;
    rd_cycle[ 8630] = 1'b1;  wr_cycle[ 8630] = 1'b0;  addr_rom[ 8630]='h00001ee0;  wr_data_rom[ 8630]='h00000000;
    rd_cycle[ 8631] = 1'b0;  wr_cycle[ 8631] = 1'b1;  addr_rom[ 8631]='h00002c80;  wr_data_rom[ 8631]='h00000f58;
    rd_cycle[ 8632] = 1'b1;  wr_cycle[ 8632] = 1'b0;  addr_rom[ 8632]='h00000928;  wr_data_rom[ 8632]='h00000000;
    rd_cycle[ 8633] = 1'b1;  wr_cycle[ 8633] = 1'b0;  addr_rom[ 8633]='h00000050;  wr_data_rom[ 8633]='h00000000;
    rd_cycle[ 8634] = 1'b1;  wr_cycle[ 8634] = 1'b0;  addr_rom[ 8634]='h00002a34;  wr_data_rom[ 8634]='h00000000;
    rd_cycle[ 8635] = 1'b1;  wr_cycle[ 8635] = 1'b0;  addr_rom[ 8635]='h00002be8;  wr_data_rom[ 8635]='h00000000;
    rd_cycle[ 8636] = 1'b1;  wr_cycle[ 8636] = 1'b0;  addr_rom[ 8636]='h00000118;  wr_data_rom[ 8636]='h00000000;
    rd_cycle[ 8637] = 1'b0;  wr_cycle[ 8637] = 1'b1;  addr_rom[ 8637]='h000011c0;  wr_data_rom[ 8637]='h0000053c;
    rd_cycle[ 8638] = 1'b0;  wr_cycle[ 8638] = 1'b1;  addr_rom[ 8638]='h00002d6c;  wr_data_rom[ 8638]='h00003265;
    rd_cycle[ 8639] = 1'b0;  wr_cycle[ 8639] = 1'b1;  addr_rom[ 8639]='h00001504;  wr_data_rom[ 8639]='h000032f9;
    rd_cycle[ 8640] = 1'b1;  wr_cycle[ 8640] = 1'b0;  addr_rom[ 8640]='h00000108;  wr_data_rom[ 8640]='h00000000;
    rd_cycle[ 8641] = 1'b0;  wr_cycle[ 8641] = 1'b1;  addr_rom[ 8641]='h00003698;  wr_data_rom[ 8641]='h00000ce3;
    rd_cycle[ 8642] = 1'b0;  wr_cycle[ 8642] = 1'b1;  addr_rom[ 8642]='h00000e70;  wr_data_rom[ 8642]='h00003a54;
    rd_cycle[ 8643] = 1'b0;  wr_cycle[ 8643] = 1'b1;  addr_rom[ 8643]='h000015b8;  wr_data_rom[ 8643]='h0000110a;
    rd_cycle[ 8644] = 1'b0;  wr_cycle[ 8644] = 1'b1;  addr_rom[ 8644]='h00001768;  wr_data_rom[ 8644]='h0000217c;
    rd_cycle[ 8645] = 1'b0;  wr_cycle[ 8645] = 1'b1;  addr_rom[ 8645]='h0000149c;  wr_data_rom[ 8645]='h00000326;
    rd_cycle[ 8646] = 1'b0;  wr_cycle[ 8646] = 1'b1;  addr_rom[ 8646]='h00000978;  wr_data_rom[ 8646]='h00003e8c;
    rd_cycle[ 8647] = 1'b1;  wr_cycle[ 8647] = 1'b0;  addr_rom[ 8647]='h00001b2c;  wr_data_rom[ 8647]='h00000000;
    rd_cycle[ 8648] = 1'b0;  wr_cycle[ 8648] = 1'b1;  addr_rom[ 8648]='h00000b14;  wr_data_rom[ 8648]='h000023be;
    rd_cycle[ 8649] = 1'b1;  wr_cycle[ 8649] = 1'b0;  addr_rom[ 8649]='h000002fc;  wr_data_rom[ 8649]='h00000000;
    rd_cycle[ 8650] = 1'b1;  wr_cycle[ 8650] = 1'b0;  addr_rom[ 8650]='h000004b0;  wr_data_rom[ 8650]='h00000000;
    rd_cycle[ 8651] = 1'b1;  wr_cycle[ 8651] = 1'b0;  addr_rom[ 8651]='h000033f0;  wr_data_rom[ 8651]='h00000000;
    rd_cycle[ 8652] = 1'b1;  wr_cycle[ 8652] = 1'b0;  addr_rom[ 8652]='h00000078;  wr_data_rom[ 8652]='h00000000;
    rd_cycle[ 8653] = 1'b0;  wr_cycle[ 8653] = 1'b1;  addr_rom[ 8653]='h00000734;  wr_data_rom[ 8653]='h00002009;
    rd_cycle[ 8654] = 1'b0;  wr_cycle[ 8654] = 1'b1;  addr_rom[ 8654]='h000002f4;  wr_data_rom[ 8654]='h00003603;
    rd_cycle[ 8655] = 1'b1;  wr_cycle[ 8655] = 1'b0;  addr_rom[ 8655]='h00002d74;  wr_data_rom[ 8655]='h00000000;
    rd_cycle[ 8656] = 1'b1;  wr_cycle[ 8656] = 1'b0;  addr_rom[ 8656]='h00001574;  wr_data_rom[ 8656]='h00000000;
    rd_cycle[ 8657] = 1'b1;  wr_cycle[ 8657] = 1'b0;  addr_rom[ 8657]='h00000c68;  wr_data_rom[ 8657]='h00000000;
    rd_cycle[ 8658] = 1'b0;  wr_cycle[ 8658] = 1'b1;  addr_rom[ 8658]='h000017bc;  wr_data_rom[ 8658]='h000017fb;
    rd_cycle[ 8659] = 1'b1;  wr_cycle[ 8659] = 1'b0;  addr_rom[ 8659]='h00001b04;  wr_data_rom[ 8659]='h00000000;
    rd_cycle[ 8660] = 1'b0;  wr_cycle[ 8660] = 1'b1;  addr_rom[ 8660]='h00001268;  wr_data_rom[ 8660]='h00003142;
    rd_cycle[ 8661] = 1'b1;  wr_cycle[ 8661] = 1'b0;  addr_rom[ 8661]='h00003b08;  wr_data_rom[ 8661]='h00000000;
    rd_cycle[ 8662] = 1'b1;  wr_cycle[ 8662] = 1'b0;  addr_rom[ 8662]='h00000958;  wr_data_rom[ 8662]='h00000000;
    rd_cycle[ 8663] = 1'b0;  wr_cycle[ 8663] = 1'b1;  addr_rom[ 8663]='h00003878;  wr_data_rom[ 8663]='h000006e6;
    rd_cycle[ 8664] = 1'b0;  wr_cycle[ 8664] = 1'b1;  addr_rom[ 8664]='h00002bc8;  wr_data_rom[ 8664]='h0000024b;
    rd_cycle[ 8665] = 1'b1;  wr_cycle[ 8665] = 1'b0;  addr_rom[ 8665]='h00001820;  wr_data_rom[ 8665]='h00000000;
    rd_cycle[ 8666] = 1'b0;  wr_cycle[ 8666] = 1'b1;  addr_rom[ 8666]='h00002ee8;  wr_data_rom[ 8666]='h00001816;
    rd_cycle[ 8667] = 1'b0;  wr_cycle[ 8667] = 1'b1;  addr_rom[ 8667]='h00000de0;  wr_data_rom[ 8667]='h00001f1b;
    rd_cycle[ 8668] = 1'b0;  wr_cycle[ 8668] = 1'b1;  addr_rom[ 8668]='h00001c8c;  wr_data_rom[ 8668]='h00002c0b;
    rd_cycle[ 8669] = 1'b1;  wr_cycle[ 8669] = 1'b0;  addr_rom[ 8669]='h000002fc;  wr_data_rom[ 8669]='h00000000;
    rd_cycle[ 8670] = 1'b0;  wr_cycle[ 8670] = 1'b1;  addr_rom[ 8670]='h00002a38;  wr_data_rom[ 8670]='h00001771;
    rd_cycle[ 8671] = 1'b0;  wr_cycle[ 8671] = 1'b1;  addr_rom[ 8671]='h00000d10;  wr_data_rom[ 8671]='h000006b1;
    rd_cycle[ 8672] = 1'b1;  wr_cycle[ 8672] = 1'b0;  addr_rom[ 8672]='h00001274;  wr_data_rom[ 8672]='h00000000;
    rd_cycle[ 8673] = 1'b0;  wr_cycle[ 8673] = 1'b1;  addr_rom[ 8673]='h00000284;  wr_data_rom[ 8673]='h00002e1e;
    rd_cycle[ 8674] = 1'b1;  wr_cycle[ 8674] = 1'b0;  addr_rom[ 8674]='h00002d1c;  wr_data_rom[ 8674]='h00000000;
    rd_cycle[ 8675] = 1'b1;  wr_cycle[ 8675] = 1'b0;  addr_rom[ 8675]='h000020d8;  wr_data_rom[ 8675]='h00000000;
    rd_cycle[ 8676] = 1'b0;  wr_cycle[ 8676] = 1'b1;  addr_rom[ 8676]='h00000094;  wr_data_rom[ 8676]='h000030ba;
    rd_cycle[ 8677] = 1'b1;  wr_cycle[ 8677] = 1'b0;  addr_rom[ 8677]='h00002008;  wr_data_rom[ 8677]='h00000000;
    rd_cycle[ 8678] = 1'b0;  wr_cycle[ 8678] = 1'b1;  addr_rom[ 8678]='h00003990;  wr_data_rom[ 8678]='h00003af5;
    rd_cycle[ 8679] = 1'b0;  wr_cycle[ 8679] = 1'b1;  addr_rom[ 8679]='h00003374;  wr_data_rom[ 8679]='h00001ebe;
    rd_cycle[ 8680] = 1'b1;  wr_cycle[ 8680] = 1'b0;  addr_rom[ 8680]='h00000594;  wr_data_rom[ 8680]='h00000000;
    rd_cycle[ 8681] = 1'b0;  wr_cycle[ 8681] = 1'b1;  addr_rom[ 8681]='h00000cfc;  wr_data_rom[ 8681]='h000004a0;
    rd_cycle[ 8682] = 1'b1;  wr_cycle[ 8682] = 1'b0;  addr_rom[ 8682]='h00003b40;  wr_data_rom[ 8682]='h00000000;
    rd_cycle[ 8683] = 1'b0;  wr_cycle[ 8683] = 1'b1;  addr_rom[ 8683]='h00002b28;  wr_data_rom[ 8683]='h000018ef;
    rd_cycle[ 8684] = 1'b0;  wr_cycle[ 8684] = 1'b1;  addr_rom[ 8684]='h00000054;  wr_data_rom[ 8684]='h00001650;
    rd_cycle[ 8685] = 1'b1;  wr_cycle[ 8685] = 1'b0;  addr_rom[ 8685]='h00000948;  wr_data_rom[ 8685]='h00000000;
    rd_cycle[ 8686] = 1'b1;  wr_cycle[ 8686] = 1'b0;  addr_rom[ 8686]='h00003270;  wr_data_rom[ 8686]='h00000000;
    rd_cycle[ 8687] = 1'b0;  wr_cycle[ 8687] = 1'b1;  addr_rom[ 8687]='h00001c1c;  wr_data_rom[ 8687]='h00000f83;
    rd_cycle[ 8688] = 1'b0;  wr_cycle[ 8688] = 1'b1;  addr_rom[ 8688]='h000009d0;  wr_data_rom[ 8688]='h00000299;
    rd_cycle[ 8689] = 1'b0;  wr_cycle[ 8689] = 1'b1;  addr_rom[ 8689]='h00003180;  wr_data_rom[ 8689]='h000032a8;
    rd_cycle[ 8690] = 1'b0;  wr_cycle[ 8690] = 1'b1;  addr_rom[ 8690]='h00003d20;  wr_data_rom[ 8690]='h000014d9;
    rd_cycle[ 8691] = 1'b1;  wr_cycle[ 8691] = 1'b0;  addr_rom[ 8691]='h00002520;  wr_data_rom[ 8691]='h00000000;
    rd_cycle[ 8692] = 1'b1;  wr_cycle[ 8692] = 1'b0;  addr_rom[ 8692]='h00003e88;  wr_data_rom[ 8692]='h00000000;
    rd_cycle[ 8693] = 1'b0;  wr_cycle[ 8693] = 1'b1;  addr_rom[ 8693]='h00003608;  wr_data_rom[ 8693]='h00001c5e;
    rd_cycle[ 8694] = 1'b1;  wr_cycle[ 8694] = 1'b0;  addr_rom[ 8694]='h00002ff8;  wr_data_rom[ 8694]='h00000000;
    rd_cycle[ 8695] = 1'b0;  wr_cycle[ 8695] = 1'b1;  addr_rom[ 8695]='h00000c90;  wr_data_rom[ 8695]='h00000402;
    rd_cycle[ 8696] = 1'b0;  wr_cycle[ 8696] = 1'b1;  addr_rom[ 8696]='h000034ec;  wr_data_rom[ 8696]='h00000095;
    rd_cycle[ 8697] = 1'b1;  wr_cycle[ 8697] = 1'b0;  addr_rom[ 8697]='h00001e38;  wr_data_rom[ 8697]='h00000000;
    rd_cycle[ 8698] = 1'b0;  wr_cycle[ 8698] = 1'b1;  addr_rom[ 8698]='h00002e5c;  wr_data_rom[ 8698]='h000008e0;
    rd_cycle[ 8699] = 1'b1;  wr_cycle[ 8699] = 1'b0;  addr_rom[ 8699]='h00001f94;  wr_data_rom[ 8699]='h00000000;
    rd_cycle[ 8700] = 1'b1;  wr_cycle[ 8700] = 1'b0;  addr_rom[ 8700]='h00002a48;  wr_data_rom[ 8700]='h00000000;
    rd_cycle[ 8701] = 1'b0;  wr_cycle[ 8701] = 1'b1;  addr_rom[ 8701]='h000008d4;  wr_data_rom[ 8701]='h000019eb;
    rd_cycle[ 8702] = 1'b1;  wr_cycle[ 8702] = 1'b0;  addr_rom[ 8702]='h000030e0;  wr_data_rom[ 8702]='h00000000;
    rd_cycle[ 8703] = 1'b1;  wr_cycle[ 8703] = 1'b0;  addr_rom[ 8703]='h00000600;  wr_data_rom[ 8703]='h00000000;
    rd_cycle[ 8704] = 1'b0;  wr_cycle[ 8704] = 1'b1;  addr_rom[ 8704]='h00001424;  wr_data_rom[ 8704]='h00001e7f;
    rd_cycle[ 8705] = 1'b1;  wr_cycle[ 8705] = 1'b0;  addr_rom[ 8705]='h00000454;  wr_data_rom[ 8705]='h00000000;
    rd_cycle[ 8706] = 1'b0;  wr_cycle[ 8706] = 1'b1;  addr_rom[ 8706]='h00002bc8;  wr_data_rom[ 8706]='h00002c62;
    rd_cycle[ 8707] = 1'b0;  wr_cycle[ 8707] = 1'b1;  addr_rom[ 8707]='h00003050;  wr_data_rom[ 8707]='h00002731;
    rd_cycle[ 8708] = 1'b1;  wr_cycle[ 8708] = 1'b0;  addr_rom[ 8708]='h00002924;  wr_data_rom[ 8708]='h00000000;
    rd_cycle[ 8709] = 1'b1;  wr_cycle[ 8709] = 1'b0;  addr_rom[ 8709]='h00002f14;  wr_data_rom[ 8709]='h00000000;
    rd_cycle[ 8710] = 1'b1;  wr_cycle[ 8710] = 1'b0;  addr_rom[ 8710]='h00000508;  wr_data_rom[ 8710]='h00000000;
    rd_cycle[ 8711] = 1'b0;  wr_cycle[ 8711] = 1'b1;  addr_rom[ 8711]='h000033b0;  wr_data_rom[ 8711]='h000028d4;
    rd_cycle[ 8712] = 1'b0;  wr_cycle[ 8712] = 1'b1;  addr_rom[ 8712]='h00001074;  wr_data_rom[ 8712]='h00000def;
    rd_cycle[ 8713] = 1'b1;  wr_cycle[ 8713] = 1'b0;  addr_rom[ 8713]='h00003910;  wr_data_rom[ 8713]='h00000000;
    rd_cycle[ 8714] = 1'b1;  wr_cycle[ 8714] = 1'b0;  addr_rom[ 8714]='h00002fa0;  wr_data_rom[ 8714]='h00000000;
    rd_cycle[ 8715] = 1'b1;  wr_cycle[ 8715] = 1'b0;  addr_rom[ 8715]='h000029e0;  wr_data_rom[ 8715]='h00000000;
    rd_cycle[ 8716] = 1'b1;  wr_cycle[ 8716] = 1'b0;  addr_rom[ 8716]='h00002bf4;  wr_data_rom[ 8716]='h00000000;
    rd_cycle[ 8717] = 1'b1;  wr_cycle[ 8717] = 1'b0;  addr_rom[ 8717]='h000019e8;  wr_data_rom[ 8717]='h00000000;
    rd_cycle[ 8718] = 1'b1;  wr_cycle[ 8718] = 1'b0;  addr_rom[ 8718]='h000007b4;  wr_data_rom[ 8718]='h00000000;
    rd_cycle[ 8719] = 1'b0;  wr_cycle[ 8719] = 1'b1;  addr_rom[ 8719]='h00003bcc;  wr_data_rom[ 8719]='h00003cc8;
    rd_cycle[ 8720] = 1'b1;  wr_cycle[ 8720] = 1'b0;  addr_rom[ 8720]='h00000804;  wr_data_rom[ 8720]='h00000000;
    rd_cycle[ 8721] = 1'b1;  wr_cycle[ 8721] = 1'b0;  addr_rom[ 8721]='h00003b7c;  wr_data_rom[ 8721]='h00000000;
    rd_cycle[ 8722] = 1'b0;  wr_cycle[ 8722] = 1'b1;  addr_rom[ 8722]='h0000385c;  wr_data_rom[ 8722]='h00000fcd;
    rd_cycle[ 8723] = 1'b1;  wr_cycle[ 8723] = 1'b0;  addr_rom[ 8723]='h00000eb4;  wr_data_rom[ 8723]='h00000000;
    rd_cycle[ 8724] = 1'b1;  wr_cycle[ 8724] = 1'b0;  addr_rom[ 8724]='h00002d40;  wr_data_rom[ 8724]='h00000000;
    rd_cycle[ 8725] = 1'b1;  wr_cycle[ 8725] = 1'b0;  addr_rom[ 8725]='h00002c28;  wr_data_rom[ 8725]='h00000000;
    rd_cycle[ 8726] = 1'b0;  wr_cycle[ 8726] = 1'b1;  addr_rom[ 8726]='h00001d78;  wr_data_rom[ 8726]='h00001219;
    rd_cycle[ 8727] = 1'b1;  wr_cycle[ 8727] = 1'b0;  addr_rom[ 8727]='h00002ff8;  wr_data_rom[ 8727]='h00000000;
    rd_cycle[ 8728] = 1'b1;  wr_cycle[ 8728] = 1'b0;  addr_rom[ 8728]='h000015b0;  wr_data_rom[ 8728]='h00000000;
    rd_cycle[ 8729] = 1'b1;  wr_cycle[ 8729] = 1'b0;  addr_rom[ 8729]='h000024f8;  wr_data_rom[ 8729]='h00000000;
    rd_cycle[ 8730] = 1'b1;  wr_cycle[ 8730] = 1'b0;  addr_rom[ 8730]='h00002d44;  wr_data_rom[ 8730]='h00000000;
    rd_cycle[ 8731] = 1'b0;  wr_cycle[ 8731] = 1'b1;  addr_rom[ 8731]='h00003de0;  wr_data_rom[ 8731]='h0000237b;
    rd_cycle[ 8732] = 1'b1;  wr_cycle[ 8732] = 1'b0;  addr_rom[ 8732]='h00001674;  wr_data_rom[ 8732]='h00000000;
    rd_cycle[ 8733] = 1'b0;  wr_cycle[ 8733] = 1'b1;  addr_rom[ 8733]='h00000b44;  wr_data_rom[ 8733]='h0000223e;
    rd_cycle[ 8734] = 1'b1;  wr_cycle[ 8734] = 1'b0;  addr_rom[ 8734]='h00001f3c;  wr_data_rom[ 8734]='h00000000;
    rd_cycle[ 8735] = 1'b0;  wr_cycle[ 8735] = 1'b1;  addr_rom[ 8735]='h00002988;  wr_data_rom[ 8735]='h00003997;
    rd_cycle[ 8736] = 1'b1;  wr_cycle[ 8736] = 1'b0;  addr_rom[ 8736]='h00003380;  wr_data_rom[ 8736]='h00000000;
    rd_cycle[ 8737] = 1'b0;  wr_cycle[ 8737] = 1'b1;  addr_rom[ 8737]='h00003708;  wr_data_rom[ 8737]='h00003497;
    rd_cycle[ 8738] = 1'b0;  wr_cycle[ 8738] = 1'b1;  addr_rom[ 8738]='h00001afc;  wr_data_rom[ 8738]='h00001eaf;
    rd_cycle[ 8739] = 1'b0;  wr_cycle[ 8739] = 1'b1;  addr_rom[ 8739]='h00000684;  wr_data_rom[ 8739]='h00002fbd;
    rd_cycle[ 8740] = 1'b1;  wr_cycle[ 8740] = 1'b0;  addr_rom[ 8740]='h00002240;  wr_data_rom[ 8740]='h00000000;
    rd_cycle[ 8741] = 1'b0;  wr_cycle[ 8741] = 1'b1;  addr_rom[ 8741]='h0000173c;  wr_data_rom[ 8741]='h00002a1a;
    rd_cycle[ 8742] = 1'b0;  wr_cycle[ 8742] = 1'b1;  addr_rom[ 8742]='h00002b00;  wr_data_rom[ 8742]='h00000f32;
    rd_cycle[ 8743] = 1'b1;  wr_cycle[ 8743] = 1'b0;  addr_rom[ 8743]='h00000400;  wr_data_rom[ 8743]='h00000000;
    rd_cycle[ 8744] = 1'b0;  wr_cycle[ 8744] = 1'b1;  addr_rom[ 8744]='h000004cc;  wr_data_rom[ 8744]='h00001a87;
    rd_cycle[ 8745] = 1'b0;  wr_cycle[ 8745] = 1'b1;  addr_rom[ 8745]='h00001720;  wr_data_rom[ 8745]='h000005e8;
    rd_cycle[ 8746] = 1'b1;  wr_cycle[ 8746] = 1'b0;  addr_rom[ 8746]='h00002940;  wr_data_rom[ 8746]='h00000000;
    rd_cycle[ 8747] = 1'b1;  wr_cycle[ 8747] = 1'b0;  addr_rom[ 8747]='h0000036c;  wr_data_rom[ 8747]='h00000000;
    rd_cycle[ 8748] = 1'b1;  wr_cycle[ 8748] = 1'b0;  addr_rom[ 8748]='h000010c4;  wr_data_rom[ 8748]='h00000000;
    rd_cycle[ 8749] = 1'b0;  wr_cycle[ 8749] = 1'b1;  addr_rom[ 8749]='h00001a6c;  wr_data_rom[ 8749]='h00001591;
    rd_cycle[ 8750] = 1'b1;  wr_cycle[ 8750] = 1'b0;  addr_rom[ 8750]='h00003584;  wr_data_rom[ 8750]='h00000000;
    rd_cycle[ 8751] = 1'b1;  wr_cycle[ 8751] = 1'b0;  addr_rom[ 8751]='h000022cc;  wr_data_rom[ 8751]='h00000000;
    rd_cycle[ 8752] = 1'b1;  wr_cycle[ 8752] = 1'b0;  addr_rom[ 8752]='h0000305c;  wr_data_rom[ 8752]='h00000000;
    rd_cycle[ 8753] = 1'b0;  wr_cycle[ 8753] = 1'b1;  addr_rom[ 8753]='h000008fc;  wr_data_rom[ 8753]='h0000001f;
    rd_cycle[ 8754] = 1'b1;  wr_cycle[ 8754] = 1'b0;  addr_rom[ 8754]='h00003524;  wr_data_rom[ 8754]='h00000000;
    rd_cycle[ 8755] = 1'b0;  wr_cycle[ 8755] = 1'b1;  addr_rom[ 8755]='h00002408;  wr_data_rom[ 8755]='h00001bb8;
    rd_cycle[ 8756] = 1'b1;  wr_cycle[ 8756] = 1'b0;  addr_rom[ 8756]='h00001f58;  wr_data_rom[ 8756]='h00000000;
    rd_cycle[ 8757] = 1'b0;  wr_cycle[ 8757] = 1'b1;  addr_rom[ 8757]='h00000340;  wr_data_rom[ 8757]='h00002bdd;
    rd_cycle[ 8758] = 1'b1;  wr_cycle[ 8758] = 1'b0;  addr_rom[ 8758]='h000015e0;  wr_data_rom[ 8758]='h00000000;
    rd_cycle[ 8759] = 1'b1;  wr_cycle[ 8759] = 1'b0;  addr_rom[ 8759]='h00001f80;  wr_data_rom[ 8759]='h00000000;
    rd_cycle[ 8760] = 1'b0;  wr_cycle[ 8760] = 1'b1;  addr_rom[ 8760]='h000018f0;  wr_data_rom[ 8760]='h00001f7b;
    rd_cycle[ 8761] = 1'b1;  wr_cycle[ 8761] = 1'b0;  addr_rom[ 8761]='h00001120;  wr_data_rom[ 8761]='h00000000;
    rd_cycle[ 8762] = 1'b1;  wr_cycle[ 8762] = 1'b0;  addr_rom[ 8762]='h0000054c;  wr_data_rom[ 8762]='h00000000;
    rd_cycle[ 8763] = 1'b1;  wr_cycle[ 8763] = 1'b0;  addr_rom[ 8763]='h00000908;  wr_data_rom[ 8763]='h00000000;
    rd_cycle[ 8764] = 1'b0;  wr_cycle[ 8764] = 1'b1;  addr_rom[ 8764]='h00002318;  wr_data_rom[ 8764]='h000016e9;
    rd_cycle[ 8765] = 1'b1;  wr_cycle[ 8765] = 1'b0;  addr_rom[ 8765]='h00002504;  wr_data_rom[ 8765]='h00000000;
    rd_cycle[ 8766] = 1'b0;  wr_cycle[ 8766] = 1'b1;  addr_rom[ 8766]='h00002d3c;  wr_data_rom[ 8766]='h000011ee;
    rd_cycle[ 8767] = 1'b1;  wr_cycle[ 8767] = 1'b0;  addr_rom[ 8767]='h0000101c;  wr_data_rom[ 8767]='h00000000;
    rd_cycle[ 8768] = 1'b1;  wr_cycle[ 8768] = 1'b0;  addr_rom[ 8768]='h00003fbc;  wr_data_rom[ 8768]='h00000000;
    rd_cycle[ 8769] = 1'b1;  wr_cycle[ 8769] = 1'b0;  addr_rom[ 8769]='h000023c0;  wr_data_rom[ 8769]='h00000000;
    rd_cycle[ 8770] = 1'b1;  wr_cycle[ 8770] = 1'b0;  addr_rom[ 8770]='h0000268c;  wr_data_rom[ 8770]='h00000000;
    rd_cycle[ 8771] = 1'b1;  wr_cycle[ 8771] = 1'b0;  addr_rom[ 8771]='h00001f98;  wr_data_rom[ 8771]='h00000000;
    rd_cycle[ 8772] = 1'b0;  wr_cycle[ 8772] = 1'b1;  addr_rom[ 8772]='h00000974;  wr_data_rom[ 8772]='h00003d64;
    rd_cycle[ 8773] = 1'b1;  wr_cycle[ 8773] = 1'b0;  addr_rom[ 8773]='h0000160c;  wr_data_rom[ 8773]='h00000000;
    rd_cycle[ 8774] = 1'b1;  wr_cycle[ 8774] = 1'b0;  addr_rom[ 8774]='h00003168;  wr_data_rom[ 8774]='h00000000;
    rd_cycle[ 8775] = 1'b1;  wr_cycle[ 8775] = 1'b0;  addr_rom[ 8775]='h00003b00;  wr_data_rom[ 8775]='h00000000;
    rd_cycle[ 8776] = 1'b0;  wr_cycle[ 8776] = 1'b1;  addr_rom[ 8776]='h00001d8c;  wr_data_rom[ 8776]='h000038c4;
    rd_cycle[ 8777] = 1'b1;  wr_cycle[ 8777] = 1'b0;  addr_rom[ 8777]='h000014fc;  wr_data_rom[ 8777]='h00000000;
    rd_cycle[ 8778] = 1'b1;  wr_cycle[ 8778] = 1'b0;  addr_rom[ 8778]='h000009c0;  wr_data_rom[ 8778]='h00000000;
    rd_cycle[ 8779] = 1'b0;  wr_cycle[ 8779] = 1'b1;  addr_rom[ 8779]='h00000748;  wr_data_rom[ 8779]='h00003a89;
    rd_cycle[ 8780] = 1'b1;  wr_cycle[ 8780] = 1'b0;  addr_rom[ 8780]='h00002878;  wr_data_rom[ 8780]='h00000000;
    rd_cycle[ 8781] = 1'b1;  wr_cycle[ 8781] = 1'b0;  addr_rom[ 8781]='h00001b28;  wr_data_rom[ 8781]='h00000000;
    rd_cycle[ 8782] = 1'b0;  wr_cycle[ 8782] = 1'b1;  addr_rom[ 8782]='h00000b20;  wr_data_rom[ 8782]='h00003d27;
    rd_cycle[ 8783] = 1'b0;  wr_cycle[ 8783] = 1'b1;  addr_rom[ 8783]='h00003634;  wr_data_rom[ 8783]='h000036e8;
    rd_cycle[ 8784] = 1'b0;  wr_cycle[ 8784] = 1'b1;  addr_rom[ 8784]='h00000e8c;  wr_data_rom[ 8784]='h000035f7;
    rd_cycle[ 8785] = 1'b1;  wr_cycle[ 8785] = 1'b0;  addr_rom[ 8785]='h000021b8;  wr_data_rom[ 8785]='h00000000;
    rd_cycle[ 8786] = 1'b1;  wr_cycle[ 8786] = 1'b0;  addr_rom[ 8786]='h00003cdc;  wr_data_rom[ 8786]='h00000000;
    rd_cycle[ 8787] = 1'b0;  wr_cycle[ 8787] = 1'b1;  addr_rom[ 8787]='h000034b4;  wr_data_rom[ 8787]='h00001b48;
    rd_cycle[ 8788] = 1'b0;  wr_cycle[ 8788] = 1'b1;  addr_rom[ 8788]='h0000172c;  wr_data_rom[ 8788]='h0000388e;
    rd_cycle[ 8789] = 1'b0;  wr_cycle[ 8789] = 1'b1;  addr_rom[ 8789]='h00003050;  wr_data_rom[ 8789]='h00003ff8;
    rd_cycle[ 8790] = 1'b1;  wr_cycle[ 8790] = 1'b0;  addr_rom[ 8790]='h000020ac;  wr_data_rom[ 8790]='h00000000;
    rd_cycle[ 8791] = 1'b0;  wr_cycle[ 8791] = 1'b1;  addr_rom[ 8791]='h00003524;  wr_data_rom[ 8791]='h000005ff;
    rd_cycle[ 8792] = 1'b1;  wr_cycle[ 8792] = 1'b0;  addr_rom[ 8792]='h000039e8;  wr_data_rom[ 8792]='h00000000;
    rd_cycle[ 8793] = 1'b0;  wr_cycle[ 8793] = 1'b1;  addr_rom[ 8793]='h00001e7c;  wr_data_rom[ 8793]='h00002535;
    rd_cycle[ 8794] = 1'b0;  wr_cycle[ 8794] = 1'b1;  addr_rom[ 8794]='h00002088;  wr_data_rom[ 8794]='h00003572;
    rd_cycle[ 8795] = 1'b0;  wr_cycle[ 8795] = 1'b1;  addr_rom[ 8795]='h000029fc;  wr_data_rom[ 8795]='h00003ba5;
    rd_cycle[ 8796] = 1'b0;  wr_cycle[ 8796] = 1'b1;  addr_rom[ 8796]='h0000347c;  wr_data_rom[ 8796]='h0000385f;
    rd_cycle[ 8797] = 1'b1;  wr_cycle[ 8797] = 1'b0;  addr_rom[ 8797]='h0000325c;  wr_data_rom[ 8797]='h00000000;
    rd_cycle[ 8798] = 1'b0;  wr_cycle[ 8798] = 1'b1;  addr_rom[ 8798]='h00003c14;  wr_data_rom[ 8798]='h000034a1;
    rd_cycle[ 8799] = 1'b1;  wr_cycle[ 8799] = 1'b0;  addr_rom[ 8799]='h0000315c;  wr_data_rom[ 8799]='h00000000;
    rd_cycle[ 8800] = 1'b0;  wr_cycle[ 8800] = 1'b1;  addr_rom[ 8800]='h00003fb4;  wr_data_rom[ 8800]='h00002593;
    rd_cycle[ 8801] = 1'b0;  wr_cycle[ 8801] = 1'b1;  addr_rom[ 8801]='h000034e8;  wr_data_rom[ 8801]='h000007be;
    rd_cycle[ 8802] = 1'b0;  wr_cycle[ 8802] = 1'b1;  addr_rom[ 8802]='h00002530;  wr_data_rom[ 8802]='h00002ebe;
    rd_cycle[ 8803] = 1'b1;  wr_cycle[ 8803] = 1'b0;  addr_rom[ 8803]='h00001260;  wr_data_rom[ 8803]='h00000000;
    rd_cycle[ 8804] = 1'b1;  wr_cycle[ 8804] = 1'b0;  addr_rom[ 8804]='h000007dc;  wr_data_rom[ 8804]='h00000000;
    rd_cycle[ 8805] = 1'b1;  wr_cycle[ 8805] = 1'b0;  addr_rom[ 8805]='h0000382c;  wr_data_rom[ 8805]='h00000000;
    rd_cycle[ 8806] = 1'b1;  wr_cycle[ 8806] = 1'b0;  addr_rom[ 8806]='h00000e44;  wr_data_rom[ 8806]='h00000000;
    rd_cycle[ 8807] = 1'b1;  wr_cycle[ 8807] = 1'b0;  addr_rom[ 8807]='h000036dc;  wr_data_rom[ 8807]='h00000000;
    rd_cycle[ 8808] = 1'b0;  wr_cycle[ 8808] = 1'b1;  addr_rom[ 8808]='h00000b24;  wr_data_rom[ 8808]='h00002a01;
    rd_cycle[ 8809] = 1'b0;  wr_cycle[ 8809] = 1'b1;  addr_rom[ 8809]='h0000353c;  wr_data_rom[ 8809]='h00000211;
    rd_cycle[ 8810] = 1'b0;  wr_cycle[ 8810] = 1'b1;  addr_rom[ 8810]='h000037cc;  wr_data_rom[ 8810]='h00000f4c;
    rd_cycle[ 8811] = 1'b1;  wr_cycle[ 8811] = 1'b0;  addr_rom[ 8811]='h000015d4;  wr_data_rom[ 8811]='h00000000;
    rd_cycle[ 8812] = 1'b1;  wr_cycle[ 8812] = 1'b0;  addr_rom[ 8812]='h00000724;  wr_data_rom[ 8812]='h00000000;
    rd_cycle[ 8813] = 1'b0;  wr_cycle[ 8813] = 1'b1;  addr_rom[ 8813]='h00003890;  wr_data_rom[ 8813]='h00001173;
    rd_cycle[ 8814] = 1'b0;  wr_cycle[ 8814] = 1'b1;  addr_rom[ 8814]='h00003f5c;  wr_data_rom[ 8814]='h00001613;
    rd_cycle[ 8815] = 1'b0;  wr_cycle[ 8815] = 1'b1;  addr_rom[ 8815]='h00002754;  wr_data_rom[ 8815]='h00001a54;
    rd_cycle[ 8816] = 1'b1;  wr_cycle[ 8816] = 1'b0;  addr_rom[ 8816]='h000001d4;  wr_data_rom[ 8816]='h00000000;
    rd_cycle[ 8817] = 1'b0;  wr_cycle[ 8817] = 1'b1;  addr_rom[ 8817]='h000005a0;  wr_data_rom[ 8817]='h00000b8f;
    rd_cycle[ 8818] = 1'b0;  wr_cycle[ 8818] = 1'b1;  addr_rom[ 8818]='h00003340;  wr_data_rom[ 8818]='h00003fbe;
    rd_cycle[ 8819] = 1'b1;  wr_cycle[ 8819] = 1'b0;  addr_rom[ 8819]='h00003abc;  wr_data_rom[ 8819]='h00000000;
    rd_cycle[ 8820] = 1'b1;  wr_cycle[ 8820] = 1'b0;  addr_rom[ 8820]='h000016b4;  wr_data_rom[ 8820]='h00000000;
    rd_cycle[ 8821] = 1'b1;  wr_cycle[ 8821] = 1'b0;  addr_rom[ 8821]='h000039f4;  wr_data_rom[ 8821]='h00000000;
    rd_cycle[ 8822] = 1'b0;  wr_cycle[ 8822] = 1'b1;  addr_rom[ 8822]='h00000578;  wr_data_rom[ 8822]='h000013ac;
    rd_cycle[ 8823] = 1'b0;  wr_cycle[ 8823] = 1'b1;  addr_rom[ 8823]='h00002ea4;  wr_data_rom[ 8823]='h00001053;
    rd_cycle[ 8824] = 1'b1;  wr_cycle[ 8824] = 1'b0;  addr_rom[ 8824]='h00001094;  wr_data_rom[ 8824]='h00000000;
    rd_cycle[ 8825] = 1'b1;  wr_cycle[ 8825] = 1'b0;  addr_rom[ 8825]='h0000006c;  wr_data_rom[ 8825]='h00000000;
    rd_cycle[ 8826] = 1'b1;  wr_cycle[ 8826] = 1'b0;  addr_rom[ 8826]='h00001708;  wr_data_rom[ 8826]='h00000000;
    rd_cycle[ 8827] = 1'b1;  wr_cycle[ 8827] = 1'b0;  addr_rom[ 8827]='h00002bd0;  wr_data_rom[ 8827]='h00000000;
    rd_cycle[ 8828] = 1'b0;  wr_cycle[ 8828] = 1'b1;  addr_rom[ 8828]='h000016ec;  wr_data_rom[ 8828]='h000019ce;
    rd_cycle[ 8829] = 1'b1;  wr_cycle[ 8829] = 1'b0;  addr_rom[ 8829]='h000024a0;  wr_data_rom[ 8829]='h00000000;
    rd_cycle[ 8830] = 1'b1;  wr_cycle[ 8830] = 1'b0;  addr_rom[ 8830]='h00002e6c;  wr_data_rom[ 8830]='h00000000;
    rd_cycle[ 8831] = 1'b0;  wr_cycle[ 8831] = 1'b1;  addr_rom[ 8831]='h000009e0;  wr_data_rom[ 8831]='h00000f17;
    rd_cycle[ 8832] = 1'b1;  wr_cycle[ 8832] = 1'b0;  addr_rom[ 8832]='h00003584;  wr_data_rom[ 8832]='h00000000;
    rd_cycle[ 8833] = 1'b1;  wr_cycle[ 8833] = 1'b0;  addr_rom[ 8833]='h00001234;  wr_data_rom[ 8833]='h00000000;
    rd_cycle[ 8834] = 1'b1;  wr_cycle[ 8834] = 1'b0;  addr_rom[ 8834]='h000032d0;  wr_data_rom[ 8834]='h00000000;
    rd_cycle[ 8835] = 1'b0;  wr_cycle[ 8835] = 1'b1;  addr_rom[ 8835]='h00000cf8;  wr_data_rom[ 8835]='h00003d8b;
    rd_cycle[ 8836] = 1'b1;  wr_cycle[ 8836] = 1'b0;  addr_rom[ 8836]='h00002040;  wr_data_rom[ 8836]='h00000000;
    rd_cycle[ 8837] = 1'b0;  wr_cycle[ 8837] = 1'b1;  addr_rom[ 8837]='h0000137c;  wr_data_rom[ 8837]='h000015bc;
    rd_cycle[ 8838] = 1'b1;  wr_cycle[ 8838] = 1'b0;  addr_rom[ 8838]='h00002164;  wr_data_rom[ 8838]='h00000000;
    rd_cycle[ 8839] = 1'b0;  wr_cycle[ 8839] = 1'b1;  addr_rom[ 8839]='h00002ad4;  wr_data_rom[ 8839]='h00000bc4;
    rd_cycle[ 8840] = 1'b1;  wr_cycle[ 8840] = 1'b0;  addr_rom[ 8840]='h000030bc;  wr_data_rom[ 8840]='h00000000;
    rd_cycle[ 8841] = 1'b1;  wr_cycle[ 8841] = 1'b0;  addr_rom[ 8841]='h000029c0;  wr_data_rom[ 8841]='h00000000;
    rd_cycle[ 8842] = 1'b1;  wr_cycle[ 8842] = 1'b0;  addr_rom[ 8842]='h0000042c;  wr_data_rom[ 8842]='h00000000;
    rd_cycle[ 8843] = 1'b1;  wr_cycle[ 8843] = 1'b0;  addr_rom[ 8843]='h00003124;  wr_data_rom[ 8843]='h00000000;
    rd_cycle[ 8844] = 1'b1;  wr_cycle[ 8844] = 1'b0;  addr_rom[ 8844]='h0000372c;  wr_data_rom[ 8844]='h00000000;
    rd_cycle[ 8845] = 1'b1;  wr_cycle[ 8845] = 1'b0;  addr_rom[ 8845]='h00000814;  wr_data_rom[ 8845]='h00000000;
    rd_cycle[ 8846] = 1'b1;  wr_cycle[ 8846] = 1'b0;  addr_rom[ 8846]='h00003a88;  wr_data_rom[ 8846]='h00000000;
    rd_cycle[ 8847] = 1'b0;  wr_cycle[ 8847] = 1'b1;  addr_rom[ 8847]='h00003050;  wr_data_rom[ 8847]='h00001e80;
    rd_cycle[ 8848] = 1'b0;  wr_cycle[ 8848] = 1'b1;  addr_rom[ 8848]='h00001e58;  wr_data_rom[ 8848]='h000021ef;
    rd_cycle[ 8849] = 1'b0;  wr_cycle[ 8849] = 1'b1;  addr_rom[ 8849]='h00001d70;  wr_data_rom[ 8849]='h0000185f;
    rd_cycle[ 8850] = 1'b0;  wr_cycle[ 8850] = 1'b1;  addr_rom[ 8850]='h000023ec;  wr_data_rom[ 8850]='h00002bc9;
    rd_cycle[ 8851] = 1'b1;  wr_cycle[ 8851] = 1'b0;  addr_rom[ 8851]='h00002c2c;  wr_data_rom[ 8851]='h00000000;
    rd_cycle[ 8852] = 1'b1;  wr_cycle[ 8852] = 1'b0;  addr_rom[ 8852]='h00001598;  wr_data_rom[ 8852]='h00000000;
    rd_cycle[ 8853] = 1'b0;  wr_cycle[ 8853] = 1'b1;  addr_rom[ 8853]='h0000133c;  wr_data_rom[ 8853]='h00000636;
    rd_cycle[ 8854] = 1'b0;  wr_cycle[ 8854] = 1'b1;  addr_rom[ 8854]='h00001f84;  wr_data_rom[ 8854]='h00000789;
    rd_cycle[ 8855] = 1'b0;  wr_cycle[ 8855] = 1'b1;  addr_rom[ 8855]='h0000122c;  wr_data_rom[ 8855]='h000021bf;
    rd_cycle[ 8856] = 1'b0;  wr_cycle[ 8856] = 1'b1;  addr_rom[ 8856]='h000017ac;  wr_data_rom[ 8856]='h0000168b;
    rd_cycle[ 8857] = 1'b1;  wr_cycle[ 8857] = 1'b0;  addr_rom[ 8857]='h0000167c;  wr_data_rom[ 8857]='h00000000;
    rd_cycle[ 8858] = 1'b1;  wr_cycle[ 8858] = 1'b0;  addr_rom[ 8858]='h00002a5c;  wr_data_rom[ 8858]='h00000000;
    rd_cycle[ 8859] = 1'b0;  wr_cycle[ 8859] = 1'b1;  addr_rom[ 8859]='h00002be4;  wr_data_rom[ 8859]='h000025e9;
    rd_cycle[ 8860] = 1'b0;  wr_cycle[ 8860] = 1'b1;  addr_rom[ 8860]='h00003f9c;  wr_data_rom[ 8860]='h00001065;
    rd_cycle[ 8861] = 1'b1;  wr_cycle[ 8861] = 1'b0;  addr_rom[ 8861]='h000003fc;  wr_data_rom[ 8861]='h00000000;
    rd_cycle[ 8862] = 1'b0;  wr_cycle[ 8862] = 1'b1;  addr_rom[ 8862]='h00000a54;  wr_data_rom[ 8862]='h0000090c;
    rd_cycle[ 8863] = 1'b1;  wr_cycle[ 8863] = 1'b0;  addr_rom[ 8863]='h00001d14;  wr_data_rom[ 8863]='h00000000;
    rd_cycle[ 8864] = 1'b1;  wr_cycle[ 8864] = 1'b0;  addr_rom[ 8864]='h00001520;  wr_data_rom[ 8864]='h00000000;
    rd_cycle[ 8865] = 1'b0;  wr_cycle[ 8865] = 1'b1;  addr_rom[ 8865]='h00001a4c;  wr_data_rom[ 8865]='h00000df1;
    rd_cycle[ 8866] = 1'b0;  wr_cycle[ 8866] = 1'b1;  addr_rom[ 8866]='h00001918;  wr_data_rom[ 8866]='h00001ad8;
    rd_cycle[ 8867] = 1'b0;  wr_cycle[ 8867] = 1'b1;  addr_rom[ 8867]='h00003960;  wr_data_rom[ 8867]='h00002362;
    rd_cycle[ 8868] = 1'b1;  wr_cycle[ 8868] = 1'b0;  addr_rom[ 8868]='h00003c88;  wr_data_rom[ 8868]='h00000000;
    rd_cycle[ 8869] = 1'b1;  wr_cycle[ 8869] = 1'b0;  addr_rom[ 8869]='h000027bc;  wr_data_rom[ 8869]='h00000000;
    rd_cycle[ 8870] = 1'b0;  wr_cycle[ 8870] = 1'b1;  addr_rom[ 8870]='h00001bb0;  wr_data_rom[ 8870]='h00000bb1;
    rd_cycle[ 8871] = 1'b1;  wr_cycle[ 8871] = 1'b0;  addr_rom[ 8871]='h0000056c;  wr_data_rom[ 8871]='h00000000;
    rd_cycle[ 8872] = 1'b1;  wr_cycle[ 8872] = 1'b0;  addr_rom[ 8872]='h00002c8c;  wr_data_rom[ 8872]='h00000000;
    rd_cycle[ 8873] = 1'b0;  wr_cycle[ 8873] = 1'b1;  addr_rom[ 8873]='h000015c0;  wr_data_rom[ 8873]='h0000215b;
    rd_cycle[ 8874] = 1'b1;  wr_cycle[ 8874] = 1'b0;  addr_rom[ 8874]='h00003700;  wr_data_rom[ 8874]='h00000000;
    rd_cycle[ 8875] = 1'b1;  wr_cycle[ 8875] = 1'b0;  addr_rom[ 8875]='h00001130;  wr_data_rom[ 8875]='h00000000;
    rd_cycle[ 8876] = 1'b0;  wr_cycle[ 8876] = 1'b1;  addr_rom[ 8876]='h00001b00;  wr_data_rom[ 8876]='h00000992;
    rd_cycle[ 8877] = 1'b0;  wr_cycle[ 8877] = 1'b1;  addr_rom[ 8877]='h000011a8;  wr_data_rom[ 8877]='h0000193c;
    rd_cycle[ 8878] = 1'b0;  wr_cycle[ 8878] = 1'b1;  addr_rom[ 8878]='h00003f0c;  wr_data_rom[ 8878]='h00002e45;
    rd_cycle[ 8879] = 1'b0;  wr_cycle[ 8879] = 1'b1;  addr_rom[ 8879]='h00002c6c;  wr_data_rom[ 8879]='h00002f53;
    rd_cycle[ 8880] = 1'b0;  wr_cycle[ 8880] = 1'b1;  addr_rom[ 8880]='h000016f4;  wr_data_rom[ 8880]='h000003ae;
    rd_cycle[ 8881] = 1'b1;  wr_cycle[ 8881] = 1'b0;  addr_rom[ 8881]='h00003100;  wr_data_rom[ 8881]='h00000000;
    rd_cycle[ 8882] = 1'b1;  wr_cycle[ 8882] = 1'b0;  addr_rom[ 8882]='h000030b8;  wr_data_rom[ 8882]='h00000000;
    rd_cycle[ 8883] = 1'b0;  wr_cycle[ 8883] = 1'b1;  addr_rom[ 8883]='h00002a64;  wr_data_rom[ 8883]='h00001bd2;
    rd_cycle[ 8884] = 1'b0;  wr_cycle[ 8884] = 1'b1;  addr_rom[ 8884]='h00003ab0;  wr_data_rom[ 8884]='h00002dd0;
    rd_cycle[ 8885] = 1'b0;  wr_cycle[ 8885] = 1'b1;  addr_rom[ 8885]='h00001544;  wr_data_rom[ 8885]='h000004ec;
    rd_cycle[ 8886] = 1'b1;  wr_cycle[ 8886] = 1'b0;  addr_rom[ 8886]='h00002124;  wr_data_rom[ 8886]='h00000000;
    rd_cycle[ 8887] = 1'b0;  wr_cycle[ 8887] = 1'b1;  addr_rom[ 8887]='h00001950;  wr_data_rom[ 8887]='h000023ab;
    rd_cycle[ 8888] = 1'b0;  wr_cycle[ 8888] = 1'b1;  addr_rom[ 8888]='h000030f8;  wr_data_rom[ 8888]='h00000783;
    rd_cycle[ 8889] = 1'b1;  wr_cycle[ 8889] = 1'b0;  addr_rom[ 8889]='h00002828;  wr_data_rom[ 8889]='h00000000;
    rd_cycle[ 8890] = 1'b0;  wr_cycle[ 8890] = 1'b1;  addr_rom[ 8890]='h00002530;  wr_data_rom[ 8890]='h000002e1;
    rd_cycle[ 8891] = 1'b1;  wr_cycle[ 8891] = 1'b0;  addr_rom[ 8891]='h00001b50;  wr_data_rom[ 8891]='h00000000;
    rd_cycle[ 8892] = 1'b1;  wr_cycle[ 8892] = 1'b0;  addr_rom[ 8892]='h000023b8;  wr_data_rom[ 8892]='h00000000;
    rd_cycle[ 8893] = 1'b1;  wr_cycle[ 8893] = 1'b0;  addr_rom[ 8893]='h00003770;  wr_data_rom[ 8893]='h00000000;
    rd_cycle[ 8894] = 1'b0;  wr_cycle[ 8894] = 1'b1;  addr_rom[ 8894]='h0000006c;  wr_data_rom[ 8894]='h000039de;
    rd_cycle[ 8895] = 1'b0;  wr_cycle[ 8895] = 1'b1;  addr_rom[ 8895]='h00000f28;  wr_data_rom[ 8895]='h00002f88;
    rd_cycle[ 8896] = 1'b0;  wr_cycle[ 8896] = 1'b1;  addr_rom[ 8896]='h00002560;  wr_data_rom[ 8896]='h00001eff;
    rd_cycle[ 8897] = 1'b1;  wr_cycle[ 8897] = 1'b0;  addr_rom[ 8897]='h00003b10;  wr_data_rom[ 8897]='h00000000;
    rd_cycle[ 8898] = 1'b1;  wr_cycle[ 8898] = 1'b0;  addr_rom[ 8898]='h00002908;  wr_data_rom[ 8898]='h00000000;
    rd_cycle[ 8899] = 1'b1;  wr_cycle[ 8899] = 1'b0;  addr_rom[ 8899]='h00000080;  wr_data_rom[ 8899]='h00000000;
    rd_cycle[ 8900] = 1'b0;  wr_cycle[ 8900] = 1'b1;  addr_rom[ 8900]='h00002e9c;  wr_data_rom[ 8900]='h00003c88;
    rd_cycle[ 8901] = 1'b0;  wr_cycle[ 8901] = 1'b1;  addr_rom[ 8901]='h000014d0;  wr_data_rom[ 8901]='h0000099a;
    rd_cycle[ 8902] = 1'b1;  wr_cycle[ 8902] = 1'b0;  addr_rom[ 8902]='h00003640;  wr_data_rom[ 8902]='h00000000;
    rd_cycle[ 8903] = 1'b1;  wr_cycle[ 8903] = 1'b0;  addr_rom[ 8903]='h00001c2c;  wr_data_rom[ 8903]='h00000000;
    rd_cycle[ 8904] = 1'b0;  wr_cycle[ 8904] = 1'b1;  addr_rom[ 8904]='h0000135c;  wr_data_rom[ 8904]='h00000023;
    rd_cycle[ 8905] = 1'b0;  wr_cycle[ 8905] = 1'b1;  addr_rom[ 8905]='h00001e94;  wr_data_rom[ 8905]='h00000170;
    rd_cycle[ 8906] = 1'b1;  wr_cycle[ 8906] = 1'b0;  addr_rom[ 8906]='h0000246c;  wr_data_rom[ 8906]='h00000000;
    rd_cycle[ 8907] = 1'b0;  wr_cycle[ 8907] = 1'b1;  addr_rom[ 8907]='h00003c7c;  wr_data_rom[ 8907]='h00002db8;
    rd_cycle[ 8908] = 1'b1;  wr_cycle[ 8908] = 1'b0;  addr_rom[ 8908]='h0000133c;  wr_data_rom[ 8908]='h00000000;
    rd_cycle[ 8909] = 1'b1;  wr_cycle[ 8909] = 1'b0;  addr_rom[ 8909]='h000007c8;  wr_data_rom[ 8909]='h00000000;
    rd_cycle[ 8910] = 1'b0;  wr_cycle[ 8910] = 1'b1;  addr_rom[ 8910]='h000034b4;  wr_data_rom[ 8910]='h00003937;
    rd_cycle[ 8911] = 1'b1;  wr_cycle[ 8911] = 1'b0;  addr_rom[ 8911]='h000037f0;  wr_data_rom[ 8911]='h00000000;
    rd_cycle[ 8912] = 1'b0;  wr_cycle[ 8912] = 1'b1;  addr_rom[ 8912]='h00001950;  wr_data_rom[ 8912]='h00002337;
    rd_cycle[ 8913] = 1'b0;  wr_cycle[ 8913] = 1'b1;  addr_rom[ 8913]='h0000284c;  wr_data_rom[ 8913]='h00000c5d;
    rd_cycle[ 8914] = 1'b1;  wr_cycle[ 8914] = 1'b0;  addr_rom[ 8914]='h00001040;  wr_data_rom[ 8914]='h00000000;
    rd_cycle[ 8915] = 1'b0;  wr_cycle[ 8915] = 1'b1;  addr_rom[ 8915]='h00001fb8;  wr_data_rom[ 8915]='h000036a5;
    rd_cycle[ 8916] = 1'b0;  wr_cycle[ 8916] = 1'b1;  addr_rom[ 8916]='h00003aa0;  wr_data_rom[ 8916]='h0000341a;
    rd_cycle[ 8917] = 1'b0;  wr_cycle[ 8917] = 1'b1;  addr_rom[ 8917]='h00003dd4;  wr_data_rom[ 8917]='h00002ed2;
    rd_cycle[ 8918] = 1'b0;  wr_cycle[ 8918] = 1'b1;  addr_rom[ 8918]='h0000162c;  wr_data_rom[ 8918]='h000027c3;
    rd_cycle[ 8919] = 1'b1;  wr_cycle[ 8919] = 1'b0;  addr_rom[ 8919]='h00003488;  wr_data_rom[ 8919]='h00000000;
    rd_cycle[ 8920] = 1'b1;  wr_cycle[ 8920] = 1'b0;  addr_rom[ 8920]='h00003ba4;  wr_data_rom[ 8920]='h00000000;
    rd_cycle[ 8921] = 1'b1;  wr_cycle[ 8921] = 1'b0;  addr_rom[ 8921]='h00002790;  wr_data_rom[ 8921]='h00000000;
    rd_cycle[ 8922] = 1'b1;  wr_cycle[ 8922] = 1'b0;  addr_rom[ 8922]='h00003ca8;  wr_data_rom[ 8922]='h00000000;
    rd_cycle[ 8923] = 1'b1;  wr_cycle[ 8923] = 1'b0;  addr_rom[ 8923]='h000028c0;  wr_data_rom[ 8923]='h00000000;
    rd_cycle[ 8924] = 1'b0;  wr_cycle[ 8924] = 1'b1;  addr_rom[ 8924]='h00000d08;  wr_data_rom[ 8924]='h00000cbc;
    rd_cycle[ 8925] = 1'b0;  wr_cycle[ 8925] = 1'b1;  addr_rom[ 8925]='h00000ce8;  wr_data_rom[ 8925]='h000032ff;
    rd_cycle[ 8926] = 1'b1;  wr_cycle[ 8926] = 1'b0;  addr_rom[ 8926]='h000001f4;  wr_data_rom[ 8926]='h00000000;
    rd_cycle[ 8927] = 1'b1;  wr_cycle[ 8927] = 1'b0;  addr_rom[ 8927]='h000018b4;  wr_data_rom[ 8927]='h00000000;
    rd_cycle[ 8928] = 1'b0;  wr_cycle[ 8928] = 1'b1;  addr_rom[ 8928]='h00002118;  wr_data_rom[ 8928]='h0000059a;
    rd_cycle[ 8929] = 1'b0;  wr_cycle[ 8929] = 1'b1;  addr_rom[ 8929]='h00002320;  wr_data_rom[ 8929]='h000000f7;
    rd_cycle[ 8930] = 1'b0;  wr_cycle[ 8930] = 1'b1;  addr_rom[ 8930]='h00000ff4;  wr_data_rom[ 8930]='h000015df;
    rd_cycle[ 8931] = 1'b0;  wr_cycle[ 8931] = 1'b1;  addr_rom[ 8931]='h000027fc;  wr_data_rom[ 8931]='h00003bbb;
    rd_cycle[ 8932] = 1'b0;  wr_cycle[ 8932] = 1'b1;  addr_rom[ 8932]='h00003e30;  wr_data_rom[ 8932]='h00002008;
    rd_cycle[ 8933] = 1'b0;  wr_cycle[ 8933] = 1'b1;  addr_rom[ 8933]='h00000ad0;  wr_data_rom[ 8933]='h000031fd;
    rd_cycle[ 8934] = 1'b0;  wr_cycle[ 8934] = 1'b1;  addr_rom[ 8934]='h000018dc;  wr_data_rom[ 8934]='h00003af4;
    rd_cycle[ 8935] = 1'b1;  wr_cycle[ 8935] = 1'b0;  addr_rom[ 8935]='h00003d64;  wr_data_rom[ 8935]='h00000000;
    rd_cycle[ 8936] = 1'b0;  wr_cycle[ 8936] = 1'b1;  addr_rom[ 8936]='h000003a8;  wr_data_rom[ 8936]='h000033d4;
    rd_cycle[ 8937] = 1'b0;  wr_cycle[ 8937] = 1'b1;  addr_rom[ 8937]='h000015ec;  wr_data_rom[ 8937]='h00002960;
    rd_cycle[ 8938] = 1'b0;  wr_cycle[ 8938] = 1'b1;  addr_rom[ 8938]='h0000115c;  wr_data_rom[ 8938]='h000029db;
    rd_cycle[ 8939] = 1'b1;  wr_cycle[ 8939] = 1'b0;  addr_rom[ 8939]='h00002bd0;  wr_data_rom[ 8939]='h00000000;
    rd_cycle[ 8940] = 1'b1;  wr_cycle[ 8940] = 1'b0;  addr_rom[ 8940]='h0000215c;  wr_data_rom[ 8940]='h00000000;
    rd_cycle[ 8941] = 1'b0;  wr_cycle[ 8941] = 1'b1;  addr_rom[ 8941]='h000033c8;  wr_data_rom[ 8941]='h000015c4;
    rd_cycle[ 8942] = 1'b0;  wr_cycle[ 8942] = 1'b1;  addr_rom[ 8942]='h000014e4;  wr_data_rom[ 8942]='h00002c3a;
    rd_cycle[ 8943] = 1'b0;  wr_cycle[ 8943] = 1'b1;  addr_rom[ 8943]='h0000245c;  wr_data_rom[ 8943]='h00002051;
    rd_cycle[ 8944] = 1'b0;  wr_cycle[ 8944] = 1'b1;  addr_rom[ 8944]='h000002e4;  wr_data_rom[ 8944]='h000015a1;
    rd_cycle[ 8945] = 1'b1;  wr_cycle[ 8945] = 1'b0;  addr_rom[ 8945]='h00003290;  wr_data_rom[ 8945]='h00000000;
    rd_cycle[ 8946] = 1'b1;  wr_cycle[ 8946] = 1'b0;  addr_rom[ 8946]='h00001d28;  wr_data_rom[ 8946]='h00000000;
    rd_cycle[ 8947] = 1'b0;  wr_cycle[ 8947] = 1'b1;  addr_rom[ 8947]='h00002c7c;  wr_data_rom[ 8947]='h000002ad;
    rd_cycle[ 8948] = 1'b1;  wr_cycle[ 8948] = 1'b0;  addr_rom[ 8948]='h00002a4c;  wr_data_rom[ 8948]='h00000000;
    rd_cycle[ 8949] = 1'b0;  wr_cycle[ 8949] = 1'b1;  addr_rom[ 8949]='h0000166c;  wr_data_rom[ 8949]='h000015bb;
    rd_cycle[ 8950] = 1'b0;  wr_cycle[ 8950] = 1'b1;  addr_rom[ 8950]='h00002454;  wr_data_rom[ 8950]='h00003d6d;
    rd_cycle[ 8951] = 1'b1;  wr_cycle[ 8951] = 1'b0;  addr_rom[ 8951]='h0000383c;  wr_data_rom[ 8951]='h00000000;
    rd_cycle[ 8952] = 1'b0;  wr_cycle[ 8952] = 1'b1;  addr_rom[ 8952]='h0000311c;  wr_data_rom[ 8952]='h00001a57;
    rd_cycle[ 8953] = 1'b1;  wr_cycle[ 8953] = 1'b0;  addr_rom[ 8953]='h000034a8;  wr_data_rom[ 8953]='h00000000;
    rd_cycle[ 8954] = 1'b0;  wr_cycle[ 8954] = 1'b1;  addr_rom[ 8954]='h000027e4;  wr_data_rom[ 8954]='h00002b38;
    rd_cycle[ 8955] = 1'b0;  wr_cycle[ 8955] = 1'b1;  addr_rom[ 8955]='h00003b5c;  wr_data_rom[ 8955]='h00000789;
    rd_cycle[ 8956] = 1'b0;  wr_cycle[ 8956] = 1'b1;  addr_rom[ 8956]='h0000346c;  wr_data_rom[ 8956]='h00003660;
    rd_cycle[ 8957] = 1'b1;  wr_cycle[ 8957] = 1'b0;  addr_rom[ 8957]='h00000f88;  wr_data_rom[ 8957]='h00000000;
    rd_cycle[ 8958] = 1'b0;  wr_cycle[ 8958] = 1'b1;  addr_rom[ 8958]='h000007a8;  wr_data_rom[ 8958]='h000017b3;
    rd_cycle[ 8959] = 1'b0;  wr_cycle[ 8959] = 1'b1;  addr_rom[ 8959]='h00003694;  wr_data_rom[ 8959]='h00001614;
    rd_cycle[ 8960] = 1'b1;  wr_cycle[ 8960] = 1'b0;  addr_rom[ 8960]='h000028b4;  wr_data_rom[ 8960]='h00000000;
    rd_cycle[ 8961] = 1'b0;  wr_cycle[ 8961] = 1'b1;  addr_rom[ 8961]='h0000327c;  wr_data_rom[ 8961]='h00003b0f;
    rd_cycle[ 8962] = 1'b1;  wr_cycle[ 8962] = 1'b0;  addr_rom[ 8962]='h0000286c;  wr_data_rom[ 8962]='h00000000;
    rd_cycle[ 8963] = 1'b1;  wr_cycle[ 8963] = 1'b0;  addr_rom[ 8963]='h00001ea8;  wr_data_rom[ 8963]='h00000000;
    rd_cycle[ 8964] = 1'b1;  wr_cycle[ 8964] = 1'b0;  addr_rom[ 8964]='h00001764;  wr_data_rom[ 8964]='h00000000;
    rd_cycle[ 8965] = 1'b1;  wr_cycle[ 8965] = 1'b0;  addr_rom[ 8965]='h00001ab8;  wr_data_rom[ 8965]='h00000000;
    rd_cycle[ 8966] = 1'b1;  wr_cycle[ 8966] = 1'b0;  addr_rom[ 8966]='h0000222c;  wr_data_rom[ 8966]='h00000000;
    rd_cycle[ 8967] = 1'b0;  wr_cycle[ 8967] = 1'b1;  addr_rom[ 8967]='h000027e4;  wr_data_rom[ 8967]='h00001a9f;
    rd_cycle[ 8968] = 1'b0;  wr_cycle[ 8968] = 1'b1;  addr_rom[ 8968]='h0000134c;  wr_data_rom[ 8968]='h00001697;
    rd_cycle[ 8969] = 1'b1;  wr_cycle[ 8969] = 1'b0;  addr_rom[ 8969]='h000008dc;  wr_data_rom[ 8969]='h00000000;
    rd_cycle[ 8970] = 1'b1;  wr_cycle[ 8970] = 1'b0;  addr_rom[ 8970]='h000028ec;  wr_data_rom[ 8970]='h00000000;
    rd_cycle[ 8971] = 1'b1;  wr_cycle[ 8971] = 1'b0;  addr_rom[ 8971]='h00002bcc;  wr_data_rom[ 8971]='h00000000;
    rd_cycle[ 8972] = 1'b0;  wr_cycle[ 8972] = 1'b1;  addr_rom[ 8972]='h00001e0c;  wr_data_rom[ 8972]='h00000d0d;
    rd_cycle[ 8973] = 1'b0;  wr_cycle[ 8973] = 1'b1;  addr_rom[ 8973]='h00000fac;  wr_data_rom[ 8973]='h00001aaa;
    rd_cycle[ 8974] = 1'b1;  wr_cycle[ 8974] = 1'b0;  addr_rom[ 8974]='h00003cd0;  wr_data_rom[ 8974]='h00000000;
    rd_cycle[ 8975] = 1'b0;  wr_cycle[ 8975] = 1'b1;  addr_rom[ 8975]='h00000740;  wr_data_rom[ 8975]='h00001229;
    rd_cycle[ 8976] = 1'b0;  wr_cycle[ 8976] = 1'b1;  addr_rom[ 8976]='h000039e4;  wr_data_rom[ 8976]='h000020aa;
    rd_cycle[ 8977] = 1'b0;  wr_cycle[ 8977] = 1'b1;  addr_rom[ 8977]='h00000c58;  wr_data_rom[ 8977]='h0000114e;
    rd_cycle[ 8978] = 1'b0;  wr_cycle[ 8978] = 1'b1;  addr_rom[ 8978]='h000000b8;  wr_data_rom[ 8978]='h0000272b;
    rd_cycle[ 8979] = 1'b1;  wr_cycle[ 8979] = 1'b0;  addr_rom[ 8979]='h00003990;  wr_data_rom[ 8979]='h00000000;
    rd_cycle[ 8980] = 1'b0;  wr_cycle[ 8980] = 1'b1;  addr_rom[ 8980]='h000032cc;  wr_data_rom[ 8980]='h00003e85;
    rd_cycle[ 8981] = 1'b0;  wr_cycle[ 8981] = 1'b1;  addr_rom[ 8981]='h00000ddc;  wr_data_rom[ 8981]='h00000e1c;
    rd_cycle[ 8982] = 1'b0;  wr_cycle[ 8982] = 1'b1;  addr_rom[ 8982]='h00001034;  wr_data_rom[ 8982]='h000011fb;
    rd_cycle[ 8983] = 1'b0;  wr_cycle[ 8983] = 1'b1;  addr_rom[ 8983]='h00002cc8;  wr_data_rom[ 8983]='h000010aa;
    rd_cycle[ 8984] = 1'b0;  wr_cycle[ 8984] = 1'b1;  addr_rom[ 8984]='h00002a94;  wr_data_rom[ 8984]='h000007ad;
    rd_cycle[ 8985] = 1'b1;  wr_cycle[ 8985] = 1'b0;  addr_rom[ 8985]='h00002abc;  wr_data_rom[ 8985]='h00000000;
    rd_cycle[ 8986] = 1'b0;  wr_cycle[ 8986] = 1'b1;  addr_rom[ 8986]='h00003a64;  wr_data_rom[ 8986]='h00003636;
    rd_cycle[ 8987] = 1'b1;  wr_cycle[ 8987] = 1'b0;  addr_rom[ 8987]='h00000c10;  wr_data_rom[ 8987]='h00000000;
    rd_cycle[ 8988] = 1'b0;  wr_cycle[ 8988] = 1'b1;  addr_rom[ 8988]='h00003d74;  wr_data_rom[ 8988]='h00000263;
    rd_cycle[ 8989] = 1'b0;  wr_cycle[ 8989] = 1'b1;  addr_rom[ 8989]='h000009f0;  wr_data_rom[ 8989]='h00000d4e;
    rd_cycle[ 8990] = 1'b1;  wr_cycle[ 8990] = 1'b0;  addr_rom[ 8990]='h000018e4;  wr_data_rom[ 8990]='h00000000;
    rd_cycle[ 8991] = 1'b1;  wr_cycle[ 8991] = 1'b0;  addr_rom[ 8991]='h00000468;  wr_data_rom[ 8991]='h00000000;
    rd_cycle[ 8992] = 1'b0;  wr_cycle[ 8992] = 1'b1;  addr_rom[ 8992]='h00000dec;  wr_data_rom[ 8992]='h000010c1;
    rd_cycle[ 8993] = 1'b0;  wr_cycle[ 8993] = 1'b1;  addr_rom[ 8993]='h0000316c;  wr_data_rom[ 8993]='h000001b9;
    rd_cycle[ 8994] = 1'b1;  wr_cycle[ 8994] = 1'b0;  addr_rom[ 8994]='h000027c8;  wr_data_rom[ 8994]='h00000000;
    rd_cycle[ 8995] = 1'b1;  wr_cycle[ 8995] = 1'b0;  addr_rom[ 8995]='h00001da8;  wr_data_rom[ 8995]='h00000000;
    rd_cycle[ 8996] = 1'b1;  wr_cycle[ 8996] = 1'b0;  addr_rom[ 8996]='h00001d44;  wr_data_rom[ 8996]='h00000000;
    rd_cycle[ 8997] = 1'b1;  wr_cycle[ 8997] = 1'b0;  addr_rom[ 8997]='h000033b0;  wr_data_rom[ 8997]='h00000000;
    rd_cycle[ 8998] = 1'b1;  wr_cycle[ 8998] = 1'b0;  addr_rom[ 8998]='h000016ac;  wr_data_rom[ 8998]='h00000000;
    rd_cycle[ 8999] = 1'b1;  wr_cycle[ 8999] = 1'b0;  addr_rom[ 8999]='h00000a00;  wr_data_rom[ 8999]='h00000000;
    rd_cycle[ 9000] = 1'b0;  wr_cycle[ 9000] = 1'b1;  addr_rom[ 9000]='h00002498;  wr_data_rom[ 9000]='h00003fad;
    rd_cycle[ 9001] = 1'b1;  wr_cycle[ 9001] = 1'b0;  addr_rom[ 9001]='h00000acc;  wr_data_rom[ 9001]='h00000000;
    rd_cycle[ 9002] = 1'b1;  wr_cycle[ 9002] = 1'b0;  addr_rom[ 9002]='h00002ba0;  wr_data_rom[ 9002]='h00000000;
    rd_cycle[ 9003] = 1'b0;  wr_cycle[ 9003] = 1'b1;  addr_rom[ 9003]='h000019d4;  wr_data_rom[ 9003]='h00003fb8;
    rd_cycle[ 9004] = 1'b0;  wr_cycle[ 9004] = 1'b1;  addr_rom[ 9004]='h00001efc;  wr_data_rom[ 9004]='h0000060a;
    rd_cycle[ 9005] = 1'b0;  wr_cycle[ 9005] = 1'b1;  addr_rom[ 9005]='h000032f8;  wr_data_rom[ 9005]='h000000fd;
    rd_cycle[ 9006] = 1'b1;  wr_cycle[ 9006] = 1'b0;  addr_rom[ 9006]='h00002c88;  wr_data_rom[ 9006]='h00000000;
    rd_cycle[ 9007] = 1'b1;  wr_cycle[ 9007] = 1'b0;  addr_rom[ 9007]='h00002108;  wr_data_rom[ 9007]='h00000000;
    rd_cycle[ 9008] = 1'b0;  wr_cycle[ 9008] = 1'b1;  addr_rom[ 9008]='h00002134;  wr_data_rom[ 9008]='h00002e7c;
    rd_cycle[ 9009] = 1'b1;  wr_cycle[ 9009] = 1'b0;  addr_rom[ 9009]='h00000f0c;  wr_data_rom[ 9009]='h00000000;
    rd_cycle[ 9010] = 1'b1;  wr_cycle[ 9010] = 1'b0;  addr_rom[ 9010]='h00001da0;  wr_data_rom[ 9010]='h00000000;
    rd_cycle[ 9011] = 1'b1;  wr_cycle[ 9011] = 1'b0;  addr_rom[ 9011]='h00003524;  wr_data_rom[ 9011]='h00000000;
    rd_cycle[ 9012] = 1'b0;  wr_cycle[ 9012] = 1'b1;  addr_rom[ 9012]='h00000afc;  wr_data_rom[ 9012]='h00002431;
    rd_cycle[ 9013] = 1'b0;  wr_cycle[ 9013] = 1'b1;  addr_rom[ 9013]='h00001c48;  wr_data_rom[ 9013]='h00000c3a;
    rd_cycle[ 9014] = 1'b0;  wr_cycle[ 9014] = 1'b1;  addr_rom[ 9014]='h0000122c;  wr_data_rom[ 9014]='h00002f41;
    rd_cycle[ 9015] = 1'b1;  wr_cycle[ 9015] = 1'b0;  addr_rom[ 9015]='h0000329c;  wr_data_rom[ 9015]='h00000000;
    rd_cycle[ 9016] = 1'b0;  wr_cycle[ 9016] = 1'b1;  addr_rom[ 9016]='h00000d50;  wr_data_rom[ 9016]='h000030fb;
    rd_cycle[ 9017] = 1'b1;  wr_cycle[ 9017] = 1'b0;  addr_rom[ 9017]='h000025c0;  wr_data_rom[ 9017]='h00000000;
    rd_cycle[ 9018] = 1'b0;  wr_cycle[ 9018] = 1'b1;  addr_rom[ 9018]='h00003d48;  wr_data_rom[ 9018]='h00000323;
    rd_cycle[ 9019] = 1'b0;  wr_cycle[ 9019] = 1'b1;  addr_rom[ 9019]='h00002168;  wr_data_rom[ 9019]='h00002c20;
    rd_cycle[ 9020] = 1'b0;  wr_cycle[ 9020] = 1'b1;  addr_rom[ 9020]='h00002a78;  wr_data_rom[ 9020]='h00003f28;
    rd_cycle[ 9021] = 1'b0;  wr_cycle[ 9021] = 1'b1;  addr_rom[ 9021]='h0000332c;  wr_data_rom[ 9021]='h000039ae;
    rd_cycle[ 9022] = 1'b0;  wr_cycle[ 9022] = 1'b1;  addr_rom[ 9022]='h00000aa8;  wr_data_rom[ 9022]='h00003789;
    rd_cycle[ 9023] = 1'b1;  wr_cycle[ 9023] = 1'b0;  addr_rom[ 9023]='h00003508;  wr_data_rom[ 9023]='h00000000;
    rd_cycle[ 9024] = 1'b1;  wr_cycle[ 9024] = 1'b0;  addr_rom[ 9024]='h00002c7c;  wr_data_rom[ 9024]='h00000000;
    rd_cycle[ 9025] = 1'b1;  wr_cycle[ 9025] = 1'b0;  addr_rom[ 9025]='h00001278;  wr_data_rom[ 9025]='h00000000;
    rd_cycle[ 9026] = 1'b1;  wr_cycle[ 9026] = 1'b0;  addr_rom[ 9026]='h00002508;  wr_data_rom[ 9026]='h00000000;
    rd_cycle[ 9027] = 1'b0;  wr_cycle[ 9027] = 1'b1;  addr_rom[ 9027]='h000026e0;  wr_data_rom[ 9027]='h00003f70;
    rd_cycle[ 9028] = 1'b1;  wr_cycle[ 9028] = 1'b0;  addr_rom[ 9028]='h00001da0;  wr_data_rom[ 9028]='h00000000;
    rd_cycle[ 9029] = 1'b0;  wr_cycle[ 9029] = 1'b1;  addr_rom[ 9029]='h00002da8;  wr_data_rom[ 9029]='h000019db;
    rd_cycle[ 9030] = 1'b0;  wr_cycle[ 9030] = 1'b1;  addr_rom[ 9030]='h0000334c;  wr_data_rom[ 9030]='h00000b3f;
    rd_cycle[ 9031] = 1'b0;  wr_cycle[ 9031] = 1'b1;  addr_rom[ 9031]='h0000209c;  wr_data_rom[ 9031]='h00002851;
    rd_cycle[ 9032] = 1'b0;  wr_cycle[ 9032] = 1'b1;  addr_rom[ 9032]='h00000388;  wr_data_rom[ 9032]='h00001bed;
    rd_cycle[ 9033] = 1'b0;  wr_cycle[ 9033] = 1'b1;  addr_rom[ 9033]='h00002d10;  wr_data_rom[ 9033]='h00000d3b;
    rd_cycle[ 9034] = 1'b0;  wr_cycle[ 9034] = 1'b1;  addr_rom[ 9034]='h00002f5c;  wr_data_rom[ 9034]='h0000023a;
    rd_cycle[ 9035] = 1'b0;  wr_cycle[ 9035] = 1'b1;  addr_rom[ 9035]='h00002c7c;  wr_data_rom[ 9035]='h0000231d;
    rd_cycle[ 9036] = 1'b0;  wr_cycle[ 9036] = 1'b1;  addr_rom[ 9036]='h0000370c;  wr_data_rom[ 9036]='h0000291b;
    rd_cycle[ 9037] = 1'b0;  wr_cycle[ 9037] = 1'b1;  addr_rom[ 9037]='h00002ca8;  wr_data_rom[ 9037]='h00002e1c;
    rd_cycle[ 9038] = 1'b1;  wr_cycle[ 9038] = 1'b0;  addr_rom[ 9038]='h00000ea4;  wr_data_rom[ 9038]='h00000000;
    rd_cycle[ 9039] = 1'b0;  wr_cycle[ 9039] = 1'b1;  addr_rom[ 9039]='h00001da0;  wr_data_rom[ 9039]='h0000355c;
    rd_cycle[ 9040] = 1'b1;  wr_cycle[ 9040] = 1'b0;  addr_rom[ 9040]='h00000c04;  wr_data_rom[ 9040]='h00000000;
    rd_cycle[ 9041] = 1'b0;  wr_cycle[ 9041] = 1'b1;  addr_rom[ 9041]='h00001138;  wr_data_rom[ 9041]='h00002d68;
    rd_cycle[ 9042] = 1'b1;  wr_cycle[ 9042] = 1'b0;  addr_rom[ 9042]='h00002418;  wr_data_rom[ 9042]='h00000000;
    rd_cycle[ 9043] = 1'b0;  wr_cycle[ 9043] = 1'b1;  addr_rom[ 9043]='h00003898;  wr_data_rom[ 9043]='h0000370f;
    rd_cycle[ 9044] = 1'b1;  wr_cycle[ 9044] = 1'b0;  addr_rom[ 9044]='h00002f98;  wr_data_rom[ 9044]='h00000000;
    rd_cycle[ 9045] = 1'b1;  wr_cycle[ 9045] = 1'b0;  addr_rom[ 9045]='h00003098;  wr_data_rom[ 9045]='h00000000;
    rd_cycle[ 9046] = 1'b1;  wr_cycle[ 9046] = 1'b0;  addr_rom[ 9046]='h000002a0;  wr_data_rom[ 9046]='h00000000;
    rd_cycle[ 9047] = 1'b0;  wr_cycle[ 9047] = 1'b1;  addr_rom[ 9047]='h00003b5c;  wr_data_rom[ 9047]='h0000166f;
    rd_cycle[ 9048] = 1'b0;  wr_cycle[ 9048] = 1'b1;  addr_rom[ 9048]='h00001be4;  wr_data_rom[ 9048]='h0000374b;
    rd_cycle[ 9049] = 1'b1;  wr_cycle[ 9049] = 1'b0;  addr_rom[ 9049]='h00001e78;  wr_data_rom[ 9049]='h00000000;
    rd_cycle[ 9050] = 1'b0;  wr_cycle[ 9050] = 1'b1;  addr_rom[ 9050]='h0000298c;  wr_data_rom[ 9050]='h000005a3;
    rd_cycle[ 9051] = 1'b1;  wr_cycle[ 9051] = 1'b0;  addr_rom[ 9051]='h00001ba8;  wr_data_rom[ 9051]='h00000000;
    rd_cycle[ 9052] = 1'b1;  wr_cycle[ 9052] = 1'b0;  addr_rom[ 9052]='h00002040;  wr_data_rom[ 9052]='h00000000;
    rd_cycle[ 9053] = 1'b1;  wr_cycle[ 9053] = 1'b0;  addr_rom[ 9053]='h00002380;  wr_data_rom[ 9053]='h00000000;
    rd_cycle[ 9054] = 1'b1;  wr_cycle[ 9054] = 1'b0;  addr_rom[ 9054]='h000037b4;  wr_data_rom[ 9054]='h00000000;
    rd_cycle[ 9055] = 1'b0;  wr_cycle[ 9055] = 1'b1;  addr_rom[ 9055]='h00002f80;  wr_data_rom[ 9055]='h00002b3a;
    rd_cycle[ 9056] = 1'b0;  wr_cycle[ 9056] = 1'b1;  addr_rom[ 9056]='h00002b98;  wr_data_rom[ 9056]='h000011b4;
    rd_cycle[ 9057] = 1'b1;  wr_cycle[ 9057] = 1'b0;  addr_rom[ 9057]='h000004b4;  wr_data_rom[ 9057]='h00000000;
    rd_cycle[ 9058] = 1'b0;  wr_cycle[ 9058] = 1'b1;  addr_rom[ 9058]='h00003708;  wr_data_rom[ 9058]='h00001c9f;
    rd_cycle[ 9059] = 1'b0;  wr_cycle[ 9059] = 1'b1;  addr_rom[ 9059]='h00000744;  wr_data_rom[ 9059]='h00000291;
    rd_cycle[ 9060] = 1'b0;  wr_cycle[ 9060] = 1'b1;  addr_rom[ 9060]='h000037c8;  wr_data_rom[ 9060]='h00001b24;
    rd_cycle[ 9061] = 1'b1;  wr_cycle[ 9061] = 1'b0;  addr_rom[ 9061]='h00000858;  wr_data_rom[ 9061]='h00000000;
    rd_cycle[ 9062] = 1'b0;  wr_cycle[ 9062] = 1'b1;  addr_rom[ 9062]='h00003418;  wr_data_rom[ 9062]='h000002d1;
    rd_cycle[ 9063] = 1'b1;  wr_cycle[ 9063] = 1'b0;  addr_rom[ 9063]='h0000136c;  wr_data_rom[ 9063]='h00000000;
    rd_cycle[ 9064] = 1'b1;  wr_cycle[ 9064] = 1'b0;  addr_rom[ 9064]='h00000b30;  wr_data_rom[ 9064]='h00000000;
    rd_cycle[ 9065] = 1'b1;  wr_cycle[ 9065] = 1'b0;  addr_rom[ 9065]='h000015d0;  wr_data_rom[ 9065]='h00000000;
    rd_cycle[ 9066] = 1'b1;  wr_cycle[ 9066] = 1'b0;  addr_rom[ 9066]='h000012f8;  wr_data_rom[ 9066]='h00000000;
    rd_cycle[ 9067] = 1'b1;  wr_cycle[ 9067] = 1'b0;  addr_rom[ 9067]='h0000115c;  wr_data_rom[ 9067]='h00000000;
    rd_cycle[ 9068] = 1'b0;  wr_cycle[ 9068] = 1'b1;  addr_rom[ 9068]='h00000e8c;  wr_data_rom[ 9068]='h00001f44;
    rd_cycle[ 9069] = 1'b1;  wr_cycle[ 9069] = 1'b0;  addr_rom[ 9069]='h000018b4;  wr_data_rom[ 9069]='h00000000;
    rd_cycle[ 9070] = 1'b1;  wr_cycle[ 9070] = 1'b0;  addr_rom[ 9070]='h00000efc;  wr_data_rom[ 9070]='h00000000;
    rd_cycle[ 9071] = 1'b1;  wr_cycle[ 9071] = 1'b0;  addr_rom[ 9071]='h00003750;  wr_data_rom[ 9071]='h00000000;
    rd_cycle[ 9072] = 1'b1;  wr_cycle[ 9072] = 1'b0;  addr_rom[ 9072]='h00002b1c;  wr_data_rom[ 9072]='h00000000;
    rd_cycle[ 9073] = 1'b0;  wr_cycle[ 9073] = 1'b1;  addr_rom[ 9073]='h00001d80;  wr_data_rom[ 9073]='h000019bd;
    rd_cycle[ 9074] = 1'b0;  wr_cycle[ 9074] = 1'b1;  addr_rom[ 9074]='h00001ccc;  wr_data_rom[ 9074]='h00003930;
    rd_cycle[ 9075] = 1'b1;  wr_cycle[ 9075] = 1'b0;  addr_rom[ 9075]='h00003bd0;  wr_data_rom[ 9075]='h00000000;
    rd_cycle[ 9076] = 1'b1;  wr_cycle[ 9076] = 1'b0;  addr_rom[ 9076]='h00001b38;  wr_data_rom[ 9076]='h00000000;
    rd_cycle[ 9077] = 1'b0;  wr_cycle[ 9077] = 1'b1;  addr_rom[ 9077]='h00003b68;  wr_data_rom[ 9077]='h0000119c;
    rd_cycle[ 9078] = 1'b0;  wr_cycle[ 9078] = 1'b1;  addr_rom[ 9078]='h00001cd8;  wr_data_rom[ 9078]='h00003b26;
    rd_cycle[ 9079] = 1'b0;  wr_cycle[ 9079] = 1'b1;  addr_rom[ 9079]='h000023f8;  wr_data_rom[ 9079]='h00000d4a;
    rd_cycle[ 9080] = 1'b0;  wr_cycle[ 9080] = 1'b1;  addr_rom[ 9080]='h00002808;  wr_data_rom[ 9080]='h0000053d;
    rd_cycle[ 9081] = 1'b1;  wr_cycle[ 9081] = 1'b0;  addr_rom[ 9081]='h00000c4c;  wr_data_rom[ 9081]='h00000000;
    rd_cycle[ 9082] = 1'b1;  wr_cycle[ 9082] = 1'b0;  addr_rom[ 9082]='h00000248;  wr_data_rom[ 9082]='h00000000;
    rd_cycle[ 9083] = 1'b0;  wr_cycle[ 9083] = 1'b1;  addr_rom[ 9083]='h000029e0;  wr_data_rom[ 9083]='h00002312;
    rd_cycle[ 9084] = 1'b1;  wr_cycle[ 9084] = 1'b0;  addr_rom[ 9084]='h000035c0;  wr_data_rom[ 9084]='h00000000;
    rd_cycle[ 9085] = 1'b0;  wr_cycle[ 9085] = 1'b1;  addr_rom[ 9085]='h000015ac;  wr_data_rom[ 9085]='h00003189;
    rd_cycle[ 9086] = 1'b0;  wr_cycle[ 9086] = 1'b1;  addr_rom[ 9086]='h00000758;  wr_data_rom[ 9086]='h00000a7f;
    rd_cycle[ 9087] = 1'b1;  wr_cycle[ 9087] = 1'b0;  addr_rom[ 9087]='h000021d4;  wr_data_rom[ 9087]='h00000000;
    rd_cycle[ 9088] = 1'b0;  wr_cycle[ 9088] = 1'b1;  addr_rom[ 9088]='h00002de0;  wr_data_rom[ 9088]='h00002aa0;
    rd_cycle[ 9089] = 1'b1;  wr_cycle[ 9089] = 1'b0;  addr_rom[ 9089]='h00001b04;  wr_data_rom[ 9089]='h00000000;
    rd_cycle[ 9090] = 1'b0;  wr_cycle[ 9090] = 1'b1;  addr_rom[ 9090]='h0000213c;  wr_data_rom[ 9090]='h00001399;
    rd_cycle[ 9091] = 1'b0;  wr_cycle[ 9091] = 1'b1;  addr_rom[ 9091]='h00003c48;  wr_data_rom[ 9091]='h00000f1d;
    rd_cycle[ 9092] = 1'b0;  wr_cycle[ 9092] = 1'b1;  addr_rom[ 9092]='h00002a78;  wr_data_rom[ 9092]='h000030e5;
    rd_cycle[ 9093] = 1'b1;  wr_cycle[ 9093] = 1'b0;  addr_rom[ 9093]='h00001d7c;  wr_data_rom[ 9093]='h00000000;
    rd_cycle[ 9094] = 1'b0;  wr_cycle[ 9094] = 1'b1;  addr_rom[ 9094]='h00001114;  wr_data_rom[ 9094]='h00000812;
    rd_cycle[ 9095] = 1'b1;  wr_cycle[ 9095] = 1'b0;  addr_rom[ 9095]='h00002c08;  wr_data_rom[ 9095]='h00000000;
    rd_cycle[ 9096] = 1'b0;  wr_cycle[ 9096] = 1'b1;  addr_rom[ 9096]='h00001758;  wr_data_rom[ 9096]='h0000217d;
    rd_cycle[ 9097] = 1'b0;  wr_cycle[ 9097] = 1'b1;  addr_rom[ 9097]='h00002048;  wr_data_rom[ 9097]='h000034cd;
    rd_cycle[ 9098] = 1'b0;  wr_cycle[ 9098] = 1'b1;  addr_rom[ 9098]='h00002fac;  wr_data_rom[ 9098]='h00003ca3;
    rd_cycle[ 9099] = 1'b0;  wr_cycle[ 9099] = 1'b1;  addr_rom[ 9099]='h00001b14;  wr_data_rom[ 9099]='h00002079;
    rd_cycle[ 9100] = 1'b1;  wr_cycle[ 9100] = 1'b0;  addr_rom[ 9100]='h000035bc;  wr_data_rom[ 9100]='h00000000;
    rd_cycle[ 9101] = 1'b0;  wr_cycle[ 9101] = 1'b1;  addr_rom[ 9101]='h00003784;  wr_data_rom[ 9101]='h00002dd8;
    rd_cycle[ 9102] = 1'b1;  wr_cycle[ 9102] = 1'b0;  addr_rom[ 9102]='h00000024;  wr_data_rom[ 9102]='h00000000;
    rd_cycle[ 9103] = 1'b0;  wr_cycle[ 9103] = 1'b1;  addr_rom[ 9103]='h00002ad8;  wr_data_rom[ 9103]='h000016bb;
    rd_cycle[ 9104] = 1'b0;  wr_cycle[ 9104] = 1'b1;  addr_rom[ 9104]='h00003328;  wr_data_rom[ 9104]='h000000f1;
    rd_cycle[ 9105] = 1'b0;  wr_cycle[ 9105] = 1'b1;  addr_rom[ 9105]='h00001f40;  wr_data_rom[ 9105]='h00001c71;
    rd_cycle[ 9106] = 1'b0;  wr_cycle[ 9106] = 1'b1;  addr_rom[ 9106]='h0000252c;  wr_data_rom[ 9106]='h0000052d;
    rd_cycle[ 9107] = 1'b0;  wr_cycle[ 9107] = 1'b1;  addr_rom[ 9107]='h00001158;  wr_data_rom[ 9107]='h00000490;
    rd_cycle[ 9108] = 1'b0;  wr_cycle[ 9108] = 1'b1;  addr_rom[ 9108]='h00000bec;  wr_data_rom[ 9108]='h000039f9;
    rd_cycle[ 9109] = 1'b0;  wr_cycle[ 9109] = 1'b1;  addr_rom[ 9109]='h00003eb0;  wr_data_rom[ 9109]='h00002b85;
    rd_cycle[ 9110] = 1'b0;  wr_cycle[ 9110] = 1'b1;  addr_rom[ 9110]='h000016c4;  wr_data_rom[ 9110]='h00001c1c;
    rd_cycle[ 9111] = 1'b0;  wr_cycle[ 9111] = 1'b1;  addr_rom[ 9111]='h0000332c;  wr_data_rom[ 9111]='h00000e58;
    rd_cycle[ 9112] = 1'b0;  wr_cycle[ 9112] = 1'b1;  addr_rom[ 9112]='h00002f0c;  wr_data_rom[ 9112]='h000000e3;
    rd_cycle[ 9113] = 1'b0;  wr_cycle[ 9113] = 1'b1;  addr_rom[ 9113]='h00002a30;  wr_data_rom[ 9113]='h00003e87;
    rd_cycle[ 9114] = 1'b0;  wr_cycle[ 9114] = 1'b1;  addr_rom[ 9114]='h00003088;  wr_data_rom[ 9114]='h00002ab6;
    rd_cycle[ 9115] = 1'b1;  wr_cycle[ 9115] = 1'b0;  addr_rom[ 9115]='h00000c10;  wr_data_rom[ 9115]='h00000000;
    rd_cycle[ 9116] = 1'b1;  wr_cycle[ 9116] = 1'b0;  addr_rom[ 9116]='h00003cf0;  wr_data_rom[ 9116]='h00000000;
    rd_cycle[ 9117] = 1'b0;  wr_cycle[ 9117] = 1'b1;  addr_rom[ 9117]='h000023cc;  wr_data_rom[ 9117]='h0000119d;
    rd_cycle[ 9118] = 1'b0;  wr_cycle[ 9118] = 1'b1;  addr_rom[ 9118]='h00000584;  wr_data_rom[ 9118]='h00000716;
    rd_cycle[ 9119] = 1'b0;  wr_cycle[ 9119] = 1'b1;  addr_rom[ 9119]='h000000c0;  wr_data_rom[ 9119]='h00000ae1;
    rd_cycle[ 9120] = 1'b0;  wr_cycle[ 9120] = 1'b1;  addr_rom[ 9120]='h00003624;  wr_data_rom[ 9120]='h0000120f;
    rd_cycle[ 9121] = 1'b1;  wr_cycle[ 9121] = 1'b0;  addr_rom[ 9121]='h000017a0;  wr_data_rom[ 9121]='h00000000;
    rd_cycle[ 9122] = 1'b0;  wr_cycle[ 9122] = 1'b1;  addr_rom[ 9122]='h000000a8;  wr_data_rom[ 9122]='h00000b49;
    rd_cycle[ 9123] = 1'b0;  wr_cycle[ 9123] = 1'b1;  addr_rom[ 9123]='h000008fc;  wr_data_rom[ 9123]='h000036ec;
    rd_cycle[ 9124] = 1'b0;  wr_cycle[ 9124] = 1'b1;  addr_rom[ 9124]='h00003cd4;  wr_data_rom[ 9124]='h00003f3b;
    rd_cycle[ 9125] = 1'b1;  wr_cycle[ 9125] = 1'b0;  addr_rom[ 9125]='h00003dc4;  wr_data_rom[ 9125]='h00000000;
    rd_cycle[ 9126] = 1'b0;  wr_cycle[ 9126] = 1'b1;  addr_rom[ 9126]='h00001a88;  wr_data_rom[ 9126]='h00001bf7;
    rd_cycle[ 9127] = 1'b0;  wr_cycle[ 9127] = 1'b1;  addr_rom[ 9127]='h00001718;  wr_data_rom[ 9127]='h00001311;
    rd_cycle[ 9128] = 1'b1;  wr_cycle[ 9128] = 1'b0;  addr_rom[ 9128]='h00001c3c;  wr_data_rom[ 9128]='h00000000;
    rd_cycle[ 9129] = 1'b0;  wr_cycle[ 9129] = 1'b1;  addr_rom[ 9129]='h00000250;  wr_data_rom[ 9129]='h000012f9;
    rd_cycle[ 9130] = 1'b0;  wr_cycle[ 9130] = 1'b1;  addr_rom[ 9130]='h00003c40;  wr_data_rom[ 9130]='h00003d7d;
    rd_cycle[ 9131] = 1'b0;  wr_cycle[ 9131] = 1'b1;  addr_rom[ 9131]='h00002dd4;  wr_data_rom[ 9131]='h0000329c;
    rd_cycle[ 9132] = 1'b1;  wr_cycle[ 9132] = 1'b0;  addr_rom[ 9132]='h00002074;  wr_data_rom[ 9132]='h00000000;
    rd_cycle[ 9133] = 1'b1;  wr_cycle[ 9133] = 1'b0;  addr_rom[ 9133]='h000013dc;  wr_data_rom[ 9133]='h00000000;
    rd_cycle[ 9134] = 1'b1;  wr_cycle[ 9134] = 1'b0;  addr_rom[ 9134]='h00003038;  wr_data_rom[ 9134]='h00000000;
    rd_cycle[ 9135] = 1'b1;  wr_cycle[ 9135] = 1'b0;  addr_rom[ 9135]='h00003fb8;  wr_data_rom[ 9135]='h00000000;
    rd_cycle[ 9136] = 1'b0;  wr_cycle[ 9136] = 1'b1;  addr_rom[ 9136]='h00002020;  wr_data_rom[ 9136]='h00000ec6;
    rd_cycle[ 9137] = 1'b1;  wr_cycle[ 9137] = 1'b0;  addr_rom[ 9137]='h00003324;  wr_data_rom[ 9137]='h00000000;
    rd_cycle[ 9138] = 1'b0;  wr_cycle[ 9138] = 1'b1;  addr_rom[ 9138]='h000037b8;  wr_data_rom[ 9138]='h000005a6;
    rd_cycle[ 9139] = 1'b0;  wr_cycle[ 9139] = 1'b1;  addr_rom[ 9139]='h000025ec;  wr_data_rom[ 9139]='h00002cd4;
    rd_cycle[ 9140] = 1'b1;  wr_cycle[ 9140] = 1'b0;  addr_rom[ 9140]='h00000844;  wr_data_rom[ 9140]='h00000000;
    rd_cycle[ 9141] = 1'b0;  wr_cycle[ 9141] = 1'b1;  addr_rom[ 9141]='h00003f10;  wr_data_rom[ 9141]='h00001452;
    rd_cycle[ 9142] = 1'b0;  wr_cycle[ 9142] = 1'b1;  addr_rom[ 9142]='h0000353c;  wr_data_rom[ 9142]='h00003a1b;
    rd_cycle[ 9143] = 1'b1;  wr_cycle[ 9143] = 1'b0;  addr_rom[ 9143]='h00000ef8;  wr_data_rom[ 9143]='h00000000;
    rd_cycle[ 9144] = 1'b0;  wr_cycle[ 9144] = 1'b1;  addr_rom[ 9144]='h00001f08;  wr_data_rom[ 9144]='h000014cf;
    rd_cycle[ 9145] = 1'b0;  wr_cycle[ 9145] = 1'b1;  addr_rom[ 9145]='h00000be0;  wr_data_rom[ 9145]='h00003d23;
    rd_cycle[ 9146] = 1'b1;  wr_cycle[ 9146] = 1'b0;  addr_rom[ 9146]='h000030b8;  wr_data_rom[ 9146]='h00000000;
    rd_cycle[ 9147] = 1'b1;  wr_cycle[ 9147] = 1'b0;  addr_rom[ 9147]='h00003474;  wr_data_rom[ 9147]='h00000000;
    rd_cycle[ 9148] = 1'b1;  wr_cycle[ 9148] = 1'b0;  addr_rom[ 9148]='h00002424;  wr_data_rom[ 9148]='h00000000;
    rd_cycle[ 9149] = 1'b1;  wr_cycle[ 9149] = 1'b0;  addr_rom[ 9149]='h00001a9c;  wr_data_rom[ 9149]='h00000000;
    rd_cycle[ 9150] = 1'b1;  wr_cycle[ 9150] = 1'b0;  addr_rom[ 9150]='h000016e4;  wr_data_rom[ 9150]='h00000000;
    rd_cycle[ 9151] = 1'b0;  wr_cycle[ 9151] = 1'b1;  addr_rom[ 9151]='h00001e04;  wr_data_rom[ 9151]='h00000ee0;
    rd_cycle[ 9152] = 1'b1;  wr_cycle[ 9152] = 1'b0;  addr_rom[ 9152]='h0000280c;  wr_data_rom[ 9152]='h00000000;
    rd_cycle[ 9153] = 1'b0;  wr_cycle[ 9153] = 1'b1;  addr_rom[ 9153]='h00000a68;  wr_data_rom[ 9153]='h00003d35;
    rd_cycle[ 9154] = 1'b0;  wr_cycle[ 9154] = 1'b1;  addr_rom[ 9154]='h00001064;  wr_data_rom[ 9154]='h00002a32;
    rd_cycle[ 9155] = 1'b1;  wr_cycle[ 9155] = 1'b0;  addr_rom[ 9155]='h00003a14;  wr_data_rom[ 9155]='h00000000;
    rd_cycle[ 9156] = 1'b1;  wr_cycle[ 9156] = 1'b0;  addr_rom[ 9156]='h000020e0;  wr_data_rom[ 9156]='h00000000;
    rd_cycle[ 9157] = 1'b0;  wr_cycle[ 9157] = 1'b1;  addr_rom[ 9157]='h00000000;  wr_data_rom[ 9157]='h00003530;
    rd_cycle[ 9158] = 1'b1;  wr_cycle[ 9158] = 1'b0;  addr_rom[ 9158]='h00002810;  wr_data_rom[ 9158]='h00000000;
    rd_cycle[ 9159] = 1'b1;  wr_cycle[ 9159] = 1'b0;  addr_rom[ 9159]='h000014a4;  wr_data_rom[ 9159]='h00000000;
    rd_cycle[ 9160] = 1'b1;  wr_cycle[ 9160] = 1'b0;  addr_rom[ 9160]='h000026d0;  wr_data_rom[ 9160]='h00000000;
    rd_cycle[ 9161] = 1'b1;  wr_cycle[ 9161] = 1'b0;  addr_rom[ 9161]='h00002008;  wr_data_rom[ 9161]='h00000000;
    rd_cycle[ 9162] = 1'b1;  wr_cycle[ 9162] = 1'b0;  addr_rom[ 9162]='h00003470;  wr_data_rom[ 9162]='h00000000;
    rd_cycle[ 9163] = 1'b0;  wr_cycle[ 9163] = 1'b1;  addr_rom[ 9163]='h0000322c;  wr_data_rom[ 9163]='h00001046;
    rd_cycle[ 9164] = 1'b1;  wr_cycle[ 9164] = 1'b0;  addr_rom[ 9164]='h00002008;  wr_data_rom[ 9164]='h00000000;
    rd_cycle[ 9165] = 1'b0;  wr_cycle[ 9165] = 1'b1;  addr_rom[ 9165]='h00002b14;  wr_data_rom[ 9165]='h00003ce1;
    rd_cycle[ 9166] = 1'b1;  wr_cycle[ 9166] = 1'b0;  addr_rom[ 9166]='h000017ec;  wr_data_rom[ 9166]='h00000000;
    rd_cycle[ 9167] = 1'b1;  wr_cycle[ 9167] = 1'b0;  addr_rom[ 9167]='h000011f4;  wr_data_rom[ 9167]='h00000000;
    rd_cycle[ 9168] = 1'b0;  wr_cycle[ 9168] = 1'b1;  addr_rom[ 9168]='h00001190;  wr_data_rom[ 9168]='h00002986;
    rd_cycle[ 9169] = 1'b1;  wr_cycle[ 9169] = 1'b0;  addr_rom[ 9169]='h000034a4;  wr_data_rom[ 9169]='h00000000;
    rd_cycle[ 9170] = 1'b1;  wr_cycle[ 9170] = 1'b0;  addr_rom[ 9170]='h0000207c;  wr_data_rom[ 9170]='h00000000;
    rd_cycle[ 9171] = 1'b0;  wr_cycle[ 9171] = 1'b1;  addr_rom[ 9171]='h00002500;  wr_data_rom[ 9171]='h00001a91;
    rd_cycle[ 9172] = 1'b1;  wr_cycle[ 9172] = 1'b0;  addr_rom[ 9172]='h00001650;  wr_data_rom[ 9172]='h00000000;
    rd_cycle[ 9173] = 1'b0;  wr_cycle[ 9173] = 1'b1;  addr_rom[ 9173]='h00003420;  wr_data_rom[ 9173]='h000017ce;
    rd_cycle[ 9174] = 1'b0;  wr_cycle[ 9174] = 1'b1;  addr_rom[ 9174]='h00000fd4;  wr_data_rom[ 9174]='h0000140c;
    rd_cycle[ 9175] = 1'b0;  wr_cycle[ 9175] = 1'b1;  addr_rom[ 9175]='h00003cfc;  wr_data_rom[ 9175]='h000039a2;
    rd_cycle[ 9176] = 1'b1;  wr_cycle[ 9176] = 1'b0;  addr_rom[ 9176]='h00002ea0;  wr_data_rom[ 9176]='h00000000;
    rd_cycle[ 9177] = 1'b0;  wr_cycle[ 9177] = 1'b1;  addr_rom[ 9177]='h00002a34;  wr_data_rom[ 9177]='h0000286f;
    rd_cycle[ 9178] = 1'b0;  wr_cycle[ 9178] = 1'b1;  addr_rom[ 9178]='h00001c48;  wr_data_rom[ 9178]='h00000a4a;
    rd_cycle[ 9179] = 1'b0;  wr_cycle[ 9179] = 1'b1;  addr_rom[ 9179]='h00001b50;  wr_data_rom[ 9179]='h000006e0;
    rd_cycle[ 9180] = 1'b1;  wr_cycle[ 9180] = 1'b0;  addr_rom[ 9180]='h0000374c;  wr_data_rom[ 9180]='h00000000;
    rd_cycle[ 9181] = 1'b0;  wr_cycle[ 9181] = 1'b1;  addr_rom[ 9181]='h000000ec;  wr_data_rom[ 9181]='h00000b35;
    rd_cycle[ 9182] = 1'b0;  wr_cycle[ 9182] = 1'b1;  addr_rom[ 9182]='h00001d94;  wr_data_rom[ 9182]='h00000507;
    rd_cycle[ 9183] = 1'b0;  wr_cycle[ 9183] = 1'b1;  addr_rom[ 9183]='h0000026c;  wr_data_rom[ 9183]='h00000996;
    rd_cycle[ 9184] = 1'b0;  wr_cycle[ 9184] = 1'b1;  addr_rom[ 9184]='h000030dc;  wr_data_rom[ 9184]='h00000563;
    rd_cycle[ 9185] = 1'b1;  wr_cycle[ 9185] = 1'b0;  addr_rom[ 9185]='h000039c8;  wr_data_rom[ 9185]='h00000000;
    rd_cycle[ 9186] = 1'b1;  wr_cycle[ 9186] = 1'b0;  addr_rom[ 9186]='h00003a90;  wr_data_rom[ 9186]='h00000000;
    rd_cycle[ 9187] = 1'b0;  wr_cycle[ 9187] = 1'b1;  addr_rom[ 9187]='h00003d08;  wr_data_rom[ 9187]='h00000420;
    rd_cycle[ 9188] = 1'b0;  wr_cycle[ 9188] = 1'b1;  addr_rom[ 9188]='h00001838;  wr_data_rom[ 9188]='h0000057c;
    rd_cycle[ 9189] = 1'b1;  wr_cycle[ 9189] = 1'b0;  addr_rom[ 9189]='h00000af8;  wr_data_rom[ 9189]='h00000000;
    rd_cycle[ 9190] = 1'b0;  wr_cycle[ 9190] = 1'b1;  addr_rom[ 9190]='h000024b4;  wr_data_rom[ 9190]='h00002bc8;
    rd_cycle[ 9191] = 1'b0;  wr_cycle[ 9191] = 1'b1;  addr_rom[ 9191]='h00001634;  wr_data_rom[ 9191]='h00001f30;
    rd_cycle[ 9192] = 1'b0;  wr_cycle[ 9192] = 1'b1;  addr_rom[ 9192]='h0000210c;  wr_data_rom[ 9192]='h000034ff;
    rd_cycle[ 9193] = 1'b1;  wr_cycle[ 9193] = 1'b0;  addr_rom[ 9193]='h00003b6c;  wr_data_rom[ 9193]='h00000000;
    rd_cycle[ 9194] = 1'b0;  wr_cycle[ 9194] = 1'b1;  addr_rom[ 9194]='h00001d00;  wr_data_rom[ 9194]='h00001f43;
    rd_cycle[ 9195] = 1'b1;  wr_cycle[ 9195] = 1'b0;  addr_rom[ 9195]='h000004b4;  wr_data_rom[ 9195]='h00000000;
    rd_cycle[ 9196] = 1'b0;  wr_cycle[ 9196] = 1'b1;  addr_rom[ 9196]='h00002404;  wr_data_rom[ 9196]='h00002840;
    rd_cycle[ 9197] = 1'b0;  wr_cycle[ 9197] = 1'b1;  addr_rom[ 9197]='h00001d2c;  wr_data_rom[ 9197]='h00000ff4;
    rd_cycle[ 9198] = 1'b0;  wr_cycle[ 9198] = 1'b1;  addr_rom[ 9198]='h000028b4;  wr_data_rom[ 9198]='h0000378e;
    rd_cycle[ 9199] = 1'b0;  wr_cycle[ 9199] = 1'b1;  addr_rom[ 9199]='h0000026c;  wr_data_rom[ 9199]='h00001e45;
    rd_cycle[ 9200] = 1'b1;  wr_cycle[ 9200] = 1'b0;  addr_rom[ 9200]='h000008e4;  wr_data_rom[ 9200]='h00000000;
    rd_cycle[ 9201] = 1'b0;  wr_cycle[ 9201] = 1'b1;  addr_rom[ 9201]='h00000df4;  wr_data_rom[ 9201]='h0000195f;
    rd_cycle[ 9202] = 1'b1;  wr_cycle[ 9202] = 1'b0;  addr_rom[ 9202]='h000012d0;  wr_data_rom[ 9202]='h00000000;
    rd_cycle[ 9203] = 1'b0;  wr_cycle[ 9203] = 1'b1;  addr_rom[ 9203]='h00000e3c;  wr_data_rom[ 9203]='h00003cca;
    rd_cycle[ 9204] = 1'b1;  wr_cycle[ 9204] = 1'b0;  addr_rom[ 9204]='h000011f8;  wr_data_rom[ 9204]='h00000000;
    rd_cycle[ 9205] = 1'b1;  wr_cycle[ 9205] = 1'b0;  addr_rom[ 9205]='h00001204;  wr_data_rom[ 9205]='h00000000;
    rd_cycle[ 9206] = 1'b0;  wr_cycle[ 9206] = 1'b1;  addr_rom[ 9206]='h00001bbc;  wr_data_rom[ 9206]='h000025b4;
    rd_cycle[ 9207] = 1'b1;  wr_cycle[ 9207] = 1'b0;  addr_rom[ 9207]='h00000d6c;  wr_data_rom[ 9207]='h00000000;
    rd_cycle[ 9208] = 1'b1;  wr_cycle[ 9208] = 1'b0;  addr_rom[ 9208]='h00000dc8;  wr_data_rom[ 9208]='h00000000;
    rd_cycle[ 9209] = 1'b1;  wr_cycle[ 9209] = 1'b0;  addr_rom[ 9209]='h00001350;  wr_data_rom[ 9209]='h00000000;
    rd_cycle[ 9210] = 1'b1;  wr_cycle[ 9210] = 1'b0;  addr_rom[ 9210]='h000026f4;  wr_data_rom[ 9210]='h00000000;
    rd_cycle[ 9211] = 1'b1;  wr_cycle[ 9211] = 1'b0;  addr_rom[ 9211]='h000025b0;  wr_data_rom[ 9211]='h00000000;
    rd_cycle[ 9212] = 1'b0;  wr_cycle[ 9212] = 1'b1;  addr_rom[ 9212]='h00000930;  wr_data_rom[ 9212]='h00002d12;
    rd_cycle[ 9213] = 1'b0;  wr_cycle[ 9213] = 1'b1;  addr_rom[ 9213]='h00002bfc;  wr_data_rom[ 9213]='h00001d65;
    rd_cycle[ 9214] = 1'b1;  wr_cycle[ 9214] = 1'b0;  addr_rom[ 9214]='h000035d4;  wr_data_rom[ 9214]='h00000000;
    rd_cycle[ 9215] = 1'b0;  wr_cycle[ 9215] = 1'b1;  addr_rom[ 9215]='h00000288;  wr_data_rom[ 9215]='h00002e62;
    rd_cycle[ 9216] = 1'b0;  wr_cycle[ 9216] = 1'b1;  addr_rom[ 9216]='h000010b4;  wr_data_rom[ 9216]='h000034da;
    rd_cycle[ 9217] = 1'b0;  wr_cycle[ 9217] = 1'b1;  addr_rom[ 9217]='h0000154c;  wr_data_rom[ 9217]='h00002a97;
    rd_cycle[ 9218] = 1'b0;  wr_cycle[ 9218] = 1'b1;  addr_rom[ 9218]='h00000a24;  wr_data_rom[ 9218]='h00001cee;
    rd_cycle[ 9219] = 1'b0;  wr_cycle[ 9219] = 1'b1;  addr_rom[ 9219]='h00003cd8;  wr_data_rom[ 9219]='h000002dd;
    rd_cycle[ 9220] = 1'b1;  wr_cycle[ 9220] = 1'b0;  addr_rom[ 9220]='h00000b44;  wr_data_rom[ 9220]='h00000000;
    rd_cycle[ 9221] = 1'b1;  wr_cycle[ 9221] = 1'b0;  addr_rom[ 9221]='h0000038c;  wr_data_rom[ 9221]='h00000000;
    rd_cycle[ 9222] = 1'b1;  wr_cycle[ 9222] = 1'b0;  addr_rom[ 9222]='h0000040c;  wr_data_rom[ 9222]='h00000000;
    rd_cycle[ 9223] = 1'b0;  wr_cycle[ 9223] = 1'b1;  addr_rom[ 9223]='h00002a84;  wr_data_rom[ 9223]='h00003791;
    rd_cycle[ 9224] = 1'b1;  wr_cycle[ 9224] = 1'b0;  addr_rom[ 9224]='h00001848;  wr_data_rom[ 9224]='h00000000;
    rd_cycle[ 9225] = 1'b1;  wr_cycle[ 9225] = 1'b0;  addr_rom[ 9225]='h000002dc;  wr_data_rom[ 9225]='h00000000;
    rd_cycle[ 9226] = 1'b0;  wr_cycle[ 9226] = 1'b1;  addr_rom[ 9226]='h00003d08;  wr_data_rom[ 9226]='h00003bd4;
    rd_cycle[ 9227] = 1'b1;  wr_cycle[ 9227] = 1'b0;  addr_rom[ 9227]='h000034b4;  wr_data_rom[ 9227]='h00000000;
    rd_cycle[ 9228] = 1'b1;  wr_cycle[ 9228] = 1'b0;  addr_rom[ 9228]='h0000245c;  wr_data_rom[ 9228]='h00000000;
    rd_cycle[ 9229] = 1'b0;  wr_cycle[ 9229] = 1'b1;  addr_rom[ 9229]='h00002264;  wr_data_rom[ 9229]='h00001647;
    rd_cycle[ 9230] = 1'b1;  wr_cycle[ 9230] = 1'b0;  addr_rom[ 9230]='h00000fa4;  wr_data_rom[ 9230]='h00000000;
    rd_cycle[ 9231] = 1'b1;  wr_cycle[ 9231] = 1'b0;  addr_rom[ 9231]='h0000117c;  wr_data_rom[ 9231]='h00000000;
    rd_cycle[ 9232] = 1'b1;  wr_cycle[ 9232] = 1'b0;  addr_rom[ 9232]='h00000648;  wr_data_rom[ 9232]='h00000000;
    rd_cycle[ 9233] = 1'b1;  wr_cycle[ 9233] = 1'b0;  addr_rom[ 9233]='h00001f5c;  wr_data_rom[ 9233]='h00000000;
    rd_cycle[ 9234] = 1'b0;  wr_cycle[ 9234] = 1'b1;  addr_rom[ 9234]='h000030cc;  wr_data_rom[ 9234]='h0000060d;
    rd_cycle[ 9235] = 1'b0;  wr_cycle[ 9235] = 1'b1;  addr_rom[ 9235]='h000025d8;  wr_data_rom[ 9235]='h000006da;
    rd_cycle[ 9236] = 1'b1;  wr_cycle[ 9236] = 1'b0;  addr_rom[ 9236]='h000039bc;  wr_data_rom[ 9236]='h00000000;
    rd_cycle[ 9237] = 1'b0;  wr_cycle[ 9237] = 1'b1;  addr_rom[ 9237]='h0000338c;  wr_data_rom[ 9237]='h000023b5;
    rd_cycle[ 9238] = 1'b1;  wr_cycle[ 9238] = 1'b0;  addr_rom[ 9238]='h00001094;  wr_data_rom[ 9238]='h00000000;
    rd_cycle[ 9239] = 1'b0;  wr_cycle[ 9239] = 1'b1;  addr_rom[ 9239]='h000018c4;  wr_data_rom[ 9239]='h000005e7;
    rd_cycle[ 9240] = 1'b1;  wr_cycle[ 9240] = 1'b0;  addr_rom[ 9240]='h00002450;  wr_data_rom[ 9240]='h00000000;
    rd_cycle[ 9241] = 1'b0;  wr_cycle[ 9241] = 1'b1;  addr_rom[ 9241]='h00000518;  wr_data_rom[ 9241]='h000021ae;
    rd_cycle[ 9242] = 1'b0;  wr_cycle[ 9242] = 1'b1;  addr_rom[ 9242]='h000031f8;  wr_data_rom[ 9242]='h0000279f;
    rd_cycle[ 9243] = 1'b0;  wr_cycle[ 9243] = 1'b1;  addr_rom[ 9243]='h00001d74;  wr_data_rom[ 9243]='h00002a9f;
    rd_cycle[ 9244] = 1'b1;  wr_cycle[ 9244] = 1'b0;  addr_rom[ 9244]='h00002ed8;  wr_data_rom[ 9244]='h00000000;
    rd_cycle[ 9245] = 1'b0;  wr_cycle[ 9245] = 1'b1;  addr_rom[ 9245]='h00001788;  wr_data_rom[ 9245]='h000015a9;
    rd_cycle[ 9246] = 1'b1;  wr_cycle[ 9246] = 1'b0;  addr_rom[ 9246]='h000009c0;  wr_data_rom[ 9246]='h00000000;
    rd_cycle[ 9247] = 1'b0;  wr_cycle[ 9247] = 1'b1;  addr_rom[ 9247]='h00002c80;  wr_data_rom[ 9247]='h00001b8b;
    rd_cycle[ 9248] = 1'b0;  wr_cycle[ 9248] = 1'b1;  addr_rom[ 9248]='h000010f8;  wr_data_rom[ 9248]='h00002e3e;
    rd_cycle[ 9249] = 1'b1;  wr_cycle[ 9249] = 1'b0;  addr_rom[ 9249]='h00000744;  wr_data_rom[ 9249]='h00000000;
    rd_cycle[ 9250] = 1'b0;  wr_cycle[ 9250] = 1'b1;  addr_rom[ 9250]='h00003e2c;  wr_data_rom[ 9250]='h00000fb9;
    rd_cycle[ 9251] = 1'b1;  wr_cycle[ 9251] = 1'b0;  addr_rom[ 9251]='h00002c98;  wr_data_rom[ 9251]='h00000000;
    rd_cycle[ 9252] = 1'b0;  wr_cycle[ 9252] = 1'b1;  addr_rom[ 9252]='h00001d8c;  wr_data_rom[ 9252]='h00000272;
    rd_cycle[ 9253] = 1'b0;  wr_cycle[ 9253] = 1'b1;  addr_rom[ 9253]='h00001438;  wr_data_rom[ 9253]='h000010dc;
    rd_cycle[ 9254] = 1'b1;  wr_cycle[ 9254] = 1'b0;  addr_rom[ 9254]='h00001818;  wr_data_rom[ 9254]='h00000000;
    rd_cycle[ 9255] = 1'b1;  wr_cycle[ 9255] = 1'b0;  addr_rom[ 9255]='h000023d4;  wr_data_rom[ 9255]='h00000000;
    rd_cycle[ 9256] = 1'b1;  wr_cycle[ 9256] = 1'b0;  addr_rom[ 9256]='h000016a4;  wr_data_rom[ 9256]='h00000000;
    rd_cycle[ 9257] = 1'b0;  wr_cycle[ 9257] = 1'b1;  addr_rom[ 9257]='h00001370;  wr_data_rom[ 9257]='h00003f02;
    rd_cycle[ 9258] = 1'b0;  wr_cycle[ 9258] = 1'b1;  addr_rom[ 9258]='h00002800;  wr_data_rom[ 9258]='h000028e0;
    rd_cycle[ 9259] = 1'b1;  wr_cycle[ 9259] = 1'b0;  addr_rom[ 9259]='h00002ee8;  wr_data_rom[ 9259]='h00000000;
    rd_cycle[ 9260] = 1'b1;  wr_cycle[ 9260] = 1'b0;  addr_rom[ 9260]='h000018ec;  wr_data_rom[ 9260]='h00000000;
    rd_cycle[ 9261] = 1'b1;  wr_cycle[ 9261] = 1'b0;  addr_rom[ 9261]='h000039a4;  wr_data_rom[ 9261]='h00000000;
    rd_cycle[ 9262] = 1'b1;  wr_cycle[ 9262] = 1'b0;  addr_rom[ 9262]='h00003da0;  wr_data_rom[ 9262]='h00000000;
    rd_cycle[ 9263] = 1'b1;  wr_cycle[ 9263] = 1'b0;  addr_rom[ 9263]='h00000738;  wr_data_rom[ 9263]='h00000000;
    rd_cycle[ 9264] = 1'b0;  wr_cycle[ 9264] = 1'b1;  addr_rom[ 9264]='h00003718;  wr_data_rom[ 9264]='h00003f85;
    rd_cycle[ 9265] = 1'b0;  wr_cycle[ 9265] = 1'b1;  addr_rom[ 9265]='h000010f4;  wr_data_rom[ 9265]='h00000fa8;
    rd_cycle[ 9266] = 1'b1;  wr_cycle[ 9266] = 1'b0;  addr_rom[ 9266]='h000026f0;  wr_data_rom[ 9266]='h00000000;
    rd_cycle[ 9267] = 1'b1;  wr_cycle[ 9267] = 1'b0;  addr_rom[ 9267]='h000000c8;  wr_data_rom[ 9267]='h00000000;
    rd_cycle[ 9268] = 1'b1;  wr_cycle[ 9268] = 1'b0;  addr_rom[ 9268]='h00000c70;  wr_data_rom[ 9268]='h00000000;
    rd_cycle[ 9269] = 1'b1;  wr_cycle[ 9269] = 1'b0;  addr_rom[ 9269]='h00001204;  wr_data_rom[ 9269]='h00000000;
    rd_cycle[ 9270] = 1'b0;  wr_cycle[ 9270] = 1'b1;  addr_rom[ 9270]='h00002ad8;  wr_data_rom[ 9270]='h00002d51;
    rd_cycle[ 9271] = 1'b0;  wr_cycle[ 9271] = 1'b1;  addr_rom[ 9271]='h00002978;  wr_data_rom[ 9271]='h00002d02;
    rd_cycle[ 9272] = 1'b1;  wr_cycle[ 9272] = 1'b0;  addr_rom[ 9272]='h00002e7c;  wr_data_rom[ 9272]='h00000000;
    rd_cycle[ 9273] = 1'b1;  wr_cycle[ 9273] = 1'b0;  addr_rom[ 9273]='h00001048;  wr_data_rom[ 9273]='h00000000;
    rd_cycle[ 9274] = 1'b1;  wr_cycle[ 9274] = 1'b0;  addr_rom[ 9274]='h000011c0;  wr_data_rom[ 9274]='h00000000;
    rd_cycle[ 9275] = 1'b0;  wr_cycle[ 9275] = 1'b1;  addr_rom[ 9275]='h00002e9c;  wr_data_rom[ 9275]='h00003d30;
    rd_cycle[ 9276] = 1'b1;  wr_cycle[ 9276] = 1'b0;  addr_rom[ 9276]='h00000d44;  wr_data_rom[ 9276]='h00000000;
    rd_cycle[ 9277] = 1'b0;  wr_cycle[ 9277] = 1'b1;  addr_rom[ 9277]='h00000c44;  wr_data_rom[ 9277]='h00000039;
    rd_cycle[ 9278] = 1'b0;  wr_cycle[ 9278] = 1'b1;  addr_rom[ 9278]='h00002dbc;  wr_data_rom[ 9278]='h000005a0;
    rd_cycle[ 9279] = 1'b1;  wr_cycle[ 9279] = 1'b0;  addr_rom[ 9279]='h00003654;  wr_data_rom[ 9279]='h00000000;
    rd_cycle[ 9280] = 1'b1;  wr_cycle[ 9280] = 1'b0;  addr_rom[ 9280]='h00003204;  wr_data_rom[ 9280]='h00000000;
    rd_cycle[ 9281] = 1'b0;  wr_cycle[ 9281] = 1'b1;  addr_rom[ 9281]='h00002768;  wr_data_rom[ 9281]='h00002ce0;
    rd_cycle[ 9282] = 1'b1;  wr_cycle[ 9282] = 1'b0;  addr_rom[ 9282]='h00000808;  wr_data_rom[ 9282]='h00000000;
    rd_cycle[ 9283] = 1'b1;  wr_cycle[ 9283] = 1'b0;  addr_rom[ 9283]='h00001fc0;  wr_data_rom[ 9283]='h00000000;
    rd_cycle[ 9284] = 1'b0;  wr_cycle[ 9284] = 1'b1;  addr_rom[ 9284]='h00001bc0;  wr_data_rom[ 9284]='h0000118b;
    rd_cycle[ 9285] = 1'b1;  wr_cycle[ 9285] = 1'b0;  addr_rom[ 9285]='h00002e74;  wr_data_rom[ 9285]='h00000000;
    rd_cycle[ 9286] = 1'b1;  wr_cycle[ 9286] = 1'b0;  addr_rom[ 9286]='h000002d0;  wr_data_rom[ 9286]='h00000000;
    rd_cycle[ 9287] = 1'b1;  wr_cycle[ 9287] = 1'b0;  addr_rom[ 9287]='h00002ae0;  wr_data_rom[ 9287]='h00000000;
    rd_cycle[ 9288] = 1'b1;  wr_cycle[ 9288] = 1'b0;  addr_rom[ 9288]='h000014c8;  wr_data_rom[ 9288]='h00000000;
    rd_cycle[ 9289] = 1'b0;  wr_cycle[ 9289] = 1'b1;  addr_rom[ 9289]='h0000354c;  wr_data_rom[ 9289]='h00000bd6;
    rd_cycle[ 9290] = 1'b1;  wr_cycle[ 9290] = 1'b0;  addr_rom[ 9290]='h000035dc;  wr_data_rom[ 9290]='h00000000;
    rd_cycle[ 9291] = 1'b1;  wr_cycle[ 9291] = 1'b0;  addr_rom[ 9291]='h00002cc0;  wr_data_rom[ 9291]='h00000000;
    rd_cycle[ 9292] = 1'b1;  wr_cycle[ 9292] = 1'b0;  addr_rom[ 9292]='h000007fc;  wr_data_rom[ 9292]='h00000000;
    rd_cycle[ 9293] = 1'b0;  wr_cycle[ 9293] = 1'b1;  addr_rom[ 9293]='h000012b0;  wr_data_rom[ 9293]='h00003b0c;
    rd_cycle[ 9294] = 1'b1;  wr_cycle[ 9294] = 1'b0;  addr_rom[ 9294]='h00001354;  wr_data_rom[ 9294]='h00000000;
    rd_cycle[ 9295] = 1'b1;  wr_cycle[ 9295] = 1'b0;  addr_rom[ 9295]='h000023d8;  wr_data_rom[ 9295]='h00000000;
    rd_cycle[ 9296] = 1'b0;  wr_cycle[ 9296] = 1'b1;  addr_rom[ 9296]='h00001c90;  wr_data_rom[ 9296]='h000000ed;
    rd_cycle[ 9297] = 1'b0;  wr_cycle[ 9297] = 1'b1;  addr_rom[ 9297]='h0000262c;  wr_data_rom[ 9297]='h00003b13;
    rd_cycle[ 9298] = 1'b0;  wr_cycle[ 9298] = 1'b1;  addr_rom[ 9298]='h00003a14;  wr_data_rom[ 9298]='h000025d1;
    rd_cycle[ 9299] = 1'b1;  wr_cycle[ 9299] = 1'b0;  addr_rom[ 9299]='h00001d04;  wr_data_rom[ 9299]='h00000000;
    rd_cycle[ 9300] = 1'b1;  wr_cycle[ 9300] = 1'b0;  addr_rom[ 9300]='h00003bb8;  wr_data_rom[ 9300]='h00000000;
    rd_cycle[ 9301] = 1'b1;  wr_cycle[ 9301] = 1'b0;  addr_rom[ 9301]='h0000353c;  wr_data_rom[ 9301]='h00000000;
    rd_cycle[ 9302] = 1'b0;  wr_cycle[ 9302] = 1'b1;  addr_rom[ 9302]='h000030f0;  wr_data_rom[ 9302]='h00003ff3;
    rd_cycle[ 9303] = 1'b0;  wr_cycle[ 9303] = 1'b1;  addr_rom[ 9303]='h00003b04;  wr_data_rom[ 9303]='h000029a9;
    rd_cycle[ 9304] = 1'b0;  wr_cycle[ 9304] = 1'b1;  addr_rom[ 9304]='h00001944;  wr_data_rom[ 9304]='h00003907;
    rd_cycle[ 9305] = 1'b0;  wr_cycle[ 9305] = 1'b1;  addr_rom[ 9305]='h0000222c;  wr_data_rom[ 9305]='h00000366;
    rd_cycle[ 9306] = 1'b0;  wr_cycle[ 9306] = 1'b1;  addr_rom[ 9306]='h0000037c;  wr_data_rom[ 9306]='h00000a04;
    rd_cycle[ 9307] = 1'b0;  wr_cycle[ 9307] = 1'b1;  addr_rom[ 9307]='h000012dc;  wr_data_rom[ 9307]='h00002da5;
    rd_cycle[ 9308] = 1'b0;  wr_cycle[ 9308] = 1'b1;  addr_rom[ 9308]='h00000500;  wr_data_rom[ 9308]='h00001ebc;
    rd_cycle[ 9309] = 1'b0;  wr_cycle[ 9309] = 1'b1;  addr_rom[ 9309]='h00001790;  wr_data_rom[ 9309]='h0000253c;
    rd_cycle[ 9310] = 1'b1;  wr_cycle[ 9310] = 1'b0;  addr_rom[ 9310]='h00003558;  wr_data_rom[ 9310]='h00000000;
    rd_cycle[ 9311] = 1'b1;  wr_cycle[ 9311] = 1'b0;  addr_rom[ 9311]='h000002bc;  wr_data_rom[ 9311]='h00000000;
    rd_cycle[ 9312] = 1'b0;  wr_cycle[ 9312] = 1'b1;  addr_rom[ 9312]='h00002074;  wr_data_rom[ 9312]='h0000100e;
    rd_cycle[ 9313] = 1'b0;  wr_cycle[ 9313] = 1'b1;  addr_rom[ 9313]='h00000ea8;  wr_data_rom[ 9313]='h00002094;
    rd_cycle[ 9314] = 1'b0;  wr_cycle[ 9314] = 1'b1;  addr_rom[ 9314]='h0000243c;  wr_data_rom[ 9314]='h000032a9;
    rd_cycle[ 9315] = 1'b0;  wr_cycle[ 9315] = 1'b1;  addr_rom[ 9315]='h00000090;  wr_data_rom[ 9315]='h00000c9f;
    rd_cycle[ 9316] = 1'b1;  wr_cycle[ 9316] = 1'b0;  addr_rom[ 9316]='h00002b78;  wr_data_rom[ 9316]='h00000000;
    rd_cycle[ 9317] = 1'b0;  wr_cycle[ 9317] = 1'b1;  addr_rom[ 9317]='h00002b00;  wr_data_rom[ 9317]='h0000364d;
    rd_cycle[ 9318] = 1'b0;  wr_cycle[ 9318] = 1'b1;  addr_rom[ 9318]='h00003988;  wr_data_rom[ 9318]='h000016b8;
    rd_cycle[ 9319] = 1'b0;  wr_cycle[ 9319] = 1'b1;  addr_rom[ 9319]='h00003f94;  wr_data_rom[ 9319]='h000028eb;
    rd_cycle[ 9320] = 1'b1;  wr_cycle[ 9320] = 1'b0;  addr_rom[ 9320]='h00002170;  wr_data_rom[ 9320]='h00000000;
    rd_cycle[ 9321] = 1'b0;  wr_cycle[ 9321] = 1'b1;  addr_rom[ 9321]='h00000e44;  wr_data_rom[ 9321]='h0000231f;
    rd_cycle[ 9322] = 1'b0;  wr_cycle[ 9322] = 1'b1;  addr_rom[ 9322]='h000029a0;  wr_data_rom[ 9322]='h000033aa;
    rd_cycle[ 9323] = 1'b1;  wr_cycle[ 9323] = 1'b0;  addr_rom[ 9323]='h00000a0c;  wr_data_rom[ 9323]='h00000000;
    rd_cycle[ 9324] = 1'b0;  wr_cycle[ 9324] = 1'b1;  addr_rom[ 9324]='h00001f54;  wr_data_rom[ 9324]='h00002c23;
    rd_cycle[ 9325] = 1'b0;  wr_cycle[ 9325] = 1'b1;  addr_rom[ 9325]='h00000340;  wr_data_rom[ 9325]='h00000f83;
    rd_cycle[ 9326] = 1'b1;  wr_cycle[ 9326] = 1'b0;  addr_rom[ 9326]='h00000484;  wr_data_rom[ 9326]='h00000000;
    rd_cycle[ 9327] = 1'b0;  wr_cycle[ 9327] = 1'b1;  addr_rom[ 9327]='h00003618;  wr_data_rom[ 9327]='h00001ca5;
    rd_cycle[ 9328] = 1'b0;  wr_cycle[ 9328] = 1'b1;  addr_rom[ 9328]='h00002878;  wr_data_rom[ 9328]='h00002211;
    rd_cycle[ 9329] = 1'b0;  wr_cycle[ 9329] = 1'b1;  addr_rom[ 9329]='h000004d4;  wr_data_rom[ 9329]='h000001e0;
    rd_cycle[ 9330] = 1'b1;  wr_cycle[ 9330] = 1'b0;  addr_rom[ 9330]='h00002a14;  wr_data_rom[ 9330]='h00000000;
    rd_cycle[ 9331] = 1'b0;  wr_cycle[ 9331] = 1'b1;  addr_rom[ 9331]='h00003cac;  wr_data_rom[ 9331]='h000033c5;
    rd_cycle[ 9332] = 1'b1;  wr_cycle[ 9332] = 1'b0;  addr_rom[ 9332]='h00002860;  wr_data_rom[ 9332]='h00000000;
    rd_cycle[ 9333] = 1'b0;  wr_cycle[ 9333] = 1'b1;  addr_rom[ 9333]='h00002aec;  wr_data_rom[ 9333]='h0000023d;
    rd_cycle[ 9334] = 1'b0;  wr_cycle[ 9334] = 1'b1;  addr_rom[ 9334]='h00003328;  wr_data_rom[ 9334]='h000002bc;
    rd_cycle[ 9335] = 1'b0;  wr_cycle[ 9335] = 1'b1;  addr_rom[ 9335]='h00003f34;  wr_data_rom[ 9335]='h000014c8;
    rd_cycle[ 9336] = 1'b1;  wr_cycle[ 9336] = 1'b0;  addr_rom[ 9336]='h0000238c;  wr_data_rom[ 9336]='h00000000;
    rd_cycle[ 9337] = 1'b1;  wr_cycle[ 9337] = 1'b0;  addr_rom[ 9337]='h00003544;  wr_data_rom[ 9337]='h00000000;
    rd_cycle[ 9338] = 1'b0;  wr_cycle[ 9338] = 1'b1;  addr_rom[ 9338]='h00002404;  wr_data_rom[ 9338]='h00003a49;
    rd_cycle[ 9339] = 1'b1;  wr_cycle[ 9339] = 1'b0;  addr_rom[ 9339]='h00003980;  wr_data_rom[ 9339]='h00000000;
    rd_cycle[ 9340] = 1'b1;  wr_cycle[ 9340] = 1'b0;  addr_rom[ 9340]='h00000628;  wr_data_rom[ 9340]='h00000000;
    rd_cycle[ 9341] = 1'b1;  wr_cycle[ 9341] = 1'b0;  addr_rom[ 9341]='h00003a08;  wr_data_rom[ 9341]='h00000000;
    rd_cycle[ 9342] = 1'b0;  wr_cycle[ 9342] = 1'b1;  addr_rom[ 9342]='h00000344;  wr_data_rom[ 9342]='h000014f2;
    rd_cycle[ 9343] = 1'b0;  wr_cycle[ 9343] = 1'b1;  addr_rom[ 9343]='h00003928;  wr_data_rom[ 9343]='h00001b02;
    rd_cycle[ 9344] = 1'b0;  wr_cycle[ 9344] = 1'b1;  addr_rom[ 9344]='h00000e60;  wr_data_rom[ 9344]='h000030f6;
    rd_cycle[ 9345] = 1'b0;  wr_cycle[ 9345] = 1'b1;  addr_rom[ 9345]='h00001a08;  wr_data_rom[ 9345]='h00000690;
    rd_cycle[ 9346] = 1'b0;  wr_cycle[ 9346] = 1'b1;  addr_rom[ 9346]='h00003b20;  wr_data_rom[ 9346]='h000001b0;
    rd_cycle[ 9347] = 1'b1;  wr_cycle[ 9347] = 1'b0;  addr_rom[ 9347]='h0000234c;  wr_data_rom[ 9347]='h00000000;
    rd_cycle[ 9348] = 1'b1;  wr_cycle[ 9348] = 1'b0;  addr_rom[ 9348]='h000007bc;  wr_data_rom[ 9348]='h00000000;
    rd_cycle[ 9349] = 1'b0;  wr_cycle[ 9349] = 1'b1;  addr_rom[ 9349]='h000038b4;  wr_data_rom[ 9349]='h00000c2d;
    rd_cycle[ 9350] = 1'b1;  wr_cycle[ 9350] = 1'b0;  addr_rom[ 9350]='h00002754;  wr_data_rom[ 9350]='h00000000;
    rd_cycle[ 9351] = 1'b0;  wr_cycle[ 9351] = 1'b1;  addr_rom[ 9351]='h00002268;  wr_data_rom[ 9351]='h00000ec2;
    rd_cycle[ 9352] = 1'b1;  wr_cycle[ 9352] = 1'b0;  addr_rom[ 9352]='h00002730;  wr_data_rom[ 9352]='h00000000;
    rd_cycle[ 9353] = 1'b0;  wr_cycle[ 9353] = 1'b1;  addr_rom[ 9353]='h00002ce4;  wr_data_rom[ 9353]='h00001a34;
    rd_cycle[ 9354] = 1'b1;  wr_cycle[ 9354] = 1'b0;  addr_rom[ 9354]='h00003818;  wr_data_rom[ 9354]='h00000000;
    rd_cycle[ 9355] = 1'b1;  wr_cycle[ 9355] = 1'b0;  addr_rom[ 9355]='h00003808;  wr_data_rom[ 9355]='h00000000;
    rd_cycle[ 9356] = 1'b0;  wr_cycle[ 9356] = 1'b1;  addr_rom[ 9356]='h0000312c;  wr_data_rom[ 9356]='h000033b2;
    rd_cycle[ 9357] = 1'b0;  wr_cycle[ 9357] = 1'b1;  addr_rom[ 9357]='h00003c84;  wr_data_rom[ 9357]='h00003a3d;
    rd_cycle[ 9358] = 1'b1;  wr_cycle[ 9358] = 1'b0;  addr_rom[ 9358]='h00000208;  wr_data_rom[ 9358]='h00000000;
    rd_cycle[ 9359] = 1'b1;  wr_cycle[ 9359] = 1'b0;  addr_rom[ 9359]='h00003d74;  wr_data_rom[ 9359]='h00000000;
    rd_cycle[ 9360] = 1'b1;  wr_cycle[ 9360] = 1'b0;  addr_rom[ 9360]='h00000108;  wr_data_rom[ 9360]='h00000000;
    rd_cycle[ 9361] = 1'b0;  wr_cycle[ 9361] = 1'b1;  addr_rom[ 9361]='h000027cc;  wr_data_rom[ 9361]='h00001302;
    rd_cycle[ 9362] = 1'b0;  wr_cycle[ 9362] = 1'b1;  addr_rom[ 9362]='h0000197c;  wr_data_rom[ 9362]='h00002d7b;
    rd_cycle[ 9363] = 1'b1;  wr_cycle[ 9363] = 1'b0;  addr_rom[ 9363]='h00001be0;  wr_data_rom[ 9363]='h00000000;
    rd_cycle[ 9364] = 1'b1;  wr_cycle[ 9364] = 1'b0;  addr_rom[ 9364]='h000026d0;  wr_data_rom[ 9364]='h00000000;
    rd_cycle[ 9365] = 1'b0;  wr_cycle[ 9365] = 1'b1;  addr_rom[ 9365]='h00001fa8;  wr_data_rom[ 9365]='h000015d8;
    rd_cycle[ 9366] = 1'b0;  wr_cycle[ 9366] = 1'b1;  addr_rom[ 9366]='h00001d30;  wr_data_rom[ 9366]='h00003940;
    rd_cycle[ 9367] = 1'b0;  wr_cycle[ 9367] = 1'b1;  addr_rom[ 9367]='h00001034;  wr_data_rom[ 9367]='h00001cc6;
    rd_cycle[ 9368] = 1'b1;  wr_cycle[ 9368] = 1'b0;  addr_rom[ 9368]='h00000d60;  wr_data_rom[ 9368]='h00000000;
    rd_cycle[ 9369] = 1'b1;  wr_cycle[ 9369] = 1'b0;  addr_rom[ 9369]='h00000478;  wr_data_rom[ 9369]='h00000000;
    rd_cycle[ 9370] = 1'b0;  wr_cycle[ 9370] = 1'b1;  addr_rom[ 9370]='h000025c0;  wr_data_rom[ 9370]='h00002400;
    rd_cycle[ 9371] = 1'b0;  wr_cycle[ 9371] = 1'b1;  addr_rom[ 9371]='h00003664;  wr_data_rom[ 9371]='h00000d5e;
    rd_cycle[ 9372] = 1'b0;  wr_cycle[ 9372] = 1'b1;  addr_rom[ 9372]='h0000191c;  wr_data_rom[ 9372]='h000016d5;
    rd_cycle[ 9373] = 1'b1;  wr_cycle[ 9373] = 1'b0;  addr_rom[ 9373]='h00002f4c;  wr_data_rom[ 9373]='h00000000;
    rd_cycle[ 9374] = 1'b0;  wr_cycle[ 9374] = 1'b1;  addr_rom[ 9374]='h000002cc;  wr_data_rom[ 9374]='h00002e88;
    rd_cycle[ 9375] = 1'b0;  wr_cycle[ 9375] = 1'b1;  addr_rom[ 9375]='h00000138;  wr_data_rom[ 9375]='h00000432;
    rd_cycle[ 9376] = 1'b0;  wr_cycle[ 9376] = 1'b1;  addr_rom[ 9376]='h000006c8;  wr_data_rom[ 9376]='h00003e80;
    rd_cycle[ 9377] = 1'b1;  wr_cycle[ 9377] = 1'b0;  addr_rom[ 9377]='h0000375c;  wr_data_rom[ 9377]='h00000000;
    rd_cycle[ 9378] = 1'b1;  wr_cycle[ 9378] = 1'b0;  addr_rom[ 9378]='h00002ac8;  wr_data_rom[ 9378]='h00000000;
    rd_cycle[ 9379] = 1'b1;  wr_cycle[ 9379] = 1'b0;  addr_rom[ 9379]='h00000318;  wr_data_rom[ 9379]='h00000000;
    rd_cycle[ 9380] = 1'b0;  wr_cycle[ 9380] = 1'b1;  addr_rom[ 9380]='h000003d8;  wr_data_rom[ 9380]='h000029a0;
    rd_cycle[ 9381] = 1'b1;  wr_cycle[ 9381] = 1'b0;  addr_rom[ 9381]='h000005fc;  wr_data_rom[ 9381]='h00000000;
    rd_cycle[ 9382] = 1'b1;  wr_cycle[ 9382] = 1'b0;  addr_rom[ 9382]='h00003efc;  wr_data_rom[ 9382]='h00000000;
    rd_cycle[ 9383] = 1'b1;  wr_cycle[ 9383] = 1'b0;  addr_rom[ 9383]='h000016c8;  wr_data_rom[ 9383]='h00000000;
    rd_cycle[ 9384] = 1'b0;  wr_cycle[ 9384] = 1'b1;  addr_rom[ 9384]='h00003988;  wr_data_rom[ 9384]='h00000164;
    rd_cycle[ 9385] = 1'b0;  wr_cycle[ 9385] = 1'b1;  addr_rom[ 9385]='h000001e4;  wr_data_rom[ 9385]='h0000151e;
    rd_cycle[ 9386] = 1'b1;  wr_cycle[ 9386] = 1'b0;  addr_rom[ 9386]='h0000046c;  wr_data_rom[ 9386]='h00000000;
    rd_cycle[ 9387] = 1'b0;  wr_cycle[ 9387] = 1'b1;  addr_rom[ 9387]='h00003fd8;  wr_data_rom[ 9387]='h0000105d;
    rd_cycle[ 9388] = 1'b1;  wr_cycle[ 9388] = 1'b0;  addr_rom[ 9388]='h000030e0;  wr_data_rom[ 9388]='h00000000;
    rd_cycle[ 9389] = 1'b0;  wr_cycle[ 9389] = 1'b1;  addr_rom[ 9389]='h00002010;  wr_data_rom[ 9389]='h00002d97;
    rd_cycle[ 9390] = 1'b1;  wr_cycle[ 9390] = 1'b0;  addr_rom[ 9390]='h00001d60;  wr_data_rom[ 9390]='h00000000;
    rd_cycle[ 9391] = 1'b0;  wr_cycle[ 9391] = 1'b1;  addr_rom[ 9391]='h000024bc;  wr_data_rom[ 9391]='h00002ebe;
    rd_cycle[ 9392] = 1'b1;  wr_cycle[ 9392] = 1'b0;  addr_rom[ 9392]='h00003064;  wr_data_rom[ 9392]='h00000000;
    rd_cycle[ 9393] = 1'b0;  wr_cycle[ 9393] = 1'b1;  addr_rom[ 9393]='h00003de0;  wr_data_rom[ 9393]='h00003b99;
    rd_cycle[ 9394] = 1'b1;  wr_cycle[ 9394] = 1'b0;  addr_rom[ 9394]='h000037f0;  wr_data_rom[ 9394]='h00000000;
    rd_cycle[ 9395] = 1'b1;  wr_cycle[ 9395] = 1'b0;  addr_rom[ 9395]='h000019f0;  wr_data_rom[ 9395]='h00000000;
    rd_cycle[ 9396] = 1'b0;  wr_cycle[ 9396] = 1'b1;  addr_rom[ 9396]='h00002674;  wr_data_rom[ 9396]='h00001587;
    rd_cycle[ 9397] = 1'b0;  wr_cycle[ 9397] = 1'b1;  addr_rom[ 9397]='h00000eec;  wr_data_rom[ 9397]='h000039d2;
    rd_cycle[ 9398] = 1'b0;  wr_cycle[ 9398] = 1'b1;  addr_rom[ 9398]='h0000264c;  wr_data_rom[ 9398]='h00002358;
    rd_cycle[ 9399] = 1'b1;  wr_cycle[ 9399] = 1'b0;  addr_rom[ 9399]='h00001f4c;  wr_data_rom[ 9399]='h00000000;
    rd_cycle[ 9400] = 1'b1;  wr_cycle[ 9400] = 1'b0;  addr_rom[ 9400]='h00002d70;  wr_data_rom[ 9400]='h00000000;
    rd_cycle[ 9401] = 1'b0;  wr_cycle[ 9401] = 1'b1;  addr_rom[ 9401]='h0000188c;  wr_data_rom[ 9401]='h000009bd;
    rd_cycle[ 9402] = 1'b1;  wr_cycle[ 9402] = 1'b0;  addr_rom[ 9402]='h0000355c;  wr_data_rom[ 9402]='h00000000;
    rd_cycle[ 9403] = 1'b0;  wr_cycle[ 9403] = 1'b1;  addr_rom[ 9403]='h00003304;  wr_data_rom[ 9403]='h0000397c;
    rd_cycle[ 9404] = 1'b1;  wr_cycle[ 9404] = 1'b0;  addr_rom[ 9404]='h00002f68;  wr_data_rom[ 9404]='h00000000;
    rd_cycle[ 9405] = 1'b1;  wr_cycle[ 9405] = 1'b0;  addr_rom[ 9405]='h00003384;  wr_data_rom[ 9405]='h00000000;
    rd_cycle[ 9406] = 1'b1;  wr_cycle[ 9406] = 1'b0;  addr_rom[ 9406]='h00001ab0;  wr_data_rom[ 9406]='h00000000;
    rd_cycle[ 9407] = 1'b0;  wr_cycle[ 9407] = 1'b1;  addr_rom[ 9407]='h00003374;  wr_data_rom[ 9407]='h00001ca9;
    rd_cycle[ 9408] = 1'b0;  wr_cycle[ 9408] = 1'b1;  addr_rom[ 9408]='h00001340;  wr_data_rom[ 9408]='h00003534;
    rd_cycle[ 9409] = 1'b0;  wr_cycle[ 9409] = 1'b1;  addr_rom[ 9409]='h000031d8;  wr_data_rom[ 9409]='h00001ad5;
    rd_cycle[ 9410] = 1'b0;  wr_cycle[ 9410] = 1'b1;  addr_rom[ 9410]='h000025ec;  wr_data_rom[ 9410]='h000019cf;
    rd_cycle[ 9411] = 1'b0;  wr_cycle[ 9411] = 1'b1;  addr_rom[ 9411]='h00003ec0;  wr_data_rom[ 9411]='h00000908;
    rd_cycle[ 9412] = 1'b0;  wr_cycle[ 9412] = 1'b1;  addr_rom[ 9412]='h00003d10;  wr_data_rom[ 9412]='h00001992;
    rd_cycle[ 9413] = 1'b1;  wr_cycle[ 9413] = 1'b0;  addr_rom[ 9413]='h000024f8;  wr_data_rom[ 9413]='h00000000;
    rd_cycle[ 9414] = 1'b1;  wr_cycle[ 9414] = 1'b0;  addr_rom[ 9414]='h00000ef0;  wr_data_rom[ 9414]='h00000000;
    rd_cycle[ 9415] = 1'b1;  wr_cycle[ 9415] = 1'b0;  addr_rom[ 9415]='h00001b50;  wr_data_rom[ 9415]='h00000000;
    rd_cycle[ 9416] = 1'b0;  wr_cycle[ 9416] = 1'b1;  addr_rom[ 9416]='h00001368;  wr_data_rom[ 9416]='h00001c56;
    rd_cycle[ 9417] = 1'b1;  wr_cycle[ 9417] = 1'b0;  addr_rom[ 9417]='h00002d0c;  wr_data_rom[ 9417]='h00000000;
    rd_cycle[ 9418] = 1'b1;  wr_cycle[ 9418] = 1'b0;  addr_rom[ 9418]='h0000059c;  wr_data_rom[ 9418]='h00000000;
    rd_cycle[ 9419] = 1'b1;  wr_cycle[ 9419] = 1'b0;  addr_rom[ 9419]='h000015c4;  wr_data_rom[ 9419]='h00000000;
    rd_cycle[ 9420] = 1'b0;  wr_cycle[ 9420] = 1'b1;  addr_rom[ 9420]='h00001e0c;  wr_data_rom[ 9420]='h00003ebf;
    rd_cycle[ 9421] = 1'b0;  wr_cycle[ 9421] = 1'b1;  addr_rom[ 9421]='h00000d54;  wr_data_rom[ 9421]='h00000988;
    rd_cycle[ 9422] = 1'b1;  wr_cycle[ 9422] = 1'b0;  addr_rom[ 9422]='h00002c64;  wr_data_rom[ 9422]='h00000000;
    rd_cycle[ 9423] = 1'b0;  wr_cycle[ 9423] = 1'b1;  addr_rom[ 9423]='h00000774;  wr_data_rom[ 9423]='h00002c8d;
    rd_cycle[ 9424] = 1'b1;  wr_cycle[ 9424] = 1'b0;  addr_rom[ 9424]='h0000210c;  wr_data_rom[ 9424]='h00000000;
    rd_cycle[ 9425] = 1'b1;  wr_cycle[ 9425] = 1'b0;  addr_rom[ 9425]='h00003d90;  wr_data_rom[ 9425]='h00000000;
    rd_cycle[ 9426] = 1'b0;  wr_cycle[ 9426] = 1'b1;  addr_rom[ 9426]='h000004a0;  wr_data_rom[ 9426]='h000035c6;
    rd_cycle[ 9427] = 1'b1;  wr_cycle[ 9427] = 1'b0;  addr_rom[ 9427]='h00000de0;  wr_data_rom[ 9427]='h00000000;
    rd_cycle[ 9428] = 1'b1;  wr_cycle[ 9428] = 1'b0;  addr_rom[ 9428]='h0000240c;  wr_data_rom[ 9428]='h00000000;
    rd_cycle[ 9429] = 1'b1;  wr_cycle[ 9429] = 1'b0;  addr_rom[ 9429]='h00003d34;  wr_data_rom[ 9429]='h00000000;
    rd_cycle[ 9430] = 1'b1;  wr_cycle[ 9430] = 1'b0;  addr_rom[ 9430]='h000033a8;  wr_data_rom[ 9430]='h00000000;
    rd_cycle[ 9431] = 1'b0;  wr_cycle[ 9431] = 1'b1;  addr_rom[ 9431]='h00000d70;  wr_data_rom[ 9431]='h0000109a;
    rd_cycle[ 9432] = 1'b1;  wr_cycle[ 9432] = 1'b0;  addr_rom[ 9432]='h00002b94;  wr_data_rom[ 9432]='h00000000;
    rd_cycle[ 9433] = 1'b0;  wr_cycle[ 9433] = 1'b1;  addr_rom[ 9433]='h000027d0;  wr_data_rom[ 9433]='h000037fe;
    rd_cycle[ 9434] = 1'b0;  wr_cycle[ 9434] = 1'b1;  addr_rom[ 9434]='h00003488;  wr_data_rom[ 9434]='h00002a0c;
    rd_cycle[ 9435] = 1'b1;  wr_cycle[ 9435] = 1'b0;  addr_rom[ 9435]='h00001388;  wr_data_rom[ 9435]='h00000000;
    rd_cycle[ 9436] = 1'b0;  wr_cycle[ 9436] = 1'b1;  addr_rom[ 9436]='h0000273c;  wr_data_rom[ 9436]='h00001073;
    rd_cycle[ 9437] = 1'b0;  wr_cycle[ 9437] = 1'b1;  addr_rom[ 9437]='h000006b4;  wr_data_rom[ 9437]='h00000b69;
    rd_cycle[ 9438] = 1'b1;  wr_cycle[ 9438] = 1'b0;  addr_rom[ 9438]='h000033f0;  wr_data_rom[ 9438]='h00000000;
    rd_cycle[ 9439] = 1'b1;  wr_cycle[ 9439] = 1'b0;  addr_rom[ 9439]='h00000444;  wr_data_rom[ 9439]='h00000000;
    rd_cycle[ 9440] = 1'b1;  wr_cycle[ 9440] = 1'b0;  addr_rom[ 9440]='h0000166c;  wr_data_rom[ 9440]='h00000000;
    rd_cycle[ 9441] = 1'b1;  wr_cycle[ 9441] = 1'b0;  addr_rom[ 9441]='h00001928;  wr_data_rom[ 9441]='h00000000;
    rd_cycle[ 9442] = 1'b1;  wr_cycle[ 9442] = 1'b0;  addr_rom[ 9442]='h0000357c;  wr_data_rom[ 9442]='h00000000;
    rd_cycle[ 9443] = 1'b1;  wr_cycle[ 9443] = 1'b0;  addr_rom[ 9443]='h0000016c;  wr_data_rom[ 9443]='h00000000;
    rd_cycle[ 9444] = 1'b0;  wr_cycle[ 9444] = 1'b1;  addr_rom[ 9444]='h00003448;  wr_data_rom[ 9444]='h00001c6e;
    rd_cycle[ 9445] = 1'b0;  wr_cycle[ 9445] = 1'b1;  addr_rom[ 9445]='h00000bb0;  wr_data_rom[ 9445]='h00003d74;
    rd_cycle[ 9446] = 1'b0;  wr_cycle[ 9446] = 1'b1;  addr_rom[ 9446]='h00003b84;  wr_data_rom[ 9446]='h00000709;
    rd_cycle[ 9447] = 1'b1;  wr_cycle[ 9447] = 1'b0;  addr_rom[ 9447]='h000018d8;  wr_data_rom[ 9447]='h00000000;
    rd_cycle[ 9448] = 1'b0;  wr_cycle[ 9448] = 1'b1;  addr_rom[ 9448]='h00000294;  wr_data_rom[ 9448]='h00003416;
    rd_cycle[ 9449] = 1'b1;  wr_cycle[ 9449] = 1'b0;  addr_rom[ 9449]='h00002d50;  wr_data_rom[ 9449]='h00000000;
    rd_cycle[ 9450] = 1'b1;  wr_cycle[ 9450] = 1'b0;  addr_rom[ 9450]='h00001774;  wr_data_rom[ 9450]='h00000000;
    rd_cycle[ 9451] = 1'b0;  wr_cycle[ 9451] = 1'b1;  addr_rom[ 9451]='h000009cc;  wr_data_rom[ 9451]='h000017c0;
    rd_cycle[ 9452] = 1'b1;  wr_cycle[ 9452] = 1'b0;  addr_rom[ 9452]='h00001680;  wr_data_rom[ 9452]='h00000000;
    rd_cycle[ 9453] = 1'b1;  wr_cycle[ 9453] = 1'b0;  addr_rom[ 9453]='h00003e44;  wr_data_rom[ 9453]='h00000000;
    rd_cycle[ 9454] = 1'b1;  wr_cycle[ 9454] = 1'b0;  addr_rom[ 9454]='h00002bdc;  wr_data_rom[ 9454]='h00000000;
    rd_cycle[ 9455] = 1'b0;  wr_cycle[ 9455] = 1'b1;  addr_rom[ 9455]='h000009bc;  wr_data_rom[ 9455]='h0000326f;
    rd_cycle[ 9456] = 1'b1;  wr_cycle[ 9456] = 1'b0;  addr_rom[ 9456]='h000019f8;  wr_data_rom[ 9456]='h00000000;
    rd_cycle[ 9457] = 1'b0;  wr_cycle[ 9457] = 1'b1;  addr_rom[ 9457]='h00000340;  wr_data_rom[ 9457]='h0000168d;
    rd_cycle[ 9458] = 1'b0;  wr_cycle[ 9458] = 1'b1;  addr_rom[ 9458]='h00003028;  wr_data_rom[ 9458]='h000001b8;
    rd_cycle[ 9459] = 1'b0;  wr_cycle[ 9459] = 1'b1;  addr_rom[ 9459]='h00000680;  wr_data_rom[ 9459]='h000001f0;
    rd_cycle[ 9460] = 1'b0;  wr_cycle[ 9460] = 1'b1;  addr_rom[ 9460]='h0000104c;  wr_data_rom[ 9460]='h00001c2f;
    rd_cycle[ 9461] = 1'b1;  wr_cycle[ 9461] = 1'b0;  addr_rom[ 9461]='h0000195c;  wr_data_rom[ 9461]='h00000000;
    rd_cycle[ 9462] = 1'b1;  wr_cycle[ 9462] = 1'b0;  addr_rom[ 9462]='h000037c0;  wr_data_rom[ 9462]='h00000000;
    rd_cycle[ 9463] = 1'b1;  wr_cycle[ 9463] = 1'b0;  addr_rom[ 9463]='h0000043c;  wr_data_rom[ 9463]='h00000000;
    rd_cycle[ 9464] = 1'b0;  wr_cycle[ 9464] = 1'b1;  addr_rom[ 9464]='h00002414;  wr_data_rom[ 9464]='h000003fe;
    rd_cycle[ 9465] = 1'b0;  wr_cycle[ 9465] = 1'b1;  addr_rom[ 9465]='h00001910;  wr_data_rom[ 9465]='h000009a6;
    rd_cycle[ 9466] = 1'b0;  wr_cycle[ 9466] = 1'b1;  addr_rom[ 9466]='h00001228;  wr_data_rom[ 9466]='h0000143d;
    rd_cycle[ 9467] = 1'b0;  wr_cycle[ 9467] = 1'b1;  addr_rom[ 9467]='h000010f8;  wr_data_rom[ 9467]='h00002bee;
    rd_cycle[ 9468] = 1'b1;  wr_cycle[ 9468] = 1'b0;  addr_rom[ 9468]='h000026f4;  wr_data_rom[ 9468]='h00000000;
    rd_cycle[ 9469] = 1'b0;  wr_cycle[ 9469] = 1'b1;  addr_rom[ 9469]='h00003ed0;  wr_data_rom[ 9469]='h0000015e;
    rd_cycle[ 9470] = 1'b0;  wr_cycle[ 9470] = 1'b1;  addr_rom[ 9470]='h00001884;  wr_data_rom[ 9470]='h000017ef;
    rd_cycle[ 9471] = 1'b0;  wr_cycle[ 9471] = 1'b1;  addr_rom[ 9471]='h0000251c;  wr_data_rom[ 9471]='h00002c08;
    rd_cycle[ 9472] = 1'b0;  wr_cycle[ 9472] = 1'b1;  addr_rom[ 9472]='h00002224;  wr_data_rom[ 9472]='h00000326;
    rd_cycle[ 9473] = 1'b0;  wr_cycle[ 9473] = 1'b1;  addr_rom[ 9473]='h00000f50;  wr_data_rom[ 9473]='h0000158e;
    rd_cycle[ 9474] = 1'b1;  wr_cycle[ 9474] = 1'b0;  addr_rom[ 9474]='h00002a5c;  wr_data_rom[ 9474]='h00000000;
    rd_cycle[ 9475] = 1'b1;  wr_cycle[ 9475] = 1'b0;  addr_rom[ 9475]='h00000234;  wr_data_rom[ 9475]='h00000000;
    rd_cycle[ 9476] = 1'b0;  wr_cycle[ 9476] = 1'b1;  addr_rom[ 9476]='h00001ccc;  wr_data_rom[ 9476]='h00001536;
    rd_cycle[ 9477] = 1'b0;  wr_cycle[ 9477] = 1'b1;  addr_rom[ 9477]='h0000063c;  wr_data_rom[ 9477]='h00001deb;
    rd_cycle[ 9478] = 1'b0;  wr_cycle[ 9478] = 1'b1;  addr_rom[ 9478]='h00001500;  wr_data_rom[ 9478]='h00002d08;
    rd_cycle[ 9479] = 1'b1;  wr_cycle[ 9479] = 1'b0;  addr_rom[ 9479]='h000033d4;  wr_data_rom[ 9479]='h00000000;
    rd_cycle[ 9480] = 1'b1;  wr_cycle[ 9480] = 1'b0;  addr_rom[ 9480]='h00003628;  wr_data_rom[ 9480]='h00000000;
    rd_cycle[ 9481] = 1'b0;  wr_cycle[ 9481] = 1'b1;  addr_rom[ 9481]='h00000934;  wr_data_rom[ 9481]='h0000260f;
    rd_cycle[ 9482] = 1'b1;  wr_cycle[ 9482] = 1'b0;  addr_rom[ 9482]='h00000130;  wr_data_rom[ 9482]='h00000000;
    rd_cycle[ 9483] = 1'b0;  wr_cycle[ 9483] = 1'b1;  addr_rom[ 9483]='h00001084;  wr_data_rom[ 9483]='h0000196f;
    rd_cycle[ 9484] = 1'b1;  wr_cycle[ 9484] = 1'b0;  addr_rom[ 9484]='h00001558;  wr_data_rom[ 9484]='h00000000;
    rd_cycle[ 9485] = 1'b1;  wr_cycle[ 9485] = 1'b0;  addr_rom[ 9485]='h00000688;  wr_data_rom[ 9485]='h00000000;
    rd_cycle[ 9486] = 1'b1;  wr_cycle[ 9486] = 1'b0;  addr_rom[ 9486]='h00003214;  wr_data_rom[ 9486]='h00000000;
    rd_cycle[ 9487] = 1'b0;  wr_cycle[ 9487] = 1'b1;  addr_rom[ 9487]='h00003e94;  wr_data_rom[ 9487]='h00001798;
    rd_cycle[ 9488] = 1'b1;  wr_cycle[ 9488] = 1'b0;  addr_rom[ 9488]='h00002348;  wr_data_rom[ 9488]='h00000000;
    rd_cycle[ 9489] = 1'b1;  wr_cycle[ 9489] = 1'b0;  addr_rom[ 9489]='h00002334;  wr_data_rom[ 9489]='h00000000;
    rd_cycle[ 9490] = 1'b1;  wr_cycle[ 9490] = 1'b0;  addr_rom[ 9490]='h00003358;  wr_data_rom[ 9490]='h00000000;
    rd_cycle[ 9491] = 1'b1;  wr_cycle[ 9491] = 1'b0;  addr_rom[ 9491]='h0000225c;  wr_data_rom[ 9491]='h00000000;
    rd_cycle[ 9492] = 1'b1;  wr_cycle[ 9492] = 1'b0;  addr_rom[ 9492]='h0000270c;  wr_data_rom[ 9492]='h00000000;
    rd_cycle[ 9493] = 1'b0;  wr_cycle[ 9493] = 1'b1;  addr_rom[ 9493]='h000025b8;  wr_data_rom[ 9493]='h00000068;
    rd_cycle[ 9494] = 1'b0;  wr_cycle[ 9494] = 1'b1;  addr_rom[ 9494]='h00002e08;  wr_data_rom[ 9494]='h00001297;
    rd_cycle[ 9495] = 1'b1;  wr_cycle[ 9495] = 1'b0;  addr_rom[ 9495]='h000011ac;  wr_data_rom[ 9495]='h00000000;
    rd_cycle[ 9496] = 1'b1;  wr_cycle[ 9496] = 1'b0;  addr_rom[ 9496]='h00000a04;  wr_data_rom[ 9496]='h00000000;
    rd_cycle[ 9497] = 1'b1;  wr_cycle[ 9497] = 1'b0;  addr_rom[ 9497]='h000017d4;  wr_data_rom[ 9497]='h00000000;
    rd_cycle[ 9498] = 1'b1;  wr_cycle[ 9498] = 1'b0;  addr_rom[ 9498]='h00001744;  wr_data_rom[ 9498]='h00000000;
    rd_cycle[ 9499] = 1'b0;  wr_cycle[ 9499] = 1'b1;  addr_rom[ 9499]='h000004c4;  wr_data_rom[ 9499]='h00000cea;
    rd_cycle[ 9500] = 1'b1;  wr_cycle[ 9500] = 1'b0;  addr_rom[ 9500]='h00002c70;  wr_data_rom[ 9500]='h00000000;
    rd_cycle[ 9501] = 1'b1;  wr_cycle[ 9501] = 1'b0;  addr_rom[ 9501]='h00002dbc;  wr_data_rom[ 9501]='h00000000;
    rd_cycle[ 9502] = 1'b1;  wr_cycle[ 9502] = 1'b0;  addr_rom[ 9502]='h00003430;  wr_data_rom[ 9502]='h00000000;
    rd_cycle[ 9503] = 1'b1;  wr_cycle[ 9503] = 1'b0;  addr_rom[ 9503]='h00003c2c;  wr_data_rom[ 9503]='h00000000;
    rd_cycle[ 9504] = 1'b1;  wr_cycle[ 9504] = 1'b0;  addr_rom[ 9504]='h00003610;  wr_data_rom[ 9504]='h00000000;
    rd_cycle[ 9505] = 1'b1;  wr_cycle[ 9505] = 1'b0;  addr_rom[ 9505]='h00001c50;  wr_data_rom[ 9505]='h00000000;
    rd_cycle[ 9506] = 1'b0;  wr_cycle[ 9506] = 1'b1;  addr_rom[ 9506]='h00003bc4;  wr_data_rom[ 9506]='h00002c34;
    rd_cycle[ 9507] = 1'b1;  wr_cycle[ 9507] = 1'b0;  addr_rom[ 9507]='h00003924;  wr_data_rom[ 9507]='h00000000;
    rd_cycle[ 9508] = 1'b1;  wr_cycle[ 9508] = 1'b0;  addr_rom[ 9508]='h00001758;  wr_data_rom[ 9508]='h00000000;
    rd_cycle[ 9509] = 1'b1;  wr_cycle[ 9509] = 1'b0;  addr_rom[ 9509]='h00002664;  wr_data_rom[ 9509]='h00000000;
    rd_cycle[ 9510] = 1'b0;  wr_cycle[ 9510] = 1'b1;  addr_rom[ 9510]='h00001108;  wr_data_rom[ 9510]='h0000166b;
    rd_cycle[ 9511] = 1'b1;  wr_cycle[ 9511] = 1'b0;  addr_rom[ 9511]='h00002c70;  wr_data_rom[ 9511]='h00000000;
    rd_cycle[ 9512] = 1'b0;  wr_cycle[ 9512] = 1'b1;  addr_rom[ 9512]='h000000e4;  wr_data_rom[ 9512]='h00001caa;
    rd_cycle[ 9513] = 1'b0;  wr_cycle[ 9513] = 1'b1;  addr_rom[ 9513]='h0000313c;  wr_data_rom[ 9513]='h000018a5;
    rd_cycle[ 9514] = 1'b1;  wr_cycle[ 9514] = 1'b0;  addr_rom[ 9514]='h00001044;  wr_data_rom[ 9514]='h00000000;
    rd_cycle[ 9515] = 1'b1;  wr_cycle[ 9515] = 1'b0;  addr_rom[ 9515]='h00001478;  wr_data_rom[ 9515]='h00000000;
    rd_cycle[ 9516] = 1'b1;  wr_cycle[ 9516] = 1'b0;  addr_rom[ 9516]='h000001dc;  wr_data_rom[ 9516]='h00000000;
    rd_cycle[ 9517] = 1'b0;  wr_cycle[ 9517] = 1'b1;  addr_rom[ 9517]='h000031f4;  wr_data_rom[ 9517]='h000023cf;
    rd_cycle[ 9518] = 1'b0;  wr_cycle[ 9518] = 1'b1;  addr_rom[ 9518]='h00003fe0;  wr_data_rom[ 9518]='h00001b95;
    rd_cycle[ 9519] = 1'b1;  wr_cycle[ 9519] = 1'b0;  addr_rom[ 9519]='h00001378;  wr_data_rom[ 9519]='h00000000;
    rd_cycle[ 9520] = 1'b0;  wr_cycle[ 9520] = 1'b1;  addr_rom[ 9520]='h00000540;  wr_data_rom[ 9520]='h0000288e;
    rd_cycle[ 9521] = 1'b1;  wr_cycle[ 9521] = 1'b0;  addr_rom[ 9521]='h000029d0;  wr_data_rom[ 9521]='h00000000;
    rd_cycle[ 9522] = 1'b0;  wr_cycle[ 9522] = 1'b1;  addr_rom[ 9522]='h00000474;  wr_data_rom[ 9522]='h00003cd1;
    rd_cycle[ 9523] = 1'b1;  wr_cycle[ 9523] = 1'b0;  addr_rom[ 9523]='h00001a34;  wr_data_rom[ 9523]='h00000000;
    rd_cycle[ 9524] = 1'b0;  wr_cycle[ 9524] = 1'b1;  addr_rom[ 9524]='h00003278;  wr_data_rom[ 9524]='h0000275f;
    rd_cycle[ 9525] = 1'b1;  wr_cycle[ 9525] = 1'b0;  addr_rom[ 9525]='h00001438;  wr_data_rom[ 9525]='h00000000;
    rd_cycle[ 9526] = 1'b1;  wr_cycle[ 9526] = 1'b0;  addr_rom[ 9526]='h00000dec;  wr_data_rom[ 9526]='h00000000;
    rd_cycle[ 9527] = 1'b0;  wr_cycle[ 9527] = 1'b1;  addr_rom[ 9527]='h00001be4;  wr_data_rom[ 9527]='h00003490;
    rd_cycle[ 9528] = 1'b1;  wr_cycle[ 9528] = 1'b0;  addr_rom[ 9528]='h00001120;  wr_data_rom[ 9528]='h00000000;
    rd_cycle[ 9529] = 1'b1;  wr_cycle[ 9529] = 1'b0;  addr_rom[ 9529]='h00001d58;  wr_data_rom[ 9529]='h00000000;
    rd_cycle[ 9530] = 1'b0;  wr_cycle[ 9530] = 1'b1;  addr_rom[ 9530]='h000037e0;  wr_data_rom[ 9530]='h00000f21;
    rd_cycle[ 9531] = 1'b1;  wr_cycle[ 9531] = 1'b0;  addr_rom[ 9531]='h00001154;  wr_data_rom[ 9531]='h00000000;
    rd_cycle[ 9532] = 1'b0;  wr_cycle[ 9532] = 1'b1;  addr_rom[ 9532]='h00002fd8;  wr_data_rom[ 9532]='h0000276e;
    rd_cycle[ 9533] = 1'b0;  wr_cycle[ 9533] = 1'b1;  addr_rom[ 9533]='h00002fd4;  wr_data_rom[ 9533]='h0000353d;
    rd_cycle[ 9534] = 1'b0;  wr_cycle[ 9534] = 1'b1;  addr_rom[ 9534]='h00001464;  wr_data_rom[ 9534]='h0000194a;
    rd_cycle[ 9535] = 1'b1;  wr_cycle[ 9535] = 1'b0;  addr_rom[ 9535]='h00003938;  wr_data_rom[ 9535]='h00000000;
    rd_cycle[ 9536] = 1'b0;  wr_cycle[ 9536] = 1'b1;  addr_rom[ 9536]='h000012bc;  wr_data_rom[ 9536]='h00001cb7;
    rd_cycle[ 9537] = 1'b1;  wr_cycle[ 9537] = 1'b0;  addr_rom[ 9537]='h00001c1c;  wr_data_rom[ 9537]='h00000000;
    rd_cycle[ 9538] = 1'b1;  wr_cycle[ 9538] = 1'b0;  addr_rom[ 9538]='h00000dbc;  wr_data_rom[ 9538]='h00000000;
    rd_cycle[ 9539] = 1'b1;  wr_cycle[ 9539] = 1'b0;  addr_rom[ 9539]='h00000864;  wr_data_rom[ 9539]='h00000000;
    rd_cycle[ 9540] = 1'b0;  wr_cycle[ 9540] = 1'b1;  addr_rom[ 9540]='h00001440;  wr_data_rom[ 9540]='h00003e28;
    rd_cycle[ 9541] = 1'b0;  wr_cycle[ 9541] = 1'b1;  addr_rom[ 9541]='h00001cbc;  wr_data_rom[ 9541]='h00002bb2;
    rd_cycle[ 9542] = 1'b0;  wr_cycle[ 9542] = 1'b1;  addr_rom[ 9542]='h00001c60;  wr_data_rom[ 9542]='h00002906;
    rd_cycle[ 9543] = 1'b0;  wr_cycle[ 9543] = 1'b1;  addr_rom[ 9543]='h0000155c;  wr_data_rom[ 9543]='h00001188;
    rd_cycle[ 9544] = 1'b1;  wr_cycle[ 9544] = 1'b0;  addr_rom[ 9544]='h00002710;  wr_data_rom[ 9544]='h00000000;
    rd_cycle[ 9545] = 1'b1;  wr_cycle[ 9545] = 1'b0;  addr_rom[ 9545]='h00003504;  wr_data_rom[ 9545]='h00000000;
    rd_cycle[ 9546] = 1'b1;  wr_cycle[ 9546] = 1'b0;  addr_rom[ 9546]='h0000200c;  wr_data_rom[ 9546]='h00000000;
    rd_cycle[ 9547] = 1'b0;  wr_cycle[ 9547] = 1'b1;  addr_rom[ 9547]='h000006f0;  wr_data_rom[ 9547]='h0000047d;
    rd_cycle[ 9548] = 1'b0;  wr_cycle[ 9548] = 1'b1;  addr_rom[ 9548]='h000017a0;  wr_data_rom[ 9548]='h0000020b;
    rd_cycle[ 9549] = 1'b0;  wr_cycle[ 9549] = 1'b1;  addr_rom[ 9549]='h00003e4c;  wr_data_rom[ 9549]='h0000248e;
    rd_cycle[ 9550] = 1'b0;  wr_cycle[ 9550] = 1'b1;  addr_rom[ 9550]='h000014ac;  wr_data_rom[ 9550]='h00000d02;
    rd_cycle[ 9551] = 1'b0;  wr_cycle[ 9551] = 1'b1;  addr_rom[ 9551]='h000028e4;  wr_data_rom[ 9551]='h000033a0;
    rd_cycle[ 9552] = 1'b1;  wr_cycle[ 9552] = 1'b0;  addr_rom[ 9552]='h000008d0;  wr_data_rom[ 9552]='h00000000;
    rd_cycle[ 9553] = 1'b0;  wr_cycle[ 9553] = 1'b1;  addr_rom[ 9553]='h00001120;  wr_data_rom[ 9553]='h0000069b;
    rd_cycle[ 9554] = 1'b1;  wr_cycle[ 9554] = 1'b0;  addr_rom[ 9554]='h0000073c;  wr_data_rom[ 9554]='h00000000;
    rd_cycle[ 9555] = 1'b0;  wr_cycle[ 9555] = 1'b1;  addr_rom[ 9555]='h000004c8;  wr_data_rom[ 9555]='h00001a9b;
    rd_cycle[ 9556] = 1'b0;  wr_cycle[ 9556] = 1'b1;  addr_rom[ 9556]='h00003dec;  wr_data_rom[ 9556]='h0000268d;
    rd_cycle[ 9557] = 1'b1;  wr_cycle[ 9557] = 1'b0;  addr_rom[ 9557]='h00000f84;  wr_data_rom[ 9557]='h00000000;
    rd_cycle[ 9558] = 1'b0;  wr_cycle[ 9558] = 1'b1;  addr_rom[ 9558]='h000007d0;  wr_data_rom[ 9558]='h000039e7;
    rd_cycle[ 9559] = 1'b0;  wr_cycle[ 9559] = 1'b1;  addr_rom[ 9559]='h00002cdc;  wr_data_rom[ 9559]='h00001ef8;
    rd_cycle[ 9560] = 1'b0;  wr_cycle[ 9560] = 1'b1;  addr_rom[ 9560]='h00003614;  wr_data_rom[ 9560]='h00000121;
    rd_cycle[ 9561] = 1'b0;  wr_cycle[ 9561] = 1'b1;  addr_rom[ 9561]='h00003bb8;  wr_data_rom[ 9561]='h00002af8;
    rd_cycle[ 9562] = 1'b0;  wr_cycle[ 9562] = 1'b1;  addr_rom[ 9562]='h00000acc;  wr_data_rom[ 9562]='h00000c24;
    rd_cycle[ 9563] = 1'b1;  wr_cycle[ 9563] = 1'b0;  addr_rom[ 9563]='h00002368;  wr_data_rom[ 9563]='h00000000;
    rd_cycle[ 9564] = 1'b1;  wr_cycle[ 9564] = 1'b0;  addr_rom[ 9564]='h00000878;  wr_data_rom[ 9564]='h00000000;
    rd_cycle[ 9565] = 1'b0;  wr_cycle[ 9565] = 1'b1;  addr_rom[ 9565]='h0000267c;  wr_data_rom[ 9565]='h00000a4b;
    rd_cycle[ 9566] = 1'b1;  wr_cycle[ 9566] = 1'b0;  addr_rom[ 9566]='h000018dc;  wr_data_rom[ 9566]='h00000000;
    rd_cycle[ 9567] = 1'b1;  wr_cycle[ 9567] = 1'b0;  addr_rom[ 9567]='h00001058;  wr_data_rom[ 9567]='h00000000;
    rd_cycle[ 9568] = 1'b1;  wr_cycle[ 9568] = 1'b0;  addr_rom[ 9568]='h0000223c;  wr_data_rom[ 9568]='h00000000;
    rd_cycle[ 9569] = 1'b1;  wr_cycle[ 9569] = 1'b0;  addr_rom[ 9569]='h00001a1c;  wr_data_rom[ 9569]='h00000000;
    rd_cycle[ 9570] = 1'b1;  wr_cycle[ 9570] = 1'b0;  addr_rom[ 9570]='h00001f68;  wr_data_rom[ 9570]='h00000000;
    rd_cycle[ 9571] = 1'b0;  wr_cycle[ 9571] = 1'b1;  addr_rom[ 9571]='h000000b8;  wr_data_rom[ 9571]='h00002c91;
    rd_cycle[ 9572] = 1'b0;  wr_cycle[ 9572] = 1'b1;  addr_rom[ 9572]='h00003b48;  wr_data_rom[ 9572]='h00001bcb;
    rd_cycle[ 9573] = 1'b1;  wr_cycle[ 9573] = 1'b0;  addr_rom[ 9573]='h000039a4;  wr_data_rom[ 9573]='h00000000;
    rd_cycle[ 9574] = 1'b0;  wr_cycle[ 9574] = 1'b1;  addr_rom[ 9574]='h00000b38;  wr_data_rom[ 9574]='h00003708;
    rd_cycle[ 9575] = 1'b0;  wr_cycle[ 9575] = 1'b1;  addr_rom[ 9575]='h00003af0;  wr_data_rom[ 9575]='h00001686;
    rd_cycle[ 9576] = 1'b0;  wr_cycle[ 9576] = 1'b1;  addr_rom[ 9576]='h000023c8;  wr_data_rom[ 9576]='h00000c06;
    rd_cycle[ 9577] = 1'b0;  wr_cycle[ 9577] = 1'b1;  addr_rom[ 9577]='h00000328;  wr_data_rom[ 9577]='h00000490;
    rd_cycle[ 9578] = 1'b1;  wr_cycle[ 9578] = 1'b0;  addr_rom[ 9578]='h0000399c;  wr_data_rom[ 9578]='h00000000;
    rd_cycle[ 9579] = 1'b0;  wr_cycle[ 9579] = 1'b1;  addr_rom[ 9579]='h000034a0;  wr_data_rom[ 9579]='h0000203c;
    rd_cycle[ 9580] = 1'b1;  wr_cycle[ 9580] = 1'b0;  addr_rom[ 9580]='h000000ac;  wr_data_rom[ 9580]='h00000000;
    rd_cycle[ 9581] = 1'b0;  wr_cycle[ 9581] = 1'b1;  addr_rom[ 9581]='h00003394;  wr_data_rom[ 9581]='h0000258c;
    rd_cycle[ 9582] = 1'b0;  wr_cycle[ 9582] = 1'b1;  addr_rom[ 9582]='h00000710;  wr_data_rom[ 9582]='h0000345b;
    rd_cycle[ 9583] = 1'b1;  wr_cycle[ 9583] = 1'b0;  addr_rom[ 9583]='h000010f4;  wr_data_rom[ 9583]='h00000000;
    rd_cycle[ 9584] = 1'b0;  wr_cycle[ 9584] = 1'b1;  addr_rom[ 9584]='h00000488;  wr_data_rom[ 9584]='h000021b0;
    rd_cycle[ 9585] = 1'b0;  wr_cycle[ 9585] = 1'b1;  addr_rom[ 9585]='h00002fdc;  wr_data_rom[ 9585]='h00001df1;
    rd_cycle[ 9586] = 1'b1;  wr_cycle[ 9586] = 1'b0;  addr_rom[ 9586]='h00000430;  wr_data_rom[ 9586]='h00000000;
    rd_cycle[ 9587] = 1'b1;  wr_cycle[ 9587] = 1'b0;  addr_rom[ 9587]='h00001cf8;  wr_data_rom[ 9587]='h00000000;
    rd_cycle[ 9588] = 1'b1;  wr_cycle[ 9588] = 1'b0;  addr_rom[ 9588]='h000002d8;  wr_data_rom[ 9588]='h00000000;
    rd_cycle[ 9589] = 1'b0;  wr_cycle[ 9589] = 1'b1;  addr_rom[ 9589]='h00002194;  wr_data_rom[ 9589]='h00000713;
    rd_cycle[ 9590] = 1'b0;  wr_cycle[ 9590] = 1'b1;  addr_rom[ 9590]='h00001900;  wr_data_rom[ 9590]='h00000719;
    rd_cycle[ 9591] = 1'b0;  wr_cycle[ 9591] = 1'b1;  addr_rom[ 9591]='h000030f0;  wr_data_rom[ 9591]='h000013ea;
    rd_cycle[ 9592] = 1'b1;  wr_cycle[ 9592] = 1'b0;  addr_rom[ 9592]='h00001720;  wr_data_rom[ 9592]='h00000000;
    rd_cycle[ 9593] = 1'b0;  wr_cycle[ 9593] = 1'b1;  addr_rom[ 9593]='h00003400;  wr_data_rom[ 9593]='h00002195;
    rd_cycle[ 9594] = 1'b1;  wr_cycle[ 9594] = 1'b0;  addr_rom[ 9594]='h000034b0;  wr_data_rom[ 9594]='h00000000;
    rd_cycle[ 9595] = 1'b0;  wr_cycle[ 9595] = 1'b1;  addr_rom[ 9595]='h00003e8c;  wr_data_rom[ 9595]='h00003fb5;
    rd_cycle[ 9596] = 1'b1;  wr_cycle[ 9596] = 1'b0;  addr_rom[ 9596]='h00003a68;  wr_data_rom[ 9596]='h00000000;
    rd_cycle[ 9597] = 1'b1;  wr_cycle[ 9597] = 1'b0;  addr_rom[ 9597]='h00001b20;  wr_data_rom[ 9597]='h00000000;
    rd_cycle[ 9598] = 1'b1;  wr_cycle[ 9598] = 1'b0;  addr_rom[ 9598]='h00003228;  wr_data_rom[ 9598]='h00000000;
    rd_cycle[ 9599] = 1'b1;  wr_cycle[ 9599] = 1'b0;  addr_rom[ 9599]='h00001e44;  wr_data_rom[ 9599]='h00000000;
    rd_cycle[ 9600] = 1'b1;  wr_cycle[ 9600] = 1'b0;  addr_rom[ 9600]='h00001e1c;  wr_data_rom[ 9600]='h00000000;
    rd_cycle[ 9601] = 1'b1;  wr_cycle[ 9601] = 1'b0;  addr_rom[ 9601]='h00000b24;  wr_data_rom[ 9601]='h00000000;
    rd_cycle[ 9602] = 1'b1;  wr_cycle[ 9602] = 1'b0;  addr_rom[ 9602]='h00002600;  wr_data_rom[ 9602]='h00000000;
    rd_cycle[ 9603] = 1'b1;  wr_cycle[ 9603] = 1'b0;  addr_rom[ 9603]='h000018a4;  wr_data_rom[ 9603]='h00000000;
    rd_cycle[ 9604] = 1'b1;  wr_cycle[ 9604] = 1'b0;  addr_rom[ 9604]='h00003dd0;  wr_data_rom[ 9604]='h00000000;
    rd_cycle[ 9605] = 1'b1;  wr_cycle[ 9605] = 1'b0;  addr_rom[ 9605]='h00003c44;  wr_data_rom[ 9605]='h00000000;
    rd_cycle[ 9606] = 1'b1;  wr_cycle[ 9606] = 1'b0;  addr_rom[ 9606]='h00003fe4;  wr_data_rom[ 9606]='h00000000;
    rd_cycle[ 9607] = 1'b0;  wr_cycle[ 9607] = 1'b1;  addr_rom[ 9607]='h000022e4;  wr_data_rom[ 9607]='h00002495;
    rd_cycle[ 9608] = 1'b0;  wr_cycle[ 9608] = 1'b1;  addr_rom[ 9608]='h000022dc;  wr_data_rom[ 9608]='h00001a94;
    rd_cycle[ 9609] = 1'b0;  wr_cycle[ 9609] = 1'b1;  addr_rom[ 9609]='h00002abc;  wr_data_rom[ 9609]='h000015fd;
    rd_cycle[ 9610] = 1'b0;  wr_cycle[ 9610] = 1'b1;  addr_rom[ 9610]='h00000b90;  wr_data_rom[ 9610]='h0000383b;
    rd_cycle[ 9611] = 1'b1;  wr_cycle[ 9611] = 1'b0;  addr_rom[ 9611]='h00000c88;  wr_data_rom[ 9611]='h00000000;
    rd_cycle[ 9612] = 1'b0;  wr_cycle[ 9612] = 1'b1;  addr_rom[ 9612]='h00003a0c;  wr_data_rom[ 9612]='h00003e6e;
    rd_cycle[ 9613] = 1'b0;  wr_cycle[ 9613] = 1'b1;  addr_rom[ 9613]='h00001474;  wr_data_rom[ 9613]='h0000251d;
    rd_cycle[ 9614] = 1'b0;  wr_cycle[ 9614] = 1'b1;  addr_rom[ 9614]='h00002bb0;  wr_data_rom[ 9614]='h00000ae0;
    rd_cycle[ 9615] = 1'b1;  wr_cycle[ 9615] = 1'b0;  addr_rom[ 9615]='h00001394;  wr_data_rom[ 9615]='h00000000;
    rd_cycle[ 9616] = 1'b0;  wr_cycle[ 9616] = 1'b1;  addr_rom[ 9616]='h00000cec;  wr_data_rom[ 9616]='h00000acd;
    rd_cycle[ 9617] = 1'b0;  wr_cycle[ 9617] = 1'b1;  addr_rom[ 9617]='h000032cc;  wr_data_rom[ 9617]='h00001468;
    rd_cycle[ 9618] = 1'b1;  wr_cycle[ 9618] = 1'b0;  addr_rom[ 9618]='h00001f54;  wr_data_rom[ 9618]='h00000000;
    rd_cycle[ 9619] = 1'b0;  wr_cycle[ 9619] = 1'b1;  addr_rom[ 9619]='h000039bc;  wr_data_rom[ 9619]='h000010ab;
    rd_cycle[ 9620] = 1'b0;  wr_cycle[ 9620] = 1'b1;  addr_rom[ 9620]='h00001c64;  wr_data_rom[ 9620]='h00002180;
    rd_cycle[ 9621] = 1'b0;  wr_cycle[ 9621] = 1'b1;  addr_rom[ 9621]='h00002434;  wr_data_rom[ 9621]='h000034cc;
    rd_cycle[ 9622] = 1'b1;  wr_cycle[ 9622] = 1'b0;  addr_rom[ 9622]='h00001d58;  wr_data_rom[ 9622]='h00000000;
    rd_cycle[ 9623] = 1'b1;  wr_cycle[ 9623] = 1'b0;  addr_rom[ 9623]='h00002ca4;  wr_data_rom[ 9623]='h00000000;
    rd_cycle[ 9624] = 1'b1;  wr_cycle[ 9624] = 1'b0;  addr_rom[ 9624]='h00003e2c;  wr_data_rom[ 9624]='h00000000;
    rd_cycle[ 9625] = 1'b0;  wr_cycle[ 9625] = 1'b1;  addr_rom[ 9625]='h000020b4;  wr_data_rom[ 9625]='h00000233;
    rd_cycle[ 9626] = 1'b0;  wr_cycle[ 9626] = 1'b1;  addr_rom[ 9626]='h000029a0;  wr_data_rom[ 9626]='h000016bd;
    rd_cycle[ 9627] = 1'b0;  wr_cycle[ 9627] = 1'b1;  addr_rom[ 9627]='h000022f8;  wr_data_rom[ 9627]='h00000f54;
    rd_cycle[ 9628] = 1'b1;  wr_cycle[ 9628] = 1'b0;  addr_rom[ 9628]='h000024a0;  wr_data_rom[ 9628]='h00000000;
    rd_cycle[ 9629] = 1'b1;  wr_cycle[ 9629] = 1'b0;  addr_rom[ 9629]='h00003f58;  wr_data_rom[ 9629]='h00000000;
    rd_cycle[ 9630] = 1'b1;  wr_cycle[ 9630] = 1'b0;  addr_rom[ 9630]='h00002d58;  wr_data_rom[ 9630]='h00000000;
    rd_cycle[ 9631] = 1'b0;  wr_cycle[ 9631] = 1'b1;  addr_rom[ 9631]='h00001694;  wr_data_rom[ 9631]='h00000c8d;
    rd_cycle[ 9632] = 1'b1;  wr_cycle[ 9632] = 1'b0;  addr_rom[ 9632]='h00001a20;  wr_data_rom[ 9632]='h00000000;
    rd_cycle[ 9633] = 1'b0;  wr_cycle[ 9633] = 1'b1;  addr_rom[ 9633]='h0000123c;  wr_data_rom[ 9633]='h00000158;
    rd_cycle[ 9634] = 1'b1;  wr_cycle[ 9634] = 1'b0;  addr_rom[ 9634]='h00000e70;  wr_data_rom[ 9634]='h00000000;
    rd_cycle[ 9635] = 1'b1;  wr_cycle[ 9635] = 1'b0;  addr_rom[ 9635]='h00003b08;  wr_data_rom[ 9635]='h00000000;
    rd_cycle[ 9636] = 1'b1;  wr_cycle[ 9636] = 1'b0;  addr_rom[ 9636]='h00002720;  wr_data_rom[ 9636]='h00000000;
    rd_cycle[ 9637] = 1'b1;  wr_cycle[ 9637] = 1'b0;  addr_rom[ 9637]='h000032d4;  wr_data_rom[ 9637]='h00000000;
    rd_cycle[ 9638] = 1'b1;  wr_cycle[ 9638] = 1'b0;  addr_rom[ 9638]='h000016dc;  wr_data_rom[ 9638]='h00000000;
    rd_cycle[ 9639] = 1'b1;  wr_cycle[ 9639] = 1'b0;  addr_rom[ 9639]='h000030b4;  wr_data_rom[ 9639]='h00000000;
    rd_cycle[ 9640] = 1'b0;  wr_cycle[ 9640] = 1'b1;  addr_rom[ 9640]='h000015cc;  wr_data_rom[ 9640]='h0000003d;
    rd_cycle[ 9641] = 1'b1;  wr_cycle[ 9641] = 1'b0;  addr_rom[ 9641]='h00003a48;  wr_data_rom[ 9641]='h00000000;
    rd_cycle[ 9642] = 1'b0;  wr_cycle[ 9642] = 1'b1;  addr_rom[ 9642]='h00002b0c;  wr_data_rom[ 9642]='h00000501;
    rd_cycle[ 9643] = 1'b0;  wr_cycle[ 9643] = 1'b1;  addr_rom[ 9643]='h00003060;  wr_data_rom[ 9643]='h000009c4;
    rd_cycle[ 9644] = 1'b0;  wr_cycle[ 9644] = 1'b1;  addr_rom[ 9644]='h00003a2c;  wr_data_rom[ 9644]='h000014b9;
    rd_cycle[ 9645] = 1'b0;  wr_cycle[ 9645] = 1'b1;  addr_rom[ 9645]='h00003dd4;  wr_data_rom[ 9645]='h00003ac2;
    rd_cycle[ 9646] = 1'b0;  wr_cycle[ 9646] = 1'b1;  addr_rom[ 9646]='h00002aa8;  wr_data_rom[ 9646]='h00001b14;
    rd_cycle[ 9647] = 1'b1;  wr_cycle[ 9647] = 1'b0;  addr_rom[ 9647]='h000032ac;  wr_data_rom[ 9647]='h00000000;
    rd_cycle[ 9648] = 1'b0;  wr_cycle[ 9648] = 1'b1;  addr_rom[ 9648]='h00002234;  wr_data_rom[ 9648]='h00001372;
    rd_cycle[ 9649] = 1'b0;  wr_cycle[ 9649] = 1'b1;  addr_rom[ 9649]='h00003ae4;  wr_data_rom[ 9649]='h00001c38;
    rd_cycle[ 9650] = 1'b1;  wr_cycle[ 9650] = 1'b0;  addr_rom[ 9650]='h000003cc;  wr_data_rom[ 9650]='h00000000;
    rd_cycle[ 9651] = 1'b1;  wr_cycle[ 9651] = 1'b0;  addr_rom[ 9651]='h000029d8;  wr_data_rom[ 9651]='h00000000;
    rd_cycle[ 9652] = 1'b0;  wr_cycle[ 9652] = 1'b1;  addr_rom[ 9652]='h00001730;  wr_data_rom[ 9652]='h00001cd7;
    rd_cycle[ 9653] = 1'b1;  wr_cycle[ 9653] = 1'b0;  addr_rom[ 9653]='h00003208;  wr_data_rom[ 9653]='h00000000;
    rd_cycle[ 9654] = 1'b0;  wr_cycle[ 9654] = 1'b1;  addr_rom[ 9654]='h000038d8;  wr_data_rom[ 9654]='h00000601;
    rd_cycle[ 9655] = 1'b1;  wr_cycle[ 9655] = 1'b0;  addr_rom[ 9655]='h00000624;  wr_data_rom[ 9655]='h00000000;
    rd_cycle[ 9656] = 1'b0;  wr_cycle[ 9656] = 1'b1;  addr_rom[ 9656]='h000005f0;  wr_data_rom[ 9656]='h00001bc2;
    rd_cycle[ 9657] = 1'b0;  wr_cycle[ 9657] = 1'b1;  addr_rom[ 9657]='h00001508;  wr_data_rom[ 9657]='h00003c69;
    rd_cycle[ 9658] = 1'b1;  wr_cycle[ 9658] = 1'b0;  addr_rom[ 9658]='h000034d8;  wr_data_rom[ 9658]='h00000000;
    rd_cycle[ 9659] = 1'b1;  wr_cycle[ 9659] = 1'b0;  addr_rom[ 9659]='h000020c4;  wr_data_rom[ 9659]='h00000000;
    rd_cycle[ 9660] = 1'b0;  wr_cycle[ 9660] = 1'b1;  addr_rom[ 9660]='h00003b74;  wr_data_rom[ 9660]='h00001368;
    rd_cycle[ 9661] = 1'b0;  wr_cycle[ 9661] = 1'b1;  addr_rom[ 9661]='h000035ec;  wr_data_rom[ 9661]='h00002cb7;
    rd_cycle[ 9662] = 1'b1;  wr_cycle[ 9662] = 1'b0;  addr_rom[ 9662]='h00000bd4;  wr_data_rom[ 9662]='h00000000;
    rd_cycle[ 9663] = 1'b0;  wr_cycle[ 9663] = 1'b1;  addr_rom[ 9663]='h000027fc;  wr_data_rom[ 9663]='h00001c67;
    rd_cycle[ 9664] = 1'b0;  wr_cycle[ 9664] = 1'b1;  addr_rom[ 9664]='h00000578;  wr_data_rom[ 9664]='h00001622;
    rd_cycle[ 9665] = 1'b0;  wr_cycle[ 9665] = 1'b1;  addr_rom[ 9665]='h00000b74;  wr_data_rom[ 9665]='h00000e53;
    rd_cycle[ 9666] = 1'b1;  wr_cycle[ 9666] = 1'b0;  addr_rom[ 9666]='h00002e40;  wr_data_rom[ 9666]='h00000000;
    rd_cycle[ 9667] = 1'b1;  wr_cycle[ 9667] = 1'b0;  addr_rom[ 9667]='h00000130;  wr_data_rom[ 9667]='h00000000;
    rd_cycle[ 9668] = 1'b1;  wr_cycle[ 9668] = 1'b0;  addr_rom[ 9668]='h00003480;  wr_data_rom[ 9668]='h00000000;
    rd_cycle[ 9669] = 1'b0;  wr_cycle[ 9669] = 1'b1;  addr_rom[ 9669]='h000029e0;  wr_data_rom[ 9669]='h00001cff;
    rd_cycle[ 9670] = 1'b1;  wr_cycle[ 9670] = 1'b0;  addr_rom[ 9670]='h00002a18;  wr_data_rom[ 9670]='h00000000;
    rd_cycle[ 9671] = 1'b0;  wr_cycle[ 9671] = 1'b1;  addr_rom[ 9671]='h000035e4;  wr_data_rom[ 9671]='h0000118e;
    rd_cycle[ 9672] = 1'b1;  wr_cycle[ 9672] = 1'b0;  addr_rom[ 9672]='h00003f48;  wr_data_rom[ 9672]='h00000000;
    rd_cycle[ 9673] = 1'b0;  wr_cycle[ 9673] = 1'b1;  addr_rom[ 9673]='h00001ab0;  wr_data_rom[ 9673]='h00001cbf;
    rd_cycle[ 9674] = 1'b1;  wr_cycle[ 9674] = 1'b0;  addr_rom[ 9674]='h0000183c;  wr_data_rom[ 9674]='h00000000;
    rd_cycle[ 9675] = 1'b0;  wr_cycle[ 9675] = 1'b1;  addr_rom[ 9675]='h00003340;  wr_data_rom[ 9675]='h000001cd;
    rd_cycle[ 9676] = 1'b1;  wr_cycle[ 9676] = 1'b0;  addr_rom[ 9676]='h00000234;  wr_data_rom[ 9676]='h00000000;
    rd_cycle[ 9677] = 1'b0;  wr_cycle[ 9677] = 1'b1;  addr_rom[ 9677]='h00000db8;  wr_data_rom[ 9677]='h00001c82;
    rd_cycle[ 9678] = 1'b0;  wr_cycle[ 9678] = 1'b1;  addr_rom[ 9678]='h00000360;  wr_data_rom[ 9678]='h00001c4a;
    rd_cycle[ 9679] = 1'b1;  wr_cycle[ 9679] = 1'b0;  addr_rom[ 9679]='h00003e28;  wr_data_rom[ 9679]='h00000000;
    rd_cycle[ 9680] = 1'b0;  wr_cycle[ 9680] = 1'b1;  addr_rom[ 9680]='h00001e60;  wr_data_rom[ 9680]='h00001d6f;
    rd_cycle[ 9681] = 1'b0;  wr_cycle[ 9681] = 1'b1;  addr_rom[ 9681]='h00003050;  wr_data_rom[ 9681]='h000022bc;
    rd_cycle[ 9682] = 1'b1;  wr_cycle[ 9682] = 1'b0;  addr_rom[ 9682]='h000026b4;  wr_data_rom[ 9682]='h00000000;
    rd_cycle[ 9683] = 1'b0;  wr_cycle[ 9683] = 1'b1;  addr_rom[ 9683]='h00002cd8;  wr_data_rom[ 9683]='h000006a4;
    rd_cycle[ 9684] = 1'b0;  wr_cycle[ 9684] = 1'b1;  addr_rom[ 9684]='h00002694;  wr_data_rom[ 9684]='h00000928;
    rd_cycle[ 9685] = 1'b1;  wr_cycle[ 9685] = 1'b0;  addr_rom[ 9685]='h0000161c;  wr_data_rom[ 9685]='h00000000;
    rd_cycle[ 9686] = 1'b1;  wr_cycle[ 9686] = 1'b0;  addr_rom[ 9686]='h0000055c;  wr_data_rom[ 9686]='h00000000;
    rd_cycle[ 9687] = 1'b0;  wr_cycle[ 9687] = 1'b1;  addr_rom[ 9687]='h00000a4c;  wr_data_rom[ 9687]='h000026af;
    rd_cycle[ 9688] = 1'b1;  wr_cycle[ 9688] = 1'b0;  addr_rom[ 9688]='h00002594;  wr_data_rom[ 9688]='h00000000;
    rd_cycle[ 9689] = 1'b1;  wr_cycle[ 9689] = 1'b0;  addr_rom[ 9689]='h00002000;  wr_data_rom[ 9689]='h00000000;
    rd_cycle[ 9690] = 1'b1;  wr_cycle[ 9690] = 1'b0;  addr_rom[ 9690]='h000031fc;  wr_data_rom[ 9690]='h00000000;
    rd_cycle[ 9691] = 1'b1;  wr_cycle[ 9691] = 1'b0;  addr_rom[ 9691]='h00002aa8;  wr_data_rom[ 9691]='h00000000;
    rd_cycle[ 9692] = 1'b1;  wr_cycle[ 9692] = 1'b0;  addr_rom[ 9692]='h00000bb8;  wr_data_rom[ 9692]='h00000000;
    rd_cycle[ 9693] = 1'b0;  wr_cycle[ 9693] = 1'b1;  addr_rom[ 9693]='h00001208;  wr_data_rom[ 9693]='h00003585;
    rd_cycle[ 9694] = 1'b0;  wr_cycle[ 9694] = 1'b1;  addr_rom[ 9694]='h00003320;  wr_data_rom[ 9694]='h00001da2;
    rd_cycle[ 9695] = 1'b1;  wr_cycle[ 9695] = 1'b0;  addr_rom[ 9695]='h00000eb0;  wr_data_rom[ 9695]='h00000000;
    rd_cycle[ 9696] = 1'b1;  wr_cycle[ 9696] = 1'b0;  addr_rom[ 9696]='h00001e48;  wr_data_rom[ 9696]='h00000000;
    rd_cycle[ 9697] = 1'b0;  wr_cycle[ 9697] = 1'b1;  addr_rom[ 9697]='h00000100;  wr_data_rom[ 9697]='h00000ebf;
    rd_cycle[ 9698] = 1'b0;  wr_cycle[ 9698] = 1'b1;  addr_rom[ 9698]='h00003424;  wr_data_rom[ 9698]='h00000b7d;
    rd_cycle[ 9699] = 1'b0;  wr_cycle[ 9699] = 1'b1;  addr_rom[ 9699]='h0000254c;  wr_data_rom[ 9699]='h00000db0;
    rd_cycle[ 9700] = 1'b1;  wr_cycle[ 9700] = 1'b0;  addr_rom[ 9700]='h000013dc;  wr_data_rom[ 9700]='h00000000;
    rd_cycle[ 9701] = 1'b1;  wr_cycle[ 9701] = 1'b0;  addr_rom[ 9701]='h00003b40;  wr_data_rom[ 9701]='h00000000;
    rd_cycle[ 9702] = 1'b0;  wr_cycle[ 9702] = 1'b1;  addr_rom[ 9702]='h000017a4;  wr_data_rom[ 9702]='h00000d21;
    rd_cycle[ 9703] = 1'b0;  wr_cycle[ 9703] = 1'b1;  addr_rom[ 9703]='h000026b8;  wr_data_rom[ 9703]='h00003410;
    rd_cycle[ 9704] = 1'b0;  wr_cycle[ 9704] = 1'b1;  addr_rom[ 9704]='h00003cd0;  wr_data_rom[ 9704]='h00000625;
    rd_cycle[ 9705] = 1'b0;  wr_cycle[ 9705] = 1'b1;  addr_rom[ 9705]='h00003050;  wr_data_rom[ 9705]='h000020d8;
    rd_cycle[ 9706] = 1'b0;  wr_cycle[ 9706] = 1'b1;  addr_rom[ 9706]='h00002198;  wr_data_rom[ 9706]='h000019a0;
    rd_cycle[ 9707] = 1'b0;  wr_cycle[ 9707] = 1'b1;  addr_rom[ 9707]='h00002858;  wr_data_rom[ 9707]='h000009f1;
    rd_cycle[ 9708] = 1'b0;  wr_cycle[ 9708] = 1'b1;  addr_rom[ 9708]='h00001960;  wr_data_rom[ 9708]='h0000352d;
    rd_cycle[ 9709] = 1'b1;  wr_cycle[ 9709] = 1'b0;  addr_rom[ 9709]='h000012d8;  wr_data_rom[ 9709]='h00000000;
    rd_cycle[ 9710] = 1'b0;  wr_cycle[ 9710] = 1'b1;  addr_rom[ 9710]='h000026ec;  wr_data_rom[ 9710]='h00000990;
    rd_cycle[ 9711] = 1'b1;  wr_cycle[ 9711] = 1'b0;  addr_rom[ 9711]='h000017f0;  wr_data_rom[ 9711]='h00000000;
    rd_cycle[ 9712] = 1'b1;  wr_cycle[ 9712] = 1'b0;  addr_rom[ 9712]='h0000168c;  wr_data_rom[ 9712]='h00000000;
    rd_cycle[ 9713] = 1'b0;  wr_cycle[ 9713] = 1'b1;  addr_rom[ 9713]='h00002064;  wr_data_rom[ 9713]='h00003fa8;
    rd_cycle[ 9714] = 1'b0;  wr_cycle[ 9714] = 1'b1;  addr_rom[ 9714]='h000021e0;  wr_data_rom[ 9714]='h0000130c;
    rd_cycle[ 9715] = 1'b1;  wr_cycle[ 9715] = 1'b0;  addr_rom[ 9715]='h00002eb4;  wr_data_rom[ 9715]='h00000000;
    rd_cycle[ 9716] = 1'b1;  wr_cycle[ 9716] = 1'b0;  addr_rom[ 9716]='h000029d4;  wr_data_rom[ 9716]='h00000000;
    rd_cycle[ 9717] = 1'b0;  wr_cycle[ 9717] = 1'b1;  addr_rom[ 9717]='h000025a8;  wr_data_rom[ 9717]='h00000617;
    rd_cycle[ 9718] = 1'b0;  wr_cycle[ 9718] = 1'b1;  addr_rom[ 9718]='h00002048;  wr_data_rom[ 9718]='h00001c35;
    rd_cycle[ 9719] = 1'b0;  wr_cycle[ 9719] = 1'b1;  addr_rom[ 9719]='h000011dc;  wr_data_rom[ 9719]='h00000a00;
    rd_cycle[ 9720] = 1'b1;  wr_cycle[ 9720] = 1'b0;  addr_rom[ 9720]='h00003e78;  wr_data_rom[ 9720]='h00000000;
    rd_cycle[ 9721] = 1'b1;  wr_cycle[ 9721] = 1'b0;  addr_rom[ 9721]='h00003a0c;  wr_data_rom[ 9721]='h00000000;
    rd_cycle[ 9722] = 1'b0;  wr_cycle[ 9722] = 1'b1;  addr_rom[ 9722]='h00000030;  wr_data_rom[ 9722]='h00002a03;
    rd_cycle[ 9723] = 1'b0;  wr_cycle[ 9723] = 1'b1;  addr_rom[ 9723]='h00003b38;  wr_data_rom[ 9723]='h0000394f;
    rd_cycle[ 9724] = 1'b1;  wr_cycle[ 9724] = 1'b0;  addr_rom[ 9724]='h000013cc;  wr_data_rom[ 9724]='h00000000;
    rd_cycle[ 9725] = 1'b1;  wr_cycle[ 9725] = 1'b0;  addr_rom[ 9725]='h00002810;  wr_data_rom[ 9725]='h00000000;
    rd_cycle[ 9726] = 1'b0;  wr_cycle[ 9726] = 1'b1;  addr_rom[ 9726]='h000024dc;  wr_data_rom[ 9726]='h00000e04;
    rd_cycle[ 9727] = 1'b0;  wr_cycle[ 9727] = 1'b1;  addr_rom[ 9727]='h00002a38;  wr_data_rom[ 9727]='h0000209b;
    rd_cycle[ 9728] = 1'b1;  wr_cycle[ 9728] = 1'b0;  addr_rom[ 9728]='h000020c8;  wr_data_rom[ 9728]='h00000000;
    rd_cycle[ 9729] = 1'b1;  wr_cycle[ 9729] = 1'b0;  addr_rom[ 9729]='h0000067c;  wr_data_rom[ 9729]='h00000000;
    rd_cycle[ 9730] = 1'b1;  wr_cycle[ 9730] = 1'b0;  addr_rom[ 9730]='h000023a4;  wr_data_rom[ 9730]='h00000000;
    rd_cycle[ 9731] = 1'b0;  wr_cycle[ 9731] = 1'b1;  addr_rom[ 9731]='h00003d34;  wr_data_rom[ 9731]='h00001999;
    rd_cycle[ 9732] = 1'b1;  wr_cycle[ 9732] = 1'b0;  addr_rom[ 9732]='h00002bbc;  wr_data_rom[ 9732]='h00000000;
    rd_cycle[ 9733] = 1'b1;  wr_cycle[ 9733] = 1'b0;  addr_rom[ 9733]='h0000100c;  wr_data_rom[ 9733]='h00000000;
    rd_cycle[ 9734] = 1'b1;  wr_cycle[ 9734] = 1'b0;  addr_rom[ 9734]='h000025a0;  wr_data_rom[ 9734]='h00000000;
    rd_cycle[ 9735] = 1'b0;  wr_cycle[ 9735] = 1'b1;  addr_rom[ 9735]='h00003aac;  wr_data_rom[ 9735]='h00001b14;
    rd_cycle[ 9736] = 1'b1;  wr_cycle[ 9736] = 1'b0;  addr_rom[ 9736]='h00002e10;  wr_data_rom[ 9736]='h00000000;
    rd_cycle[ 9737] = 1'b1;  wr_cycle[ 9737] = 1'b0;  addr_rom[ 9737]='h000018fc;  wr_data_rom[ 9737]='h00000000;
    rd_cycle[ 9738] = 1'b0;  wr_cycle[ 9738] = 1'b1;  addr_rom[ 9738]='h00001068;  wr_data_rom[ 9738]='h00001366;
    rd_cycle[ 9739] = 1'b1;  wr_cycle[ 9739] = 1'b0;  addr_rom[ 9739]='h000027b0;  wr_data_rom[ 9739]='h00000000;
    rd_cycle[ 9740] = 1'b1;  wr_cycle[ 9740] = 1'b0;  addr_rom[ 9740]='h000021d4;  wr_data_rom[ 9740]='h00000000;
    rd_cycle[ 9741] = 1'b1;  wr_cycle[ 9741] = 1'b0;  addr_rom[ 9741]='h00001b50;  wr_data_rom[ 9741]='h00000000;
    rd_cycle[ 9742] = 1'b1;  wr_cycle[ 9742] = 1'b0;  addr_rom[ 9742]='h00000b64;  wr_data_rom[ 9742]='h00000000;
    rd_cycle[ 9743] = 1'b1;  wr_cycle[ 9743] = 1'b0;  addr_rom[ 9743]='h0000303c;  wr_data_rom[ 9743]='h00000000;
    rd_cycle[ 9744] = 1'b1;  wr_cycle[ 9744] = 1'b0;  addr_rom[ 9744]='h000013b8;  wr_data_rom[ 9744]='h00000000;
    rd_cycle[ 9745] = 1'b1;  wr_cycle[ 9745] = 1'b0;  addr_rom[ 9745]='h00001418;  wr_data_rom[ 9745]='h00000000;
    rd_cycle[ 9746] = 1'b0;  wr_cycle[ 9746] = 1'b1;  addr_rom[ 9746]='h00000efc;  wr_data_rom[ 9746]='h00003ba5;
    rd_cycle[ 9747] = 1'b1;  wr_cycle[ 9747] = 1'b0;  addr_rom[ 9747]='h00000eb4;  wr_data_rom[ 9747]='h00000000;
    rd_cycle[ 9748] = 1'b1;  wr_cycle[ 9748] = 1'b0;  addr_rom[ 9748]='h00000304;  wr_data_rom[ 9748]='h00000000;
    rd_cycle[ 9749] = 1'b1;  wr_cycle[ 9749] = 1'b0;  addr_rom[ 9749]='h00002c54;  wr_data_rom[ 9749]='h00000000;
    rd_cycle[ 9750] = 1'b0;  wr_cycle[ 9750] = 1'b1;  addr_rom[ 9750]='h00002d84;  wr_data_rom[ 9750]='h00002884;
    rd_cycle[ 9751] = 1'b1;  wr_cycle[ 9751] = 1'b0;  addr_rom[ 9751]='h00003f5c;  wr_data_rom[ 9751]='h00000000;
    rd_cycle[ 9752] = 1'b1;  wr_cycle[ 9752] = 1'b0;  addr_rom[ 9752]='h00002178;  wr_data_rom[ 9752]='h00000000;
    rd_cycle[ 9753] = 1'b1;  wr_cycle[ 9753] = 1'b0;  addr_rom[ 9753]='h000009e4;  wr_data_rom[ 9753]='h00000000;
    rd_cycle[ 9754] = 1'b1;  wr_cycle[ 9754] = 1'b0;  addr_rom[ 9754]='h00001a28;  wr_data_rom[ 9754]='h00000000;
    rd_cycle[ 9755] = 1'b1;  wr_cycle[ 9755] = 1'b0;  addr_rom[ 9755]='h000002b4;  wr_data_rom[ 9755]='h00000000;
    rd_cycle[ 9756] = 1'b0;  wr_cycle[ 9756] = 1'b1;  addr_rom[ 9756]='h00002f88;  wr_data_rom[ 9756]='h00003716;
    rd_cycle[ 9757] = 1'b1;  wr_cycle[ 9757] = 1'b0;  addr_rom[ 9757]='h00003b6c;  wr_data_rom[ 9757]='h00000000;
    rd_cycle[ 9758] = 1'b0;  wr_cycle[ 9758] = 1'b1;  addr_rom[ 9758]='h00002808;  wr_data_rom[ 9758]='h00002fa1;
    rd_cycle[ 9759] = 1'b1;  wr_cycle[ 9759] = 1'b0;  addr_rom[ 9759]='h00001138;  wr_data_rom[ 9759]='h00000000;
    rd_cycle[ 9760] = 1'b1;  wr_cycle[ 9760] = 1'b0;  addr_rom[ 9760]='h00000854;  wr_data_rom[ 9760]='h00000000;
    rd_cycle[ 9761] = 1'b0;  wr_cycle[ 9761] = 1'b1;  addr_rom[ 9761]='h0000273c;  wr_data_rom[ 9761]='h000021ca;
    rd_cycle[ 9762] = 1'b0;  wr_cycle[ 9762] = 1'b1;  addr_rom[ 9762]='h00002774;  wr_data_rom[ 9762]='h00001ac5;
    rd_cycle[ 9763] = 1'b1;  wr_cycle[ 9763] = 1'b0;  addr_rom[ 9763]='h00002130;  wr_data_rom[ 9763]='h00000000;
    rd_cycle[ 9764] = 1'b1;  wr_cycle[ 9764] = 1'b0;  addr_rom[ 9764]='h00003a1c;  wr_data_rom[ 9764]='h00000000;
    rd_cycle[ 9765] = 1'b1;  wr_cycle[ 9765] = 1'b0;  addr_rom[ 9765]='h00002fac;  wr_data_rom[ 9765]='h00000000;
    rd_cycle[ 9766] = 1'b1;  wr_cycle[ 9766] = 1'b0;  addr_rom[ 9766]='h000019b4;  wr_data_rom[ 9766]='h00000000;
    rd_cycle[ 9767] = 1'b1;  wr_cycle[ 9767] = 1'b0;  addr_rom[ 9767]='h000038e8;  wr_data_rom[ 9767]='h00000000;
    rd_cycle[ 9768] = 1'b1;  wr_cycle[ 9768] = 1'b0;  addr_rom[ 9768]='h00002878;  wr_data_rom[ 9768]='h00000000;
    rd_cycle[ 9769] = 1'b0;  wr_cycle[ 9769] = 1'b1;  addr_rom[ 9769]='h00001418;  wr_data_rom[ 9769]='h00003ff5;
    rd_cycle[ 9770] = 1'b0;  wr_cycle[ 9770] = 1'b1;  addr_rom[ 9770]='h000031f4;  wr_data_rom[ 9770]='h00003f81;
    rd_cycle[ 9771] = 1'b1;  wr_cycle[ 9771] = 1'b0;  addr_rom[ 9771]='h00002c38;  wr_data_rom[ 9771]='h00000000;
    rd_cycle[ 9772] = 1'b0;  wr_cycle[ 9772] = 1'b1;  addr_rom[ 9772]='h00003664;  wr_data_rom[ 9772]='h00002a3f;
    rd_cycle[ 9773] = 1'b0;  wr_cycle[ 9773] = 1'b1;  addr_rom[ 9773]='h000030dc;  wr_data_rom[ 9773]='h00000eed;
    rd_cycle[ 9774] = 1'b0;  wr_cycle[ 9774] = 1'b1;  addr_rom[ 9774]='h00000704;  wr_data_rom[ 9774]='h00003ef8;
    rd_cycle[ 9775] = 1'b0;  wr_cycle[ 9775] = 1'b1;  addr_rom[ 9775]='h00002098;  wr_data_rom[ 9775]='h00001677;
    rd_cycle[ 9776] = 1'b0;  wr_cycle[ 9776] = 1'b1;  addr_rom[ 9776]='h000030b4;  wr_data_rom[ 9776]='h0000107c;
    rd_cycle[ 9777] = 1'b1;  wr_cycle[ 9777] = 1'b0;  addr_rom[ 9777]='h000014dc;  wr_data_rom[ 9777]='h00000000;
    rd_cycle[ 9778] = 1'b0;  wr_cycle[ 9778] = 1'b1;  addr_rom[ 9778]='h000001e8;  wr_data_rom[ 9778]='h00001c50;
    rd_cycle[ 9779] = 1'b1;  wr_cycle[ 9779] = 1'b0;  addr_rom[ 9779]='h00003728;  wr_data_rom[ 9779]='h00000000;
    rd_cycle[ 9780] = 1'b0;  wr_cycle[ 9780] = 1'b1;  addr_rom[ 9780]='h00000e4c;  wr_data_rom[ 9780]='h00003f38;
    rd_cycle[ 9781] = 1'b0;  wr_cycle[ 9781] = 1'b1;  addr_rom[ 9781]='h00003b1c;  wr_data_rom[ 9781]='h00001244;
    rd_cycle[ 9782] = 1'b0;  wr_cycle[ 9782] = 1'b1;  addr_rom[ 9782]='h00002c38;  wr_data_rom[ 9782]='h00000a6a;
    rd_cycle[ 9783] = 1'b0;  wr_cycle[ 9783] = 1'b1;  addr_rom[ 9783]='h00003ee4;  wr_data_rom[ 9783]='h00001531;
    rd_cycle[ 9784] = 1'b0;  wr_cycle[ 9784] = 1'b1;  addr_rom[ 9784]='h00000254;  wr_data_rom[ 9784]='h00003af6;
    rd_cycle[ 9785] = 1'b1;  wr_cycle[ 9785] = 1'b0;  addr_rom[ 9785]='h00002700;  wr_data_rom[ 9785]='h00000000;
    rd_cycle[ 9786] = 1'b1;  wr_cycle[ 9786] = 1'b0;  addr_rom[ 9786]='h00003e4c;  wr_data_rom[ 9786]='h00000000;
    rd_cycle[ 9787] = 1'b1;  wr_cycle[ 9787] = 1'b0;  addr_rom[ 9787]='h000010d0;  wr_data_rom[ 9787]='h00000000;
    rd_cycle[ 9788] = 1'b0;  wr_cycle[ 9788] = 1'b1;  addr_rom[ 9788]='h00003e48;  wr_data_rom[ 9788]='h00003a9c;
    rd_cycle[ 9789] = 1'b0;  wr_cycle[ 9789] = 1'b1;  addr_rom[ 9789]='h00002328;  wr_data_rom[ 9789]='h000028f3;
    rd_cycle[ 9790] = 1'b0;  wr_cycle[ 9790] = 1'b1;  addr_rom[ 9790]='h00000f6c;  wr_data_rom[ 9790]='h00001c18;
    rd_cycle[ 9791] = 1'b0;  wr_cycle[ 9791] = 1'b1;  addr_rom[ 9791]='h000035b8;  wr_data_rom[ 9791]='h00003c26;
    rd_cycle[ 9792] = 1'b1;  wr_cycle[ 9792] = 1'b0;  addr_rom[ 9792]='h000027d4;  wr_data_rom[ 9792]='h00000000;
    rd_cycle[ 9793] = 1'b0;  wr_cycle[ 9793] = 1'b1;  addr_rom[ 9793]='h000038ac;  wr_data_rom[ 9793]='h00000799;
    rd_cycle[ 9794] = 1'b1;  wr_cycle[ 9794] = 1'b0;  addr_rom[ 9794]='h00002280;  wr_data_rom[ 9794]='h00000000;
    rd_cycle[ 9795] = 1'b1;  wr_cycle[ 9795] = 1'b0;  addr_rom[ 9795]='h00001318;  wr_data_rom[ 9795]='h00000000;
    rd_cycle[ 9796] = 1'b0;  wr_cycle[ 9796] = 1'b1;  addr_rom[ 9796]='h00002a48;  wr_data_rom[ 9796]='h000000ff;
    rd_cycle[ 9797] = 1'b0;  wr_cycle[ 9797] = 1'b1;  addr_rom[ 9797]='h00002038;  wr_data_rom[ 9797]='h000002c1;
    rd_cycle[ 9798] = 1'b1;  wr_cycle[ 9798] = 1'b0;  addr_rom[ 9798]='h00000e24;  wr_data_rom[ 9798]='h00000000;
    rd_cycle[ 9799] = 1'b1;  wr_cycle[ 9799] = 1'b0;  addr_rom[ 9799]='h00002d48;  wr_data_rom[ 9799]='h00000000;
    rd_cycle[ 9800] = 1'b0;  wr_cycle[ 9800] = 1'b1;  addr_rom[ 9800]='h00003a30;  wr_data_rom[ 9800]='h00003283;
    rd_cycle[ 9801] = 1'b0;  wr_cycle[ 9801] = 1'b1;  addr_rom[ 9801]='h00001df4;  wr_data_rom[ 9801]='h000022e5;
    rd_cycle[ 9802] = 1'b1;  wr_cycle[ 9802] = 1'b0;  addr_rom[ 9802]='h00002b04;  wr_data_rom[ 9802]='h00000000;
    rd_cycle[ 9803] = 1'b0;  wr_cycle[ 9803] = 1'b1;  addr_rom[ 9803]='h000026b4;  wr_data_rom[ 9803]='h00003fa2;
    rd_cycle[ 9804] = 1'b0;  wr_cycle[ 9804] = 1'b1;  addr_rom[ 9804]='h00002258;  wr_data_rom[ 9804]='h000012be;
    rd_cycle[ 9805] = 1'b0;  wr_cycle[ 9805] = 1'b1;  addr_rom[ 9805]='h00003754;  wr_data_rom[ 9805]='h00001136;
    rd_cycle[ 9806] = 1'b1;  wr_cycle[ 9806] = 1'b0;  addr_rom[ 9806]='h00000ed8;  wr_data_rom[ 9806]='h00000000;
    rd_cycle[ 9807] = 1'b1;  wr_cycle[ 9807] = 1'b0;  addr_rom[ 9807]='h000003bc;  wr_data_rom[ 9807]='h00000000;
    rd_cycle[ 9808] = 1'b1;  wr_cycle[ 9808] = 1'b0;  addr_rom[ 9808]='h0000278c;  wr_data_rom[ 9808]='h00000000;
    rd_cycle[ 9809] = 1'b0;  wr_cycle[ 9809] = 1'b1;  addr_rom[ 9809]='h00000990;  wr_data_rom[ 9809]='h0000383d;
    rd_cycle[ 9810] = 1'b0;  wr_cycle[ 9810] = 1'b1;  addr_rom[ 9810]='h00002aa4;  wr_data_rom[ 9810]='h000039a4;
    rd_cycle[ 9811] = 1'b1;  wr_cycle[ 9811] = 1'b0;  addr_rom[ 9811]='h00001d94;  wr_data_rom[ 9811]='h00000000;
    rd_cycle[ 9812] = 1'b1;  wr_cycle[ 9812] = 1'b0;  addr_rom[ 9812]='h000014b4;  wr_data_rom[ 9812]='h00000000;
    rd_cycle[ 9813] = 1'b0;  wr_cycle[ 9813] = 1'b1;  addr_rom[ 9813]='h0000348c;  wr_data_rom[ 9813]='h000037be;
    rd_cycle[ 9814] = 1'b0;  wr_cycle[ 9814] = 1'b1;  addr_rom[ 9814]='h00002d68;  wr_data_rom[ 9814]='h0000021e;
    rd_cycle[ 9815] = 1'b1;  wr_cycle[ 9815] = 1'b0;  addr_rom[ 9815]='h00000dac;  wr_data_rom[ 9815]='h00000000;
    rd_cycle[ 9816] = 1'b1;  wr_cycle[ 9816] = 1'b0;  addr_rom[ 9816]='h00001894;  wr_data_rom[ 9816]='h00000000;
    rd_cycle[ 9817] = 1'b1;  wr_cycle[ 9817] = 1'b0;  addr_rom[ 9817]='h00002fd8;  wr_data_rom[ 9817]='h00000000;
    rd_cycle[ 9818] = 1'b1;  wr_cycle[ 9818] = 1'b0;  addr_rom[ 9818]='h0000076c;  wr_data_rom[ 9818]='h00000000;
    rd_cycle[ 9819] = 1'b0;  wr_cycle[ 9819] = 1'b1;  addr_rom[ 9819]='h00003574;  wr_data_rom[ 9819]='h00001c1a;
    rd_cycle[ 9820] = 1'b1;  wr_cycle[ 9820] = 1'b0;  addr_rom[ 9820]='h000022ac;  wr_data_rom[ 9820]='h00000000;
    rd_cycle[ 9821] = 1'b0;  wr_cycle[ 9821] = 1'b1;  addr_rom[ 9821]='h0000073c;  wr_data_rom[ 9821]='h00001888;
    rd_cycle[ 9822] = 1'b1;  wr_cycle[ 9822] = 1'b0;  addr_rom[ 9822]='h00001080;  wr_data_rom[ 9822]='h00000000;
    rd_cycle[ 9823] = 1'b0;  wr_cycle[ 9823] = 1'b1;  addr_rom[ 9823]='h00002098;  wr_data_rom[ 9823]='h000008a5;
    rd_cycle[ 9824] = 1'b0;  wr_cycle[ 9824] = 1'b1;  addr_rom[ 9824]='h000024c8;  wr_data_rom[ 9824]='h00003f6c;
    rd_cycle[ 9825] = 1'b1;  wr_cycle[ 9825] = 1'b0;  addr_rom[ 9825]='h000039c0;  wr_data_rom[ 9825]='h00000000;
    rd_cycle[ 9826] = 1'b1;  wr_cycle[ 9826] = 1'b0;  addr_rom[ 9826]='h000032d8;  wr_data_rom[ 9826]='h00000000;
    rd_cycle[ 9827] = 1'b1;  wr_cycle[ 9827] = 1'b0;  addr_rom[ 9827]='h00002e44;  wr_data_rom[ 9827]='h00000000;
    rd_cycle[ 9828] = 1'b1;  wr_cycle[ 9828] = 1'b0;  addr_rom[ 9828]='h00003620;  wr_data_rom[ 9828]='h00000000;
    rd_cycle[ 9829] = 1'b1;  wr_cycle[ 9829] = 1'b0;  addr_rom[ 9829]='h00001e48;  wr_data_rom[ 9829]='h00000000;
    rd_cycle[ 9830] = 1'b1;  wr_cycle[ 9830] = 1'b0;  addr_rom[ 9830]='h00003b70;  wr_data_rom[ 9830]='h00000000;
    rd_cycle[ 9831] = 1'b1;  wr_cycle[ 9831] = 1'b0;  addr_rom[ 9831]='h00000e7c;  wr_data_rom[ 9831]='h00000000;
    rd_cycle[ 9832] = 1'b1;  wr_cycle[ 9832] = 1'b0;  addr_rom[ 9832]='h0000235c;  wr_data_rom[ 9832]='h00000000;
    rd_cycle[ 9833] = 1'b0;  wr_cycle[ 9833] = 1'b1;  addr_rom[ 9833]='h00001884;  wr_data_rom[ 9833]='h00003fef;
    rd_cycle[ 9834] = 1'b1;  wr_cycle[ 9834] = 1'b0;  addr_rom[ 9834]='h00003ed8;  wr_data_rom[ 9834]='h00000000;
    rd_cycle[ 9835] = 1'b1;  wr_cycle[ 9835] = 1'b0;  addr_rom[ 9835]='h0000072c;  wr_data_rom[ 9835]='h00000000;
    rd_cycle[ 9836] = 1'b1;  wr_cycle[ 9836] = 1'b0;  addr_rom[ 9836]='h000033b0;  wr_data_rom[ 9836]='h00000000;
    rd_cycle[ 9837] = 1'b0;  wr_cycle[ 9837] = 1'b1;  addr_rom[ 9837]='h00001360;  wr_data_rom[ 9837]='h000038ab;
    rd_cycle[ 9838] = 1'b1;  wr_cycle[ 9838] = 1'b0;  addr_rom[ 9838]='h00001aa8;  wr_data_rom[ 9838]='h00000000;
    rd_cycle[ 9839] = 1'b1;  wr_cycle[ 9839] = 1'b0;  addr_rom[ 9839]='h00000868;  wr_data_rom[ 9839]='h00000000;
    rd_cycle[ 9840] = 1'b0;  wr_cycle[ 9840] = 1'b1;  addr_rom[ 9840]='h000014e4;  wr_data_rom[ 9840]='h000006bc;
    rd_cycle[ 9841] = 1'b1;  wr_cycle[ 9841] = 1'b0;  addr_rom[ 9841]='h0000018c;  wr_data_rom[ 9841]='h00000000;
    rd_cycle[ 9842] = 1'b1;  wr_cycle[ 9842] = 1'b0;  addr_rom[ 9842]='h00002a40;  wr_data_rom[ 9842]='h00000000;
    rd_cycle[ 9843] = 1'b0;  wr_cycle[ 9843] = 1'b1;  addr_rom[ 9843]='h00003d2c;  wr_data_rom[ 9843]='h000016c8;
    rd_cycle[ 9844] = 1'b1;  wr_cycle[ 9844] = 1'b0;  addr_rom[ 9844]='h000001c4;  wr_data_rom[ 9844]='h00000000;
    rd_cycle[ 9845] = 1'b1;  wr_cycle[ 9845] = 1'b0;  addr_rom[ 9845]='h00000a48;  wr_data_rom[ 9845]='h00000000;
    rd_cycle[ 9846] = 1'b0;  wr_cycle[ 9846] = 1'b1;  addr_rom[ 9846]='h000001a8;  wr_data_rom[ 9846]='h000030b2;
    rd_cycle[ 9847] = 1'b1;  wr_cycle[ 9847] = 1'b0;  addr_rom[ 9847]='h000017dc;  wr_data_rom[ 9847]='h00000000;
    rd_cycle[ 9848] = 1'b1;  wr_cycle[ 9848] = 1'b0;  addr_rom[ 9848]='h000010dc;  wr_data_rom[ 9848]='h00000000;
    rd_cycle[ 9849] = 1'b0;  wr_cycle[ 9849] = 1'b1;  addr_rom[ 9849]='h00002720;  wr_data_rom[ 9849]='h0000382a;
    rd_cycle[ 9850] = 1'b1;  wr_cycle[ 9850] = 1'b0;  addr_rom[ 9850]='h00001d14;  wr_data_rom[ 9850]='h00000000;
    rd_cycle[ 9851] = 1'b1;  wr_cycle[ 9851] = 1'b0;  addr_rom[ 9851]='h000036a0;  wr_data_rom[ 9851]='h00000000;
    rd_cycle[ 9852] = 1'b1;  wr_cycle[ 9852] = 1'b0;  addr_rom[ 9852]='h00003b18;  wr_data_rom[ 9852]='h00000000;
    rd_cycle[ 9853] = 1'b1;  wr_cycle[ 9853] = 1'b0;  addr_rom[ 9853]='h00003108;  wr_data_rom[ 9853]='h00000000;
    rd_cycle[ 9854] = 1'b1;  wr_cycle[ 9854] = 1'b0;  addr_rom[ 9854]='h00003c80;  wr_data_rom[ 9854]='h00000000;
    rd_cycle[ 9855] = 1'b1;  wr_cycle[ 9855] = 1'b0;  addr_rom[ 9855]='h000010a0;  wr_data_rom[ 9855]='h00000000;
    rd_cycle[ 9856] = 1'b1;  wr_cycle[ 9856] = 1'b0;  addr_rom[ 9856]='h00003f18;  wr_data_rom[ 9856]='h00000000;
    rd_cycle[ 9857] = 1'b1;  wr_cycle[ 9857] = 1'b0;  addr_rom[ 9857]='h00001a4c;  wr_data_rom[ 9857]='h00000000;
    rd_cycle[ 9858] = 1'b1;  wr_cycle[ 9858] = 1'b0;  addr_rom[ 9858]='h00002788;  wr_data_rom[ 9858]='h00000000;
    rd_cycle[ 9859] = 1'b1;  wr_cycle[ 9859] = 1'b0;  addr_rom[ 9859]='h00000070;  wr_data_rom[ 9859]='h00000000;
    rd_cycle[ 9860] = 1'b0;  wr_cycle[ 9860] = 1'b1;  addr_rom[ 9860]='h00001268;  wr_data_rom[ 9860]='h00000cdf;
    rd_cycle[ 9861] = 1'b0;  wr_cycle[ 9861] = 1'b1;  addr_rom[ 9861]='h00003628;  wr_data_rom[ 9861]='h00003941;
    rd_cycle[ 9862] = 1'b0;  wr_cycle[ 9862] = 1'b1;  addr_rom[ 9862]='h00000f18;  wr_data_rom[ 9862]='h00001958;
    rd_cycle[ 9863] = 1'b1;  wr_cycle[ 9863] = 1'b0;  addr_rom[ 9863]='h00001874;  wr_data_rom[ 9863]='h00000000;
    rd_cycle[ 9864] = 1'b1;  wr_cycle[ 9864] = 1'b0;  addr_rom[ 9864]='h00003c28;  wr_data_rom[ 9864]='h00000000;
    rd_cycle[ 9865] = 1'b0;  wr_cycle[ 9865] = 1'b1;  addr_rom[ 9865]='h00001cd0;  wr_data_rom[ 9865]='h00001638;
    rd_cycle[ 9866] = 1'b1;  wr_cycle[ 9866] = 1'b0;  addr_rom[ 9866]='h000034f4;  wr_data_rom[ 9866]='h00000000;
    rd_cycle[ 9867] = 1'b1;  wr_cycle[ 9867] = 1'b0;  addr_rom[ 9867]='h00002bc8;  wr_data_rom[ 9867]='h00000000;
    rd_cycle[ 9868] = 1'b1;  wr_cycle[ 9868] = 1'b0;  addr_rom[ 9868]='h00002f58;  wr_data_rom[ 9868]='h00000000;
    rd_cycle[ 9869] = 1'b0;  wr_cycle[ 9869] = 1'b1;  addr_rom[ 9869]='h0000056c;  wr_data_rom[ 9869]='h00002ec7;
    rd_cycle[ 9870] = 1'b1;  wr_cycle[ 9870] = 1'b0;  addr_rom[ 9870]='h00002a34;  wr_data_rom[ 9870]='h00000000;
    rd_cycle[ 9871] = 1'b0;  wr_cycle[ 9871] = 1'b1;  addr_rom[ 9871]='h00001108;  wr_data_rom[ 9871]='h000025ea;
    rd_cycle[ 9872] = 1'b0;  wr_cycle[ 9872] = 1'b1;  addr_rom[ 9872]='h0000309c;  wr_data_rom[ 9872]='h000007cf;
    rd_cycle[ 9873] = 1'b1;  wr_cycle[ 9873] = 1'b0;  addr_rom[ 9873]='h000017f8;  wr_data_rom[ 9873]='h00000000;
    rd_cycle[ 9874] = 1'b0;  wr_cycle[ 9874] = 1'b1;  addr_rom[ 9874]='h00002590;  wr_data_rom[ 9874]='h00001b32;
    rd_cycle[ 9875] = 1'b0;  wr_cycle[ 9875] = 1'b1;  addr_rom[ 9875]='h00003c88;  wr_data_rom[ 9875]='h000037ad;
    rd_cycle[ 9876] = 1'b0;  wr_cycle[ 9876] = 1'b1;  addr_rom[ 9876]='h000015c4;  wr_data_rom[ 9876]='h000036d6;
    rd_cycle[ 9877] = 1'b0;  wr_cycle[ 9877] = 1'b1;  addr_rom[ 9877]='h00001368;  wr_data_rom[ 9877]='h00003c66;
    rd_cycle[ 9878] = 1'b1;  wr_cycle[ 9878] = 1'b0;  addr_rom[ 9878]='h000038b8;  wr_data_rom[ 9878]='h00000000;
    rd_cycle[ 9879] = 1'b1;  wr_cycle[ 9879] = 1'b0;  addr_rom[ 9879]='h00002040;  wr_data_rom[ 9879]='h00000000;
    rd_cycle[ 9880] = 1'b1;  wr_cycle[ 9880] = 1'b0;  addr_rom[ 9880]='h000014f0;  wr_data_rom[ 9880]='h00000000;
    rd_cycle[ 9881] = 1'b1;  wr_cycle[ 9881] = 1'b0;  addr_rom[ 9881]='h00001524;  wr_data_rom[ 9881]='h00000000;
    rd_cycle[ 9882] = 1'b1;  wr_cycle[ 9882] = 1'b0;  addr_rom[ 9882]='h00002ac8;  wr_data_rom[ 9882]='h00000000;
    rd_cycle[ 9883] = 1'b0;  wr_cycle[ 9883] = 1'b1;  addr_rom[ 9883]='h00001bdc;  wr_data_rom[ 9883]='h000002ec;
    rd_cycle[ 9884] = 1'b0;  wr_cycle[ 9884] = 1'b1;  addr_rom[ 9884]='h00002c9c;  wr_data_rom[ 9884]='h00001d20;
    rd_cycle[ 9885] = 1'b0;  wr_cycle[ 9885] = 1'b1;  addr_rom[ 9885]='h00003570;  wr_data_rom[ 9885]='h00001622;
    rd_cycle[ 9886] = 1'b0;  wr_cycle[ 9886] = 1'b1;  addr_rom[ 9886]='h00003630;  wr_data_rom[ 9886]='h00000a48;
    rd_cycle[ 9887] = 1'b0;  wr_cycle[ 9887] = 1'b1;  addr_rom[ 9887]='h00001f54;  wr_data_rom[ 9887]='h00002d1d;
    rd_cycle[ 9888] = 1'b1;  wr_cycle[ 9888] = 1'b0;  addr_rom[ 9888]='h000020bc;  wr_data_rom[ 9888]='h00000000;
    rd_cycle[ 9889] = 1'b0;  wr_cycle[ 9889] = 1'b1;  addr_rom[ 9889]='h00002028;  wr_data_rom[ 9889]='h0000202c;
    rd_cycle[ 9890] = 1'b1;  wr_cycle[ 9890] = 1'b0;  addr_rom[ 9890]='h00002cec;  wr_data_rom[ 9890]='h00000000;
    rd_cycle[ 9891] = 1'b0;  wr_cycle[ 9891] = 1'b1;  addr_rom[ 9891]='h000031c0;  wr_data_rom[ 9891]='h00003c8e;
    rd_cycle[ 9892] = 1'b1;  wr_cycle[ 9892] = 1'b0;  addr_rom[ 9892]='h000021a4;  wr_data_rom[ 9892]='h00000000;
    rd_cycle[ 9893] = 1'b1;  wr_cycle[ 9893] = 1'b0;  addr_rom[ 9893]='h00001a98;  wr_data_rom[ 9893]='h00000000;
    rd_cycle[ 9894] = 1'b0;  wr_cycle[ 9894] = 1'b1;  addr_rom[ 9894]='h00000874;  wr_data_rom[ 9894]='h0000237a;
    rd_cycle[ 9895] = 1'b1;  wr_cycle[ 9895] = 1'b0;  addr_rom[ 9895]='h00001de0;  wr_data_rom[ 9895]='h00000000;
    rd_cycle[ 9896] = 1'b1;  wr_cycle[ 9896] = 1'b0;  addr_rom[ 9896]='h000029b8;  wr_data_rom[ 9896]='h00000000;
    rd_cycle[ 9897] = 1'b0;  wr_cycle[ 9897] = 1'b1;  addr_rom[ 9897]='h00001884;  wr_data_rom[ 9897]='h000022d9;
    rd_cycle[ 9898] = 1'b0;  wr_cycle[ 9898] = 1'b1;  addr_rom[ 9898]='h00003b6c;  wr_data_rom[ 9898]='h00003302;
    rd_cycle[ 9899] = 1'b1;  wr_cycle[ 9899] = 1'b0;  addr_rom[ 9899]='h00000620;  wr_data_rom[ 9899]='h00000000;
    rd_cycle[ 9900] = 1'b0;  wr_cycle[ 9900] = 1'b1;  addr_rom[ 9900]='h0000218c;  wr_data_rom[ 9900]='h0000275f;
    rd_cycle[ 9901] = 1'b1;  wr_cycle[ 9901] = 1'b0;  addr_rom[ 9901]='h00002e64;  wr_data_rom[ 9901]='h00000000;
    rd_cycle[ 9902] = 1'b0;  wr_cycle[ 9902] = 1'b1;  addr_rom[ 9902]='h000021ec;  wr_data_rom[ 9902]='h00000cec;
    rd_cycle[ 9903] = 1'b1;  wr_cycle[ 9903] = 1'b0;  addr_rom[ 9903]='h0000306c;  wr_data_rom[ 9903]='h00000000;
    rd_cycle[ 9904] = 1'b1;  wr_cycle[ 9904] = 1'b0;  addr_rom[ 9904]='h000029d0;  wr_data_rom[ 9904]='h00000000;
    rd_cycle[ 9905] = 1'b0;  wr_cycle[ 9905] = 1'b1;  addr_rom[ 9905]='h00002444;  wr_data_rom[ 9905]='h0000144a;
    rd_cycle[ 9906] = 1'b1;  wr_cycle[ 9906] = 1'b0;  addr_rom[ 9906]='h00000a44;  wr_data_rom[ 9906]='h00000000;
    rd_cycle[ 9907] = 1'b0;  wr_cycle[ 9907] = 1'b1;  addr_rom[ 9907]='h00002e4c;  wr_data_rom[ 9907]='h00001c8e;
    rd_cycle[ 9908] = 1'b1;  wr_cycle[ 9908] = 1'b0;  addr_rom[ 9908]='h00002420;  wr_data_rom[ 9908]='h00000000;
    rd_cycle[ 9909] = 1'b0;  wr_cycle[ 9909] = 1'b1;  addr_rom[ 9909]='h000021b8;  wr_data_rom[ 9909]='h00003d3a;
    rd_cycle[ 9910] = 1'b1;  wr_cycle[ 9910] = 1'b0;  addr_rom[ 9910]='h00000bcc;  wr_data_rom[ 9910]='h00000000;
    rd_cycle[ 9911] = 1'b1;  wr_cycle[ 9911] = 1'b0;  addr_rom[ 9911]='h00000234;  wr_data_rom[ 9911]='h00000000;
    rd_cycle[ 9912] = 1'b0;  wr_cycle[ 9912] = 1'b1;  addr_rom[ 9912]='h00000b10;  wr_data_rom[ 9912]='h0000316f;
    rd_cycle[ 9913] = 1'b0;  wr_cycle[ 9913] = 1'b1;  addr_rom[ 9913]='h00000b70;  wr_data_rom[ 9913]='h00002e87;
    rd_cycle[ 9914] = 1'b1;  wr_cycle[ 9914] = 1'b0;  addr_rom[ 9914]='h00001270;  wr_data_rom[ 9914]='h00000000;
    rd_cycle[ 9915] = 1'b0;  wr_cycle[ 9915] = 1'b1;  addr_rom[ 9915]='h000021f0;  wr_data_rom[ 9915]='h0000108e;
    rd_cycle[ 9916] = 1'b1;  wr_cycle[ 9916] = 1'b0;  addr_rom[ 9916]='h000014b4;  wr_data_rom[ 9916]='h00000000;
    rd_cycle[ 9917] = 1'b1;  wr_cycle[ 9917] = 1'b0;  addr_rom[ 9917]='h00000c78;  wr_data_rom[ 9917]='h00000000;
    rd_cycle[ 9918] = 1'b1;  wr_cycle[ 9918] = 1'b0;  addr_rom[ 9918]='h00003630;  wr_data_rom[ 9918]='h00000000;
    rd_cycle[ 9919] = 1'b1;  wr_cycle[ 9919] = 1'b0;  addr_rom[ 9919]='h00001ed4;  wr_data_rom[ 9919]='h00000000;
    rd_cycle[ 9920] = 1'b0;  wr_cycle[ 9920] = 1'b1;  addr_rom[ 9920]='h00000c38;  wr_data_rom[ 9920]='h0000271e;
    rd_cycle[ 9921] = 1'b1;  wr_cycle[ 9921] = 1'b0;  addr_rom[ 9921]='h00002940;  wr_data_rom[ 9921]='h00000000;
    rd_cycle[ 9922] = 1'b0;  wr_cycle[ 9922] = 1'b1;  addr_rom[ 9922]='h000007a0;  wr_data_rom[ 9922]='h00002db5;
    rd_cycle[ 9923] = 1'b1;  wr_cycle[ 9923] = 1'b0;  addr_rom[ 9923]='h00002948;  wr_data_rom[ 9923]='h00000000;
    rd_cycle[ 9924] = 1'b1;  wr_cycle[ 9924] = 1'b0;  addr_rom[ 9924]='h00000988;  wr_data_rom[ 9924]='h00000000;
    rd_cycle[ 9925] = 1'b1;  wr_cycle[ 9925] = 1'b0;  addr_rom[ 9925]='h00000954;  wr_data_rom[ 9925]='h00000000;
    rd_cycle[ 9926] = 1'b1;  wr_cycle[ 9926] = 1'b0;  addr_rom[ 9926]='h00001ea4;  wr_data_rom[ 9926]='h00000000;
    rd_cycle[ 9927] = 1'b1;  wr_cycle[ 9927] = 1'b0;  addr_rom[ 9927]='h00000d6c;  wr_data_rom[ 9927]='h00000000;
    rd_cycle[ 9928] = 1'b1;  wr_cycle[ 9928] = 1'b0;  addr_rom[ 9928]='h00002c08;  wr_data_rom[ 9928]='h00000000;
    rd_cycle[ 9929] = 1'b0;  wr_cycle[ 9929] = 1'b1;  addr_rom[ 9929]='h00001bac;  wr_data_rom[ 9929]='h00002e97;
    rd_cycle[ 9930] = 1'b0;  wr_cycle[ 9930] = 1'b1;  addr_rom[ 9930]='h0000371c;  wr_data_rom[ 9930]='h00001e7f;
    rd_cycle[ 9931] = 1'b1;  wr_cycle[ 9931] = 1'b0;  addr_rom[ 9931]='h0000312c;  wr_data_rom[ 9931]='h00000000;
    rd_cycle[ 9932] = 1'b0;  wr_cycle[ 9932] = 1'b1;  addr_rom[ 9932]='h00003074;  wr_data_rom[ 9932]='h000026df;
    rd_cycle[ 9933] = 1'b0;  wr_cycle[ 9933] = 1'b1;  addr_rom[ 9933]='h00002650;  wr_data_rom[ 9933]='h000036ce;
    rd_cycle[ 9934] = 1'b1;  wr_cycle[ 9934] = 1'b0;  addr_rom[ 9934]='h00002ce8;  wr_data_rom[ 9934]='h00000000;
    rd_cycle[ 9935] = 1'b1;  wr_cycle[ 9935] = 1'b0;  addr_rom[ 9935]='h0000095c;  wr_data_rom[ 9935]='h00000000;
    rd_cycle[ 9936] = 1'b1;  wr_cycle[ 9936] = 1'b0;  addr_rom[ 9936]='h00000dfc;  wr_data_rom[ 9936]='h00000000;
    rd_cycle[ 9937] = 1'b1;  wr_cycle[ 9937] = 1'b0;  addr_rom[ 9937]='h00003cf0;  wr_data_rom[ 9937]='h00000000;
    rd_cycle[ 9938] = 1'b1;  wr_cycle[ 9938] = 1'b0;  addr_rom[ 9938]='h000010c4;  wr_data_rom[ 9938]='h00000000;
    rd_cycle[ 9939] = 1'b1;  wr_cycle[ 9939] = 1'b0;  addr_rom[ 9939]='h000019ec;  wr_data_rom[ 9939]='h00000000;
    rd_cycle[ 9940] = 1'b0;  wr_cycle[ 9940] = 1'b1;  addr_rom[ 9940]='h00001874;  wr_data_rom[ 9940]='h00003d55;
    rd_cycle[ 9941] = 1'b0;  wr_cycle[ 9941] = 1'b1;  addr_rom[ 9941]='h00001298;  wr_data_rom[ 9941]='h000008e7;
    rd_cycle[ 9942] = 1'b0;  wr_cycle[ 9942] = 1'b1;  addr_rom[ 9942]='h00002d60;  wr_data_rom[ 9942]='h00000d01;
    rd_cycle[ 9943] = 1'b0;  wr_cycle[ 9943] = 1'b1;  addr_rom[ 9943]='h00001264;  wr_data_rom[ 9943]='h0000348e;
    rd_cycle[ 9944] = 1'b0;  wr_cycle[ 9944] = 1'b1;  addr_rom[ 9944]='h00002574;  wr_data_rom[ 9944]='h000036c6;
    rd_cycle[ 9945] = 1'b0;  wr_cycle[ 9945] = 1'b1;  addr_rom[ 9945]='h00000864;  wr_data_rom[ 9945]='h00001e39;
    rd_cycle[ 9946] = 1'b0;  wr_cycle[ 9946] = 1'b1;  addr_rom[ 9946]='h00001988;  wr_data_rom[ 9946]='h0000175b;
    rd_cycle[ 9947] = 1'b1;  wr_cycle[ 9947] = 1'b0;  addr_rom[ 9947]='h00003afc;  wr_data_rom[ 9947]='h00000000;
    rd_cycle[ 9948] = 1'b0;  wr_cycle[ 9948] = 1'b1;  addr_rom[ 9948]='h00002c14;  wr_data_rom[ 9948]='h00002b6d;
    rd_cycle[ 9949] = 1'b0;  wr_cycle[ 9949] = 1'b1;  addr_rom[ 9949]='h000032b4;  wr_data_rom[ 9949]='h00002a2e;
    rd_cycle[ 9950] = 1'b1;  wr_cycle[ 9950] = 1'b0;  addr_rom[ 9950]='h000028ac;  wr_data_rom[ 9950]='h00000000;
    rd_cycle[ 9951] = 1'b1;  wr_cycle[ 9951] = 1'b0;  addr_rom[ 9951]='h00003180;  wr_data_rom[ 9951]='h00000000;
    rd_cycle[ 9952] = 1'b0;  wr_cycle[ 9952] = 1'b1;  addr_rom[ 9952]='h00002ea4;  wr_data_rom[ 9952]='h00003fa9;
    rd_cycle[ 9953] = 1'b1;  wr_cycle[ 9953] = 1'b0;  addr_rom[ 9953]='h00002054;  wr_data_rom[ 9953]='h00000000;
    rd_cycle[ 9954] = 1'b1;  wr_cycle[ 9954] = 1'b0;  addr_rom[ 9954]='h00001c70;  wr_data_rom[ 9954]='h00000000;
    rd_cycle[ 9955] = 1'b0;  wr_cycle[ 9955] = 1'b1;  addr_rom[ 9955]='h00002754;  wr_data_rom[ 9955]='h00003808;
    rd_cycle[ 9956] = 1'b0;  wr_cycle[ 9956] = 1'b1;  addr_rom[ 9956]='h00000ad4;  wr_data_rom[ 9956]='h0000250e;
    rd_cycle[ 9957] = 1'b0;  wr_cycle[ 9957] = 1'b1;  addr_rom[ 9957]='h00000df8;  wr_data_rom[ 9957]='h0000075a;
    rd_cycle[ 9958] = 1'b0;  wr_cycle[ 9958] = 1'b1;  addr_rom[ 9958]='h00002118;  wr_data_rom[ 9958]='h0000132f;
    rd_cycle[ 9959] = 1'b1;  wr_cycle[ 9959] = 1'b0;  addr_rom[ 9959]='h00001ce4;  wr_data_rom[ 9959]='h00000000;
    rd_cycle[ 9960] = 1'b0;  wr_cycle[ 9960] = 1'b1;  addr_rom[ 9960]='h00000bf8;  wr_data_rom[ 9960]='h000028e4;
    rd_cycle[ 9961] = 1'b0;  wr_cycle[ 9961] = 1'b1;  addr_rom[ 9961]='h00001e84;  wr_data_rom[ 9961]='h00003cb0;
    rd_cycle[ 9962] = 1'b1;  wr_cycle[ 9962] = 1'b0;  addr_rom[ 9962]='h00003334;  wr_data_rom[ 9962]='h00000000;
    rd_cycle[ 9963] = 1'b1;  wr_cycle[ 9963] = 1'b0;  addr_rom[ 9963]='h00000378;  wr_data_rom[ 9963]='h00000000;
    rd_cycle[ 9964] = 1'b1;  wr_cycle[ 9964] = 1'b0;  addr_rom[ 9964]='h0000216c;  wr_data_rom[ 9964]='h00000000;
    rd_cycle[ 9965] = 1'b1;  wr_cycle[ 9965] = 1'b0;  addr_rom[ 9965]='h00000518;  wr_data_rom[ 9965]='h00000000;
    rd_cycle[ 9966] = 1'b1;  wr_cycle[ 9966] = 1'b0;  addr_rom[ 9966]='h0000019c;  wr_data_rom[ 9966]='h00000000;
    rd_cycle[ 9967] = 1'b1;  wr_cycle[ 9967] = 1'b0;  addr_rom[ 9967]='h000001b0;  wr_data_rom[ 9967]='h00000000;
    rd_cycle[ 9968] = 1'b0;  wr_cycle[ 9968] = 1'b1;  addr_rom[ 9968]='h00001444;  wr_data_rom[ 9968]='h000021ba;
    rd_cycle[ 9969] = 1'b1;  wr_cycle[ 9969] = 1'b0;  addr_rom[ 9969]='h00002890;  wr_data_rom[ 9969]='h00000000;
    rd_cycle[ 9970] = 1'b0;  wr_cycle[ 9970] = 1'b1;  addr_rom[ 9970]='h000028cc;  wr_data_rom[ 9970]='h00003b76;
    rd_cycle[ 9971] = 1'b0;  wr_cycle[ 9971] = 1'b1;  addr_rom[ 9971]='h0000065c;  wr_data_rom[ 9971]='h0000241c;
    rd_cycle[ 9972] = 1'b1;  wr_cycle[ 9972] = 1'b0;  addr_rom[ 9972]='h00003308;  wr_data_rom[ 9972]='h00000000;
    rd_cycle[ 9973] = 1'b0;  wr_cycle[ 9973] = 1'b1;  addr_rom[ 9973]='h000008cc;  wr_data_rom[ 9973]='h00002807;
    rd_cycle[ 9974] = 1'b1;  wr_cycle[ 9974] = 1'b0;  addr_rom[ 9974]='h00003b7c;  wr_data_rom[ 9974]='h00000000;
    rd_cycle[ 9975] = 1'b1;  wr_cycle[ 9975] = 1'b0;  addr_rom[ 9975]='h00001048;  wr_data_rom[ 9975]='h00000000;
    rd_cycle[ 9976] = 1'b0;  wr_cycle[ 9976] = 1'b1;  addr_rom[ 9976]='h00000038;  wr_data_rom[ 9976]='h00001aeb;
    rd_cycle[ 9977] = 1'b1;  wr_cycle[ 9977] = 1'b0;  addr_rom[ 9977]='h0000160c;  wr_data_rom[ 9977]='h00000000;
    rd_cycle[ 9978] = 1'b0;  wr_cycle[ 9978] = 1'b1;  addr_rom[ 9978]='h00002530;  wr_data_rom[ 9978]='h00002046;
    rd_cycle[ 9979] = 1'b1;  wr_cycle[ 9979] = 1'b0;  addr_rom[ 9979]='h00001c0c;  wr_data_rom[ 9979]='h00000000;
    rd_cycle[ 9980] = 1'b0;  wr_cycle[ 9980] = 1'b1;  addr_rom[ 9980]='h000008a0;  wr_data_rom[ 9980]='h0000204f;
    rd_cycle[ 9981] = 1'b0;  wr_cycle[ 9981] = 1'b1;  addr_rom[ 9981]='h00001b9c;  wr_data_rom[ 9981]='h00002802;
    rd_cycle[ 9982] = 1'b1;  wr_cycle[ 9982] = 1'b0;  addr_rom[ 9982]='h00001e24;  wr_data_rom[ 9982]='h00000000;
    rd_cycle[ 9983] = 1'b0;  wr_cycle[ 9983] = 1'b1;  addr_rom[ 9983]='h00003d3c;  wr_data_rom[ 9983]='h00002bff;
    rd_cycle[ 9984] = 1'b1;  wr_cycle[ 9984] = 1'b0;  addr_rom[ 9984]='h000017bc;  wr_data_rom[ 9984]='h00000000;
    rd_cycle[ 9985] = 1'b1;  wr_cycle[ 9985] = 1'b0;  addr_rom[ 9985]='h000008e8;  wr_data_rom[ 9985]='h00000000;
    rd_cycle[ 9986] = 1'b1;  wr_cycle[ 9986] = 1'b0;  addr_rom[ 9986]='h00001b78;  wr_data_rom[ 9986]='h00000000;
    rd_cycle[ 9987] = 1'b1;  wr_cycle[ 9987] = 1'b0;  addr_rom[ 9987]='h00002104;  wr_data_rom[ 9987]='h00000000;
    rd_cycle[ 9988] = 1'b1;  wr_cycle[ 9988] = 1'b0;  addr_rom[ 9988]='h00003768;  wr_data_rom[ 9988]='h00000000;
    rd_cycle[ 9989] = 1'b1;  wr_cycle[ 9989] = 1'b0;  addr_rom[ 9989]='h000007f8;  wr_data_rom[ 9989]='h00000000;
    rd_cycle[ 9990] = 1'b1;  wr_cycle[ 9990] = 1'b0;  addr_rom[ 9990]='h0000247c;  wr_data_rom[ 9990]='h00000000;
    rd_cycle[ 9991] = 1'b0;  wr_cycle[ 9991] = 1'b1;  addr_rom[ 9991]='h00002ce8;  wr_data_rom[ 9991]='h0000034f;
    rd_cycle[ 9992] = 1'b0;  wr_cycle[ 9992] = 1'b1;  addr_rom[ 9992]='h000039cc;  wr_data_rom[ 9992]='h00001338;
    rd_cycle[ 9993] = 1'b1;  wr_cycle[ 9993] = 1'b0;  addr_rom[ 9993]='h000034dc;  wr_data_rom[ 9993]='h00000000;
    rd_cycle[ 9994] = 1'b0;  wr_cycle[ 9994] = 1'b1;  addr_rom[ 9994]='h00000a40;  wr_data_rom[ 9994]='h00003fc2;
    rd_cycle[ 9995] = 1'b0;  wr_cycle[ 9995] = 1'b1;  addr_rom[ 9995]='h000024bc;  wr_data_rom[ 9995]='h00000714;
    rd_cycle[ 9996] = 1'b1;  wr_cycle[ 9996] = 1'b0;  addr_rom[ 9996]='h00001304;  wr_data_rom[ 9996]='h00000000;
    rd_cycle[ 9997] = 1'b1;  wr_cycle[ 9997] = 1'b0;  addr_rom[ 9997]='h000034e8;  wr_data_rom[ 9997]='h00000000;
    rd_cycle[ 9998] = 1'b0;  wr_cycle[ 9998] = 1'b1;  addr_rom[ 9998]='h00000258;  wr_data_rom[ 9998]='h00003ca7;
    rd_cycle[ 9999] = 1'b0;  wr_cycle[ 9999] = 1'b1;  addr_rom[ 9999]='h0000185c;  wr_data_rom[ 9999]='h000035e3;
    rd_cycle[10000] = 1'b1;  wr_cycle[10000] = 1'b0;  addr_rom[10000]='h000027c8;  wr_data_rom[10000]='h00000000;
    rd_cycle[10001] = 1'b1;  wr_cycle[10001] = 1'b0;  addr_rom[10001]='h000001f8;  wr_data_rom[10001]='h00000000;
    rd_cycle[10002] = 1'b0;  wr_cycle[10002] = 1'b1;  addr_rom[10002]='h00001ad8;  wr_data_rom[10002]='h0000323f;
    rd_cycle[10003] = 1'b0;  wr_cycle[10003] = 1'b1;  addr_rom[10003]='h000020c4;  wr_data_rom[10003]='h00003969;
    rd_cycle[10004] = 1'b1;  wr_cycle[10004] = 1'b0;  addr_rom[10004]='h000021d8;  wr_data_rom[10004]='h00000000;
    rd_cycle[10005] = 1'b1;  wr_cycle[10005] = 1'b0;  addr_rom[10005]='h00002b08;  wr_data_rom[10005]='h00000000;
    rd_cycle[10006] = 1'b0;  wr_cycle[10006] = 1'b1;  addr_rom[10006]='h00002544;  wr_data_rom[10006]='h00002b0e;
    rd_cycle[10007] = 1'b1;  wr_cycle[10007] = 1'b0;  addr_rom[10007]='h00002048;  wr_data_rom[10007]='h00000000;
    rd_cycle[10008] = 1'b0;  wr_cycle[10008] = 1'b1;  addr_rom[10008]='h000003a8;  wr_data_rom[10008]='h00001fe3;
    rd_cycle[10009] = 1'b0;  wr_cycle[10009] = 1'b1;  addr_rom[10009]='h00000488;  wr_data_rom[10009]='h00002a6e;
    rd_cycle[10010] = 1'b1;  wr_cycle[10010] = 1'b0;  addr_rom[10010]='h00000e70;  wr_data_rom[10010]='h00000000;
    rd_cycle[10011] = 1'b0;  wr_cycle[10011] = 1'b1;  addr_rom[10011]='h000021f4;  wr_data_rom[10011]='h000013f8;
    rd_cycle[10012] = 1'b0;  wr_cycle[10012] = 1'b1;  addr_rom[10012]='h00001cb0;  wr_data_rom[10012]='h00001131;
    rd_cycle[10013] = 1'b1;  wr_cycle[10013] = 1'b0;  addr_rom[10013]='h00003458;  wr_data_rom[10013]='h00000000;
    rd_cycle[10014] = 1'b0;  wr_cycle[10014] = 1'b1;  addr_rom[10014]='h00003d84;  wr_data_rom[10014]='h00000d3c;
    rd_cycle[10015] = 1'b1;  wr_cycle[10015] = 1'b0;  addr_rom[10015]='h00002d54;  wr_data_rom[10015]='h00000000;
    rd_cycle[10016] = 1'b1;  wr_cycle[10016] = 1'b0;  addr_rom[10016]='h00000934;  wr_data_rom[10016]='h00000000;
    rd_cycle[10017] = 1'b0;  wr_cycle[10017] = 1'b1;  addr_rom[10017]='h00001c28;  wr_data_rom[10017]='h000001c6;
    rd_cycle[10018] = 1'b1;  wr_cycle[10018] = 1'b0;  addr_rom[10018]='h00000434;  wr_data_rom[10018]='h00000000;
    rd_cycle[10019] = 1'b1;  wr_cycle[10019] = 1'b0;  addr_rom[10019]='h00003a0c;  wr_data_rom[10019]='h00000000;
    rd_cycle[10020] = 1'b1;  wr_cycle[10020] = 1'b0;  addr_rom[10020]='h00001598;  wr_data_rom[10020]='h00000000;
    rd_cycle[10021] = 1'b1;  wr_cycle[10021] = 1'b0;  addr_rom[10021]='h000002cc;  wr_data_rom[10021]='h00000000;
    rd_cycle[10022] = 1'b1;  wr_cycle[10022] = 1'b0;  addr_rom[10022]='h000031dc;  wr_data_rom[10022]='h00000000;
    rd_cycle[10023] = 1'b0;  wr_cycle[10023] = 1'b1;  addr_rom[10023]='h000029e4;  wr_data_rom[10023]='h00002a48;
    rd_cycle[10024] = 1'b0;  wr_cycle[10024] = 1'b1;  addr_rom[10024]='h000007d4;  wr_data_rom[10024]='h0000088b;
    rd_cycle[10025] = 1'b1;  wr_cycle[10025] = 1'b0;  addr_rom[10025]='h00001020;  wr_data_rom[10025]='h00000000;
    rd_cycle[10026] = 1'b1;  wr_cycle[10026] = 1'b0;  addr_rom[10026]='h00001c58;  wr_data_rom[10026]='h00000000;
    rd_cycle[10027] = 1'b0;  wr_cycle[10027] = 1'b1;  addr_rom[10027]='h00001898;  wr_data_rom[10027]='h000006cf;
    rd_cycle[10028] = 1'b1;  wr_cycle[10028] = 1'b0;  addr_rom[10028]='h00003e3c;  wr_data_rom[10028]='h00000000;
    rd_cycle[10029] = 1'b1;  wr_cycle[10029] = 1'b0;  addr_rom[10029]='h000033b0;  wr_data_rom[10029]='h00000000;
    rd_cycle[10030] = 1'b1;  wr_cycle[10030] = 1'b0;  addr_rom[10030]='h00000bb4;  wr_data_rom[10030]='h00000000;
    rd_cycle[10031] = 1'b1;  wr_cycle[10031] = 1'b0;  addr_rom[10031]='h000023c4;  wr_data_rom[10031]='h00000000;
    rd_cycle[10032] = 1'b0;  wr_cycle[10032] = 1'b1;  addr_rom[10032]='h00003390;  wr_data_rom[10032]='h00001b01;
    rd_cycle[10033] = 1'b0;  wr_cycle[10033] = 1'b1;  addr_rom[10033]='h000021ec;  wr_data_rom[10033]='h00000ef0;
    rd_cycle[10034] = 1'b1;  wr_cycle[10034] = 1'b0;  addr_rom[10034]='h000036c4;  wr_data_rom[10034]='h00000000;
    rd_cycle[10035] = 1'b0;  wr_cycle[10035] = 1'b1;  addr_rom[10035]='h00002164;  wr_data_rom[10035]='h0000325d;
    rd_cycle[10036] = 1'b0;  wr_cycle[10036] = 1'b1;  addr_rom[10036]='h00000b24;  wr_data_rom[10036]='h000018a2;
    rd_cycle[10037] = 1'b1;  wr_cycle[10037] = 1'b0;  addr_rom[10037]='h000034dc;  wr_data_rom[10037]='h00000000;
    rd_cycle[10038] = 1'b1;  wr_cycle[10038] = 1'b0;  addr_rom[10038]='h0000011c;  wr_data_rom[10038]='h00000000;
    rd_cycle[10039] = 1'b1;  wr_cycle[10039] = 1'b0;  addr_rom[10039]='h00003b78;  wr_data_rom[10039]='h00000000;
    rd_cycle[10040] = 1'b0;  wr_cycle[10040] = 1'b1;  addr_rom[10040]='h00001770;  wr_data_rom[10040]='h00002bf9;
    rd_cycle[10041] = 1'b0;  wr_cycle[10041] = 1'b1;  addr_rom[10041]='h00000a54;  wr_data_rom[10041]='h000032fc;
    rd_cycle[10042] = 1'b0;  wr_cycle[10042] = 1'b1;  addr_rom[10042]='h00001b74;  wr_data_rom[10042]='h00002d82;
    rd_cycle[10043] = 1'b0;  wr_cycle[10043] = 1'b1;  addr_rom[10043]='h00001f08;  wr_data_rom[10043]='h000009b5;
    rd_cycle[10044] = 1'b0;  wr_cycle[10044] = 1'b1;  addr_rom[10044]='h000038e8;  wr_data_rom[10044]='h0000061b;
    rd_cycle[10045] = 1'b1;  wr_cycle[10045] = 1'b0;  addr_rom[10045]='h00002fcc;  wr_data_rom[10045]='h00000000;
    rd_cycle[10046] = 1'b0;  wr_cycle[10046] = 1'b1;  addr_rom[10046]='h00002d60;  wr_data_rom[10046]='h00003bc3;
    rd_cycle[10047] = 1'b0;  wr_cycle[10047] = 1'b1;  addr_rom[10047]='h00001b5c;  wr_data_rom[10047]='h00000db8;
    rd_cycle[10048] = 1'b1;  wr_cycle[10048] = 1'b0;  addr_rom[10048]='h00003b18;  wr_data_rom[10048]='h00000000;
    rd_cycle[10049] = 1'b1;  wr_cycle[10049] = 1'b0;  addr_rom[10049]='h00000328;  wr_data_rom[10049]='h00000000;
    rd_cycle[10050] = 1'b1;  wr_cycle[10050] = 1'b0;  addr_rom[10050]='h000002c0;  wr_data_rom[10050]='h00000000;
    rd_cycle[10051] = 1'b1;  wr_cycle[10051] = 1'b0;  addr_rom[10051]='h0000293c;  wr_data_rom[10051]='h00000000;
    rd_cycle[10052] = 1'b0;  wr_cycle[10052] = 1'b1;  addr_rom[10052]='h00000c30;  wr_data_rom[10052]='h00000c6d;
    rd_cycle[10053] = 1'b1;  wr_cycle[10053] = 1'b0;  addr_rom[10053]='h00003cc8;  wr_data_rom[10053]='h00000000;
    rd_cycle[10054] = 1'b0;  wr_cycle[10054] = 1'b1;  addr_rom[10054]='h00003d64;  wr_data_rom[10054]='h00002b5f;
    rd_cycle[10055] = 1'b0;  wr_cycle[10055] = 1'b1;  addr_rom[10055]='h000027b4;  wr_data_rom[10055]='h00002412;
    rd_cycle[10056] = 1'b1;  wr_cycle[10056] = 1'b0;  addr_rom[10056]='h00001924;  wr_data_rom[10056]='h00000000;
    rd_cycle[10057] = 1'b0;  wr_cycle[10057] = 1'b1;  addr_rom[10057]='h00001784;  wr_data_rom[10057]='h00001d70;
    rd_cycle[10058] = 1'b0;  wr_cycle[10058] = 1'b1;  addr_rom[10058]='h00003348;  wr_data_rom[10058]='h00003707;
    rd_cycle[10059] = 1'b1;  wr_cycle[10059] = 1'b0;  addr_rom[10059]='h00001808;  wr_data_rom[10059]='h00000000;
    rd_cycle[10060] = 1'b1;  wr_cycle[10060] = 1'b0;  addr_rom[10060]='h00002a4c;  wr_data_rom[10060]='h00000000;
    rd_cycle[10061] = 1'b0;  wr_cycle[10061] = 1'b1;  addr_rom[10061]='h0000392c;  wr_data_rom[10061]='h00001b67;
    rd_cycle[10062] = 1'b1;  wr_cycle[10062] = 1'b0;  addr_rom[10062]='h00003a80;  wr_data_rom[10062]='h00000000;
    rd_cycle[10063] = 1'b1;  wr_cycle[10063] = 1'b0;  addr_rom[10063]='h00003680;  wr_data_rom[10063]='h00000000;
    rd_cycle[10064] = 1'b1;  wr_cycle[10064] = 1'b0;  addr_rom[10064]='h000037ac;  wr_data_rom[10064]='h00000000;
    rd_cycle[10065] = 1'b0;  wr_cycle[10065] = 1'b1;  addr_rom[10065]='h00002768;  wr_data_rom[10065]='h00003d39;
    rd_cycle[10066] = 1'b0;  wr_cycle[10066] = 1'b1;  addr_rom[10066]='h00002c2c;  wr_data_rom[10066]='h00003feb;
    rd_cycle[10067] = 1'b0;  wr_cycle[10067] = 1'b1;  addr_rom[10067]='h00000cd4;  wr_data_rom[10067]='h00003da4;
    rd_cycle[10068] = 1'b0;  wr_cycle[10068] = 1'b1;  addr_rom[10068]='h00003f3c;  wr_data_rom[10068]='h00000038;
    rd_cycle[10069] = 1'b1;  wr_cycle[10069] = 1'b0;  addr_rom[10069]='h000039d4;  wr_data_rom[10069]='h00000000;
    rd_cycle[10070] = 1'b0;  wr_cycle[10070] = 1'b1;  addr_rom[10070]='h00000998;  wr_data_rom[10070]='h00003be1;
    rd_cycle[10071] = 1'b1;  wr_cycle[10071] = 1'b0;  addr_rom[10071]='h00003bd8;  wr_data_rom[10071]='h00000000;
    rd_cycle[10072] = 1'b1;  wr_cycle[10072] = 1'b0;  addr_rom[10072]='h00002e3c;  wr_data_rom[10072]='h00000000;
    rd_cycle[10073] = 1'b0;  wr_cycle[10073] = 1'b1;  addr_rom[10073]='h00003ea4;  wr_data_rom[10073]='h00001b38;
    rd_cycle[10074] = 1'b0;  wr_cycle[10074] = 1'b1;  addr_rom[10074]='h00001b18;  wr_data_rom[10074]='h00000025;
    rd_cycle[10075] = 1'b0;  wr_cycle[10075] = 1'b1;  addr_rom[10075]='h00001a58;  wr_data_rom[10075]='h000010fd;
    rd_cycle[10076] = 1'b0;  wr_cycle[10076] = 1'b1;  addr_rom[10076]='h00002c6c;  wr_data_rom[10076]='h00000408;
    rd_cycle[10077] = 1'b1;  wr_cycle[10077] = 1'b0;  addr_rom[10077]='h00002554;  wr_data_rom[10077]='h00000000;
    rd_cycle[10078] = 1'b0;  wr_cycle[10078] = 1'b1;  addr_rom[10078]='h00002ed4;  wr_data_rom[10078]='h000018f4;
    rd_cycle[10079] = 1'b1;  wr_cycle[10079] = 1'b0;  addr_rom[10079]='h0000294c;  wr_data_rom[10079]='h00000000;
    rd_cycle[10080] = 1'b1;  wr_cycle[10080] = 1'b0;  addr_rom[10080]='h000001b4;  wr_data_rom[10080]='h00000000;
    rd_cycle[10081] = 1'b0;  wr_cycle[10081] = 1'b1;  addr_rom[10081]='h00001850;  wr_data_rom[10081]='h00000edf;
    rd_cycle[10082] = 1'b1;  wr_cycle[10082] = 1'b0;  addr_rom[10082]='h000006d0;  wr_data_rom[10082]='h00000000;
    rd_cycle[10083] = 1'b1;  wr_cycle[10083] = 1'b0;  addr_rom[10083]='h000038c4;  wr_data_rom[10083]='h00000000;
    rd_cycle[10084] = 1'b0;  wr_cycle[10084] = 1'b1;  addr_rom[10084]='h0000144c;  wr_data_rom[10084]='h0000164b;
    rd_cycle[10085] = 1'b1;  wr_cycle[10085] = 1'b0;  addr_rom[10085]='h0000108c;  wr_data_rom[10085]='h00000000;
    rd_cycle[10086] = 1'b0;  wr_cycle[10086] = 1'b1;  addr_rom[10086]='h00001508;  wr_data_rom[10086]='h000003ba;
    rd_cycle[10087] = 1'b1;  wr_cycle[10087] = 1'b0;  addr_rom[10087]='h00002cec;  wr_data_rom[10087]='h00000000;
    rd_cycle[10088] = 1'b0;  wr_cycle[10088] = 1'b1;  addr_rom[10088]='h0000368c;  wr_data_rom[10088]='h000002c1;
    rd_cycle[10089] = 1'b0;  wr_cycle[10089] = 1'b1;  addr_rom[10089]='h000027f8;  wr_data_rom[10089]='h00003b5e;
    rd_cycle[10090] = 1'b1;  wr_cycle[10090] = 1'b0;  addr_rom[10090]='h00001578;  wr_data_rom[10090]='h00000000;
    rd_cycle[10091] = 1'b1;  wr_cycle[10091] = 1'b0;  addr_rom[10091]='h00002cd0;  wr_data_rom[10091]='h00000000;
    rd_cycle[10092] = 1'b0;  wr_cycle[10092] = 1'b1;  addr_rom[10092]='h00002944;  wr_data_rom[10092]='h00001f7b;
    rd_cycle[10093] = 1'b0;  wr_cycle[10093] = 1'b1;  addr_rom[10093]='h00003960;  wr_data_rom[10093]='h000022db;
    rd_cycle[10094] = 1'b1;  wr_cycle[10094] = 1'b0;  addr_rom[10094]='h00003758;  wr_data_rom[10094]='h00000000;
    rd_cycle[10095] = 1'b0;  wr_cycle[10095] = 1'b1;  addr_rom[10095]='h00003b54;  wr_data_rom[10095]='h0000232a;
    rd_cycle[10096] = 1'b0;  wr_cycle[10096] = 1'b1;  addr_rom[10096]='h00003d08;  wr_data_rom[10096]='h00000620;
    rd_cycle[10097] = 1'b1;  wr_cycle[10097] = 1'b0;  addr_rom[10097]='h00000630;  wr_data_rom[10097]='h00000000;
    rd_cycle[10098] = 1'b1;  wr_cycle[10098] = 1'b0;  addr_rom[10098]='h000018f8;  wr_data_rom[10098]='h00000000;
    rd_cycle[10099] = 1'b0;  wr_cycle[10099] = 1'b1;  addr_rom[10099]='h00001dc0;  wr_data_rom[10099]='h00002e62;
    rd_cycle[10100] = 1'b0;  wr_cycle[10100] = 1'b1;  addr_rom[10100]='h00003dc8;  wr_data_rom[10100]='h00001bd3;
    rd_cycle[10101] = 1'b1;  wr_cycle[10101] = 1'b0;  addr_rom[10101]='h000010b8;  wr_data_rom[10101]='h00000000;
    rd_cycle[10102] = 1'b1;  wr_cycle[10102] = 1'b0;  addr_rom[10102]='h00001374;  wr_data_rom[10102]='h00000000;
    rd_cycle[10103] = 1'b1;  wr_cycle[10103] = 1'b0;  addr_rom[10103]='h00001824;  wr_data_rom[10103]='h00000000;
    rd_cycle[10104] = 1'b0;  wr_cycle[10104] = 1'b1;  addr_rom[10104]='h00001d98;  wr_data_rom[10104]='h0000117d;
    rd_cycle[10105] = 1'b1;  wr_cycle[10105] = 1'b0;  addr_rom[10105]='h00002334;  wr_data_rom[10105]='h00000000;
    rd_cycle[10106] = 1'b1;  wr_cycle[10106] = 1'b0;  addr_rom[10106]='h00003694;  wr_data_rom[10106]='h00000000;
    rd_cycle[10107] = 1'b0;  wr_cycle[10107] = 1'b1;  addr_rom[10107]='h00002938;  wr_data_rom[10107]='h000029b3;
    rd_cycle[10108] = 1'b1;  wr_cycle[10108] = 1'b0;  addr_rom[10108]='h00002ce8;  wr_data_rom[10108]='h00000000;
    rd_cycle[10109] = 1'b1;  wr_cycle[10109] = 1'b0;  addr_rom[10109]='h00001330;  wr_data_rom[10109]='h00000000;
    rd_cycle[10110] = 1'b0;  wr_cycle[10110] = 1'b1;  addr_rom[10110]='h000012d8;  wr_data_rom[10110]='h00002572;
    rd_cycle[10111] = 1'b0;  wr_cycle[10111] = 1'b1;  addr_rom[10111]='h00003370;  wr_data_rom[10111]='h00002488;
    rd_cycle[10112] = 1'b1;  wr_cycle[10112] = 1'b0;  addr_rom[10112]='h00002cf8;  wr_data_rom[10112]='h00000000;
    rd_cycle[10113] = 1'b1;  wr_cycle[10113] = 1'b0;  addr_rom[10113]='h00003d60;  wr_data_rom[10113]='h00000000;
    rd_cycle[10114] = 1'b1;  wr_cycle[10114] = 1'b0;  addr_rom[10114]='h000015d8;  wr_data_rom[10114]='h00000000;
    rd_cycle[10115] = 1'b0;  wr_cycle[10115] = 1'b1;  addr_rom[10115]='h00001398;  wr_data_rom[10115]='h0000298e;
    rd_cycle[10116] = 1'b0;  wr_cycle[10116] = 1'b1;  addr_rom[10116]='h0000093c;  wr_data_rom[10116]='h00001a5b;
    rd_cycle[10117] = 1'b1;  wr_cycle[10117] = 1'b0;  addr_rom[10117]='h00003060;  wr_data_rom[10117]='h00000000;
    rd_cycle[10118] = 1'b0;  wr_cycle[10118] = 1'b1;  addr_rom[10118]='h000010c8;  wr_data_rom[10118]='h00000e27;
    rd_cycle[10119] = 1'b1;  wr_cycle[10119] = 1'b0;  addr_rom[10119]='h00003d6c;  wr_data_rom[10119]='h00000000;
    rd_cycle[10120] = 1'b1;  wr_cycle[10120] = 1'b0;  addr_rom[10120]='h00002020;  wr_data_rom[10120]='h00000000;
    rd_cycle[10121] = 1'b1;  wr_cycle[10121] = 1'b0;  addr_rom[10121]='h00003270;  wr_data_rom[10121]='h00000000;
    rd_cycle[10122] = 1'b0;  wr_cycle[10122] = 1'b1;  addr_rom[10122]='h00002788;  wr_data_rom[10122]='h00003816;
    rd_cycle[10123] = 1'b1;  wr_cycle[10123] = 1'b0;  addr_rom[10123]='h00000ce4;  wr_data_rom[10123]='h00000000;
    rd_cycle[10124] = 1'b0;  wr_cycle[10124] = 1'b1;  addr_rom[10124]='h00000f40;  wr_data_rom[10124]='h00002b95;
    rd_cycle[10125] = 1'b1;  wr_cycle[10125] = 1'b0;  addr_rom[10125]='h0000156c;  wr_data_rom[10125]='h00000000;
    rd_cycle[10126] = 1'b1;  wr_cycle[10126] = 1'b0;  addr_rom[10126]='h00001da8;  wr_data_rom[10126]='h00000000;
    rd_cycle[10127] = 1'b0;  wr_cycle[10127] = 1'b1;  addr_rom[10127]='h0000312c;  wr_data_rom[10127]='h00000e3f;
    rd_cycle[10128] = 1'b0;  wr_cycle[10128] = 1'b1;  addr_rom[10128]='h00002e64;  wr_data_rom[10128]='h000009db;
    rd_cycle[10129] = 1'b0;  wr_cycle[10129] = 1'b1;  addr_rom[10129]='h00003e1c;  wr_data_rom[10129]='h0000347d;
    rd_cycle[10130] = 1'b1;  wr_cycle[10130] = 1'b0;  addr_rom[10130]='h00003794;  wr_data_rom[10130]='h00000000;
    rd_cycle[10131] = 1'b1;  wr_cycle[10131] = 1'b0;  addr_rom[10131]='h00002bb8;  wr_data_rom[10131]='h00000000;
    rd_cycle[10132] = 1'b0;  wr_cycle[10132] = 1'b1;  addr_rom[10132]='h000017c0;  wr_data_rom[10132]='h000028d4;
    rd_cycle[10133] = 1'b0;  wr_cycle[10133] = 1'b1;  addr_rom[10133]='h00000cd0;  wr_data_rom[10133]='h00002f7c;
    rd_cycle[10134] = 1'b1;  wr_cycle[10134] = 1'b0;  addr_rom[10134]='h00001878;  wr_data_rom[10134]='h00000000;
    rd_cycle[10135] = 1'b1;  wr_cycle[10135] = 1'b0;  addr_rom[10135]='h00003c88;  wr_data_rom[10135]='h00000000;
    rd_cycle[10136] = 1'b0;  wr_cycle[10136] = 1'b1;  addr_rom[10136]='h00003798;  wr_data_rom[10136]='h00003bac;
    rd_cycle[10137] = 1'b0;  wr_cycle[10137] = 1'b1;  addr_rom[10137]='h00003aec;  wr_data_rom[10137]='h00001452;
    rd_cycle[10138] = 1'b1;  wr_cycle[10138] = 1'b0;  addr_rom[10138]='h00000e54;  wr_data_rom[10138]='h00000000;
    rd_cycle[10139] = 1'b0;  wr_cycle[10139] = 1'b1;  addr_rom[10139]='h00000848;  wr_data_rom[10139]='h00003f31;
    rd_cycle[10140] = 1'b1;  wr_cycle[10140] = 1'b0;  addr_rom[10140]='h0000060c;  wr_data_rom[10140]='h00000000;
    rd_cycle[10141] = 1'b0;  wr_cycle[10141] = 1'b1;  addr_rom[10141]='h00000424;  wr_data_rom[10141]='h00000b88;
    rd_cycle[10142] = 1'b1;  wr_cycle[10142] = 1'b0;  addr_rom[10142]='h000024ec;  wr_data_rom[10142]='h00000000;
    rd_cycle[10143] = 1'b0;  wr_cycle[10143] = 1'b1;  addr_rom[10143]='h000031d4;  wr_data_rom[10143]='h0000345e;
    rd_cycle[10144] = 1'b1;  wr_cycle[10144] = 1'b0;  addr_rom[10144]='h00003e44;  wr_data_rom[10144]='h00000000;
    rd_cycle[10145] = 1'b0;  wr_cycle[10145] = 1'b1;  addr_rom[10145]='h00003fd4;  wr_data_rom[10145]='h00000d20;
    rd_cycle[10146] = 1'b0;  wr_cycle[10146] = 1'b1;  addr_rom[10146]='h00000888;  wr_data_rom[10146]='h000029d0;
    rd_cycle[10147] = 1'b0;  wr_cycle[10147] = 1'b1;  addr_rom[10147]='h0000253c;  wr_data_rom[10147]='h00003fd8;
    rd_cycle[10148] = 1'b0;  wr_cycle[10148] = 1'b1;  addr_rom[10148]='h00002090;  wr_data_rom[10148]='h000029b4;
    rd_cycle[10149] = 1'b0;  wr_cycle[10149] = 1'b1;  addr_rom[10149]='h000037f0;  wr_data_rom[10149]='h00001c06;
    rd_cycle[10150] = 1'b1;  wr_cycle[10150] = 1'b0;  addr_rom[10150]='h00003bc0;  wr_data_rom[10150]='h00000000;
    rd_cycle[10151] = 1'b0;  wr_cycle[10151] = 1'b1;  addr_rom[10151]='h00000cb4;  wr_data_rom[10151]='h0000124f;
    rd_cycle[10152] = 1'b1;  wr_cycle[10152] = 1'b0;  addr_rom[10152]='h00002e88;  wr_data_rom[10152]='h00000000;
    rd_cycle[10153] = 1'b1;  wr_cycle[10153] = 1'b0;  addr_rom[10153]='h00000eac;  wr_data_rom[10153]='h00000000;
    rd_cycle[10154] = 1'b1;  wr_cycle[10154] = 1'b0;  addr_rom[10154]='h0000369c;  wr_data_rom[10154]='h00000000;
    rd_cycle[10155] = 1'b0;  wr_cycle[10155] = 1'b1;  addr_rom[10155]='h00002738;  wr_data_rom[10155]='h00002b07;
    rd_cycle[10156] = 1'b0;  wr_cycle[10156] = 1'b1;  addr_rom[10156]='h00001734;  wr_data_rom[10156]='h0000295e;
    rd_cycle[10157] = 1'b1;  wr_cycle[10157] = 1'b0;  addr_rom[10157]='h00000628;  wr_data_rom[10157]='h00000000;
    rd_cycle[10158] = 1'b0;  wr_cycle[10158] = 1'b1;  addr_rom[10158]='h00002004;  wr_data_rom[10158]='h000015a4;
    rd_cycle[10159] = 1'b1;  wr_cycle[10159] = 1'b0;  addr_rom[10159]='h00001eac;  wr_data_rom[10159]='h00000000;
    rd_cycle[10160] = 1'b1;  wr_cycle[10160] = 1'b0;  addr_rom[10160]='h00001e78;  wr_data_rom[10160]='h00000000;
    rd_cycle[10161] = 1'b0;  wr_cycle[10161] = 1'b1;  addr_rom[10161]='h00003f1c;  wr_data_rom[10161]='h000020b8;
    rd_cycle[10162] = 1'b1;  wr_cycle[10162] = 1'b0;  addr_rom[10162]='h0000148c;  wr_data_rom[10162]='h00000000;
    rd_cycle[10163] = 1'b1;  wr_cycle[10163] = 1'b0;  addr_rom[10163]='h000014dc;  wr_data_rom[10163]='h00000000;
    rd_cycle[10164] = 1'b1;  wr_cycle[10164] = 1'b0;  addr_rom[10164]='h00001d54;  wr_data_rom[10164]='h00000000;
    rd_cycle[10165] = 1'b1;  wr_cycle[10165] = 1'b0;  addr_rom[10165]='h00001b28;  wr_data_rom[10165]='h00000000;
    rd_cycle[10166] = 1'b1;  wr_cycle[10166] = 1'b0;  addr_rom[10166]='h00000cf8;  wr_data_rom[10166]='h00000000;
    rd_cycle[10167] = 1'b1;  wr_cycle[10167] = 1'b0;  addr_rom[10167]='h00002030;  wr_data_rom[10167]='h00000000;
    rd_cycle[10168] = 1'b1;  wr_cycle[10168] = 1'b0;  addr_rom[10168]='h0000250c;  wr_data_rom[10168]='h00000000;
    rd_cycle[10169] = 1'b1;  wr_cycle[10169] = 1'b0;  addr_rom[10169]='h00000738;  wr_data_rom[10169]='h00000000;
    rd_cycle[10170] = 1'b1;  wr_cycle[10170] = 1'b0;  addr_rom[10170]='h00002610;  wr_data_rom[10170]='h00000000;
    rd_cycle[10171] = 1'b0;  wr_cycle[10171] = 1'b1;  addr_rom[10171]='h00001c30;  wr_data_rom[10171]='h00003d7a;
    rd_cycle[10172] = 1'b1;  wr_cycle[10172] = 1'b0;  addr_rom[10172]='h000016c0;  wr_data_rom[10172]='h00000000;
    rd_cycle[10173] = 1'b1;  wr_cycle[10173] = 1'b0;  addr_rom[10173]='h0000050c;  wr_data_rom[10173]='h00000000;
    rd_cycle[10174] = 1'b1;  wr_cycle[10174] = 1'b0;  addr_rom[10174]='h00003b84;  wr_data_rom[10174]='h00000000;
    rd_cycle[10175] = 1'b1;  wr_cycle[10175] = 1'b0;  addr_rom[10175]='h00000bb4;  wr_data_rom[10175]='h00000000;
    rd_cycle[10176] = 1'b0;  wr_cycle[10176] = 1'b1;  addr_rom[10176]='h00003188;  wr_data_rom[10176]='h000012e3;
    rd_cycle[10177] = 1'b1;  wr_cycle[10177] = 1'b0;  addr_rom[10177]='h000016f8;  wr_data_rom[10177]='h00000000;
    rd_cycle[10178] = 1'b0;  wr_cycle[10178] = 1'b1;  addr_rom[10178]='h0000117c;  wr_data_rom[10178]='h00003bdf;
    rd_cycle[10179] = 1'b1;  wr_cycle[10179] = 1'b0;  addr_rom[10179]='h00002fc0;  wr_data_rom[10179]='h00000000;
    rd_cycle[10180] = 1'b0;  wr_cycle[10180] = 1'b1;  addr_rom[10180]='h00003be0;  wr_data_rom[10180]='h00000737;
    rd_cycle[10181] = 1'b1;  wr_cycle[10181] = 1'b0;  addr_rom[10181]='h000010c8;  wr_data_rom[10181]='h00000000;
    rd_cycle[10182] = 1'b0;  wr_cycle[10182] = 1'b1;  addr_rom[10182]='h00000314;  wr_data_rom[10182]='h000013b5;
    rd_cycle[10183] = 1'b1;  wr_cycle[10183] = 1'b0;  addr_rom[10183]='h00001458;  wr_data_rom[10183]='h00000000;
    rd_cycle[10184] = 1'b0;  wr_cycle[10184] = 1'b1;  addr_rom[10184]='h00002cb0;  wr_data_rom[10184]='h00003a74;
    rd_cycle[10185] = 1'b0;  wr_cycle[10185] = 1'b1;  addr_rom[10185]='h00000560;  wr_data_rom[10185]='h00002c7a;
    rd_cycle[10186] = 1'b1;  wr_cycle[10186] = 1'b0;  addr_rom[10186]='h00000648;  wr_data_rom[10186]='h00000000;
    rd_cycle[10187] = 1'b0;  wr_cycle[10187] = 1'b1;  addr_rom[10187]='h000008d8;  wr_data_rom[10187]='h00002855;
    rd_cycle[10188] = 1'b1;  wr_cycle[10188] = 1'b0;  addr_rom[10188]='h00001bb8;  wr_data_rom[10188]='h00000000;
    rd_cycle[10189] = 1'b1;  wr_cycle[10189] = 1'b0;  addr_rom[10189]='h00000cfc;  wr_data_rom[10189]='h00000000;
    rd_cycle[10190] = 1'b1;  wr_cycle[10190] = 1'b0;  addr_rom[10190]='h00000e48;  wr_data_rom[10190]='h00000000;
    rd_cycle[10191] = 1'b0;  wr_cycle[10191] = 1'b1;  addr_rom[10191]='h000010e4;  wr_data_rom[10191]='h00001183;
    rd_cycle[10192] = 1'b1;  wr_cycle[10192] = 1'b0;  addr_rom[10192]='h0000007c;  wr_data_rom[10192]='h00000000;
    rd_cycle[10193] = 1'b0;  wr_cycle[10193] = 1'b1;  addr_rom[10193]='h00001a04;  wr_data_rom[10193]='h000007a7;
    rd_cycle[10194] = 1'b1;  wr_cycle[10194] = 1'b0;  addr_rom[10194]='h00000f08;  wr_data_rom[10194]='h00000000;
    rd_cycle[10195] = 1'b1;  wr_cycle[10195] = 1'b0;  addr_rom[10195]='h00000734;  wr_data_rom[10195]='h00000000;
    rd_cycle[10196] = 1'b1;  wr_cycle[10196] = 1'b0;  addr_rom[10196]='h00000730;  wr_data_rom[10196]='h00000000;
    rd_cycle[10197] = 1'b1;  wr_cycle[10197] = 1'b0;  addr_rom[10197]='h00003030;  wr_data_rom[10197]='h00000000;
    rd_cycle[10198] = 1'b0;  wr_cycle[10198] = 1'b1;  addr_rom[10198]='h00002c14;  wr_data_rom[10198]='h00001b31;
    rd_cycle[10199] = 1'b1;  wr_cycle[10199] = 1'b0;  addr_rom[10199]='h000036ac;  wr_data_rom[10199]='h00000000;
    rd_cycle[10200] = 1'b1;  wr_cycle[10200] = 1'b0;  addr_rom[10200]='h000016f0;  wr_data_rom[10200]='h00000000;
    rd_cycle[10201] = 1'b1;  wr_cycle[10201] = 1'b0;  addr_rom[10201]='h0000114c;  wr_data_rom[10201]='h00000000;
    rd_cycle[10202] = 1'b0;  wr_cycle[10202] = 1'b1;  addr_rom[10202]='h000017a4;  wr_data_rom[10202]='h0000220d;
    rd_cycle[10203] = 1'b0;  wr_cycle[10203] = 1'b1;  addr_rom[10203]='h000028ac;  wr_data_rom[10203]='h00000c10;
    rd_cycle[10204] = 1'b1;  wr_cycle[10204] = 1'b0;  addr_rom[10204]='h0000135c;  wr_data_rom[10204]='h00000000;
    rd_cycle[10205] = 1'b0;  wr_cycle[10205] = 1'b1;  addr_rom[10205]='h00000eb0;  wr_data_rom[10205]='h00003d9b;
    rd_cycle[10206] = 1'b0;  wr_cycle[10206] = 1'b1;  addr_rom[10206]='h00000398;  wr_data_rom[10206]='h000025c0;
    rd_cycle[10207] = 1'b1;  wr_cycle[10207] = 1'b0;  addr_rom[10207]='h00000d78;  wr_data_rom[10207]='h00000000;
    rd_cycle[10208] = 1'b1;  wr_cycle[10208] = 1'b0;  addr_rom[10208]='h0000155c;  wr_data_rom[10208]='h00000000;
    rd_cycle[10209] = 1'b0;  wr_cycle[10209] = 1'b1;  addr_rom[10209]='h000039f4;  wr_data_rom[10209]='h00003d23;
    rd_cycle[10210] = 1'b0;  wr_cycle[10210] = 1'b1;  addr_rom[10210]='h0000140c;  wr_data_rom[10210]='h0000339d;
    rd_cycle[10211] = 1'b0;  wr_cycle[10211] = 1'b1;  addr_rom[10211]='h00000644;  wr_data_rom[10211]='h0000188b;
    rd_cycle[10212] = 1'b0;  wr_cycle[10212] = 1'b1;  addr_rom[10212]='h00001694;  wr_data_rom[10212]='h00000292;
    rd_cycle[10213] = 1'b1;  wr_cycle[10213] = 1'b0;  addr_rom[10213]='h00003360;  wr_data_rom[10213]='h00000000;
    rd_cycle[10214] = 1'b0;  wr_cycle[10214] = 1'b1;  addr_rom[10214]='h00000ea4;  wr_data_rom[10214]='h000007ab;
    rd_cycle[10215] = 1'b1;  wr_cycle[10215] = 1'b0;  addr_rom[10215]='h00001d24;  wr_data_rom[10215]='h00000000;
    rd_cycle[10216] = 1'b0;  wr_cycle[10216] = 1'b1;  addr_rom[10216]='h00002064;  wr_data_rom[10216]='h00002dd6;
    rd_cycle[10217] = 1'b0;  wr_cycle[10217] = 1'b1;  addr_rom[10217]='h00003d14;  wr_data_rom[10217]='h00000011;
    rd_cycle[10218] = 1'b1;  wr_cycle[10218] = 1'b0;  addr_rom[10218]='h00002998;  wr_data_rom[10218]='h00000000;
    rd_cycle[10219] = 1'b0;  wr_cycle[10219] = 1'b1;  addr_rom[10219]='h00002428;  wr_data_rom[10219]='h00000a05;
    rd_cycle[10220] = 1'b0;  wr_cycle[10220] = 1'b1;  addr_rom[10220]='h0000309c;  wr_data_rom[10220]='h000007a2;
    rd_cycle[10221] = 1'b1;  wr_cycle[10221] = 1'b0;  addr_rom[10221]='h00000328;  wr_data_rom[10221]='h00000000;
    rd_cycle[10222] = 1'b1;  wr_cycle[10222] = 1'b0;  addr_rom[10222]='h000013a0;  wr_data_rom[10222]='h00000000;
    rd_cycle[10223] = 1'b0;  wr_cycle[10223] = 1'b1;  addr_rom[10223]='h0000269c;  wr_data_rom[10223]='h00002f5d;
    rd_cycle[10224] = 1'b0;  wr_cycle[10224] = 1'b1;  addr_rom[10224]='h00000338;  wr_data_rom[10224]='h00001bdd;
    rd_cycle[10225] = 1'b1;  wr_cycle[10225] = 1'b0;  addr_rom[10225]='h00000bb0;  wr_data_rom[10225]='h00000000;
    rd_cycle[10226] = 1'b1;  wr_cycle[10226] = 1'b0;  addr_rom[10226]='h00001524;  wr_data_rom[10226]='h00000000;
    rd_cycle[10227] = 1'b1;  wr_cycle[10227] = 1'b0;  addr_rom[10227]='h00002c28;  wr_data_rom[10227]='h00000000;
    rd_cycle[10228] = 1'b0;  wr_cycle[10228] = 1'b1;  addr_rom[10228]='h000022c0;  wr_data_rom[10228]='h00003571;
    rd_cycle[10229] = 1'b0;  wr_cycle[10229] = 1'b1;  addr_rom[10229]='h00002188;  wr_data_rom[10229]='h000002e3;
    rd_cycle[10230] = 1'b1;  wr_cycle[10230] = 1'b0;  addr_rom[10230]='h00001458;  wr_data_rom[10230]='h00000000;
    rd_cycle[10231] = 1'b1;  wr_cycle[10231] = 1'b0;  addr_rom[10231]='h000024c4;  wr_data_rom[10231]='h00000000;
    rd_cycle[10232] = 1'b0;  wr_cycle[10232] = 1'b1;  addr_rom[10232]='h000012f0;  wr_data_rom[10232]='h00000d13;
    rd_cycle[10233] = 1'b0;  wr_cycle[10233] = 1'b1;  addr_rom[10233]='h00000aec;  wr_data_rom[10233]='h0000071f;
    rd_cycle[10234] = 1'b1;  wr_cycle[10234] = 1'b0;  addr_rom[10234]='h00002354;  wr_data_rom[10234]='h00000000;
    rd_cycle[10235] = 1'b1;  wr_cycle[10235] = 1'b0;  addr_rom[10235]='h00000b88;  wr_data_rom[10235]='h00000000;
    rd_cycle[10236] = 1'b0;  wr_cycle[10236] = 1'b1;  addr_rom[10236]='h00003bac;  wr_data_rom[10236]='h00002a0a;
    rd_cycle[10237] = 1'b0;  wr_cycle[10237] = 1'b1;  addr_rom[10237]='h00001930;  wr_data_rom[10237]='h00002aa9;
    rd_cycle[10238] = 1'b0;  wr_cycle[10238] = 1'b1;  addr_rom[10238]='h00002bf0;  wr_data_rom[10238]='h00003baa;
    rd_cycle[10239] = 1'b1;  wr_cycle[10239] = 1'b0;  addr_rom[10239]='h00003710;  wr_data_rom[10239]='h00000000;
    rd_cycle[10240] = 1'b1;  wr_cycle[10240] = 1'b0;  addr_rom[10240]='h00001ae4;  wr_data_rom[10240]='h00000000;
    rd_cycle[10241] = 1'b1;  wr_cycle[10241] = 1'b0;  addr_rom[10241]='h00000590;  wr_data_rom[10241]='h00000000;
    rd_cycle[10242] = 1'b0;  wr_cycle[10242] = 1'b1;  addr_rom[10242]='h00001184;  wr_data_rom[10242]='h00001f86;
    rd_cycle[10243] = 1'b0;  wr_cycle[10243] = 1'b1;  addr_rom[10243]='h0000132c;  wr_data_rom[10243]='h0000298e;
    rd_cycle[10244] = 1'b1;  wr_cycle[10244] = 1'b0;  addr_rom[10244]='h00002580;  wr_data_rom[10244]='h00000000;
    rd_cycle[10245] = 1'b1;  wr_cycle[10245] = 1'b0;  addr_rom[10245]='h00002ca4;  wr_data_rom[10245]='h00000000;
    rd_cycle[10246] = 1'b0;  wr_cycle[10246] = 1'b1;  addr_rom[10246]='h00001034;  wr_data_rom[10246]='h0000282f;
    rd_cycle[10247] = 1'b1;  wr_cycle[10247] = 1'b0;  addr_rom[10247]='h00001774;  wr_data_rom[10247]='h00000000;
    rd_cycle[10248] = 1'b0;  wr_cycle[10248] = 1'b1;  addr_rom[10248]='h00001ff4;  wr_data_rom[10248]='h00003e62;
    rd_cycle[10249] = 1'b0;  wr_cycle[10249] = 1'b1;  addr_rom[10249]='h000006e4;  wr_data_rom[10249]='h00003895;
    rd_cycle[10250] = 1'b0;  wr_cycle[10250] = 1'b1;  addr_rom[10250]='h000025d0;  wr_data_rom[10250]='h00003381;
    rd_cycle[10251] = 1'b1;  wr_cycle[10251] = 1'b0;  addr_rom[10251]='h000006b4;  wr_data_rom[10251]='h00000000;
    rd_cycle[10252] = 1'b0;  wr_cycle[10252] = 1'b1;  addr_rom[10252]='h00003ab4;  wr_data_rom[10252]='h00001577;
    rd_cycle[10253] = 1'b1;  wr_cycle[10253] = 1'b0;  addr_rom[10253]='h000022fc;  wr_data_rom[10253]='h00000000;
    rd_cycle[10254] = 1'b1;  wr_cycle[10254] = 1'b0;  addr_rom[10254]='h00001da0;  wr_data_rom[10254]='h00000000;
    rd_cycle[10255] = 1'b1;  wr_cycle[10255] = 1'b0;  addr_rom[10255]='h00000a2c;  wr_data_rom[10255]='h00000000;
    rd_cycle[10256] = 1'b0;  wr_cycle[10256] = 1'b1;  addr_rom[10256]='h00001028;  wr_data_rom[10256]='h00002952;
    rd_cycle[10257] = 1'b1;  wr_cycle[10257] = 1'b0;  addr_rom[10257]='h00001e6c;  wr_data_rom[10257]='h00000000;
    rd_cycle[10258] = 1'b0;  wr_cycle[10258] = 1'b1;  addr_rom[10258]='h00003fe4;  wr_data_rom[10258]='h0000295e;
    rd_cycle[10259] = 1'b0;  wr_cycle[10259] = 1'b1;  addr_rom[10259]='h00003648;  wr_data_rom[10259]='h0000265b;
    rd_cycle[10260] = 1'b0;  wr_cycle[10260] = 1'b1;  addr_rom[10260]='h00003fac;  wr_data_rom[10260]='h00001350;
    rd_cycle[10261] = 1'b1;  wr_cycle[10261] = 1'b0;  addr_rom[10261]='h00003ee8;  wr_data_rom[10261]='h00000000;
    rd_cycle[10262] = 1'b1;  wr_cycle[10262] = 1'b0;  addr_rom[10262]='h00003a3c;  wr_data_rom[10262]='h00000000;
    rd_cycle[10263] = 1'b0;  wr_cycle[10263] = 1'b1;  addr_rom[10263]='h00002f18;  wr_data_rom[10263]='h00003800;
    rd_cycle[10264] = 1'b1;  wr_cycle[10264] = 1'b0;  addr_rom[10264]='h000039a0;  wr_data_rom[10264]='h00000000;
    rd_cycle[10265] = 1'b0;  wr_cycle[10265] = 1'b1;  addr_rom[10265]='h00002d98;  wr_data_rom[10265]='h00000cb7;
    rd_cycle[10266] = 1'b0;  wr_cycle[10266] = 1'b1;  addr_rom[10266]='h000017a0;  wr_data_rom[10266]='h00001902;
    rd_cycle[10267] = 1'b1;  wr_cycle[10267] = 1'b0;  addr_rom[10267]='h00003850;  wr_data_rom[10267]='h00000000;
    rd_cycle[10268] = 1'b1;  wr_cycle[10268] = 1'b0;  addr_rom[10268]='h000001ec;  wr_data_rom[10268]='h00000000;
    rd_cycle[10269] = 1'b1;  wr_cycle[10269] = 1'b0;  addr_rom[10269]='h00002474;  wr_data_rom[10269]='h00000000;
    rd_cycle[10270] = 1'b0;  wr_cycle[10270] = 1'b1;  addr_rom[10270]='h00002a14;  wr_data_rom[10270]='h00003105;
    rd_cycle[10271] = 1'b1;  wr_cycle[10271] = 1'b0;  addr_rom[10271]='h00002d54;  wr_data_rom[10271]='h00000000;
    rd_cycle[10272] = 1'b1;  wr_cycle[10272] = 1'b0;  addr_rom[10272]='h000017b4;  wr_data_rom[10272]='h00000000;
    rd_cycle[10273] = 1'b0;  wr_cycle[10273] = 1'b1;  addr_rom[10273]='h00003550;  wr_data_rom[10273]='h00003a0b;
    rd_cycle[10274] = 1'b0;  wr_cycle[10274] = 1'b1;  addr_rom[10274]='h00002304;  wr_data_rom[10274]='h0000116f;
    rd_cycle[10275] = 1'b0;  wr_cycle[10275] = 1'b1;  addr_rom[10275]='h00000944;  wr_data_rom[10275]='h00002c1c;
    rd_cycle[10276] = 1'b0;  wr_cycle[10276] = 1'b1;  addr_rom[10276]='h00003e3c;  wr_data_rom[10276]='h000011da;
    rd_cycle[10277] = 1'b0;  wr_cycle[10277] = 1'b1;  addr_rom[10277]='h000039e8;  wr_data_rom[10277]='h00002fe3;
    rd_cycle[10278] = 1'b1;  wr_cycle[10278] = 1'b0;  addr_rom[10278]='h00002284;  wr_data_rom[10278]='h00000000;
    rd_cycle[10279] = 1'b1;  wr_cycle[10279] = 1'b0;  addr_rom[10279]='h00000b44;  wr_data_rom[10279]='h00000000;
    rd_cycle[10280] = 1'b1;  wr_cycle[10280] = 1'b0;  addr_rom[10280]='h000014e0;  wr_data_rom[10280]='h00000000;
    rd_cycle[10281] = 1'b0;  wr_cycle[10281] = 1'b1;  addr_rom[10281]='h00001e14;  wr_data_rom[10281]='h00001e93;
    rd_cycle[10282] = 1'b0;  wr_cycle[10282] = 1'b1;  addr_rom[10282]='h00000a7c;  wr_data_rom[10282]='h000006ca;
    rd_cycle[10283] = 1'b0;  wr_cycle[10283] = 1'b1;  addr_rom[10283]='h00002b80;  wr_data_rom[10283]='h00002f6b;
    rd_cycle[10284] = 1'b0;  wr_cycle[10284] = 1'b1;  addr_rom[10284]='h000025a4;  wr_data_rom[10284]='h0000054b;
    rd_cycle[10285] = 1'b0;  wr_cycle[10285] = 1'b1;  addr_rom[10285]='h0000335c;  wr_data_rom[10285]='h00002a86;
    rd_cycle[10286] = 1'b0;  wr_cycle[10286] = 1'b1;  addr_rom[10286]='h00000204;  wr_data_rom[10286]='h00002978;
    rd_cycle[10287] = 1'b1;  wr_cycle[10287] = 1'b0;  addr_rom[10287]='h00000ed0;  wr_data_rom[10287]='h00000000;
    rd_cycle[10288] = 1'b0;  wr_cycle[10288] = 1'b1;  addr_rom[10288]='h00002dc8;  wr_data_rom[10288]='h000008cb;
    rd_cycle[10289] = 1'b1;  wr_cycle[10289] = 1'b0;  addr_rom[10289]='h000013a0;  wr_data_rom[10289]='h00000000;
    rd_cycle[10290] = 1'b0;  wr_cycle[10290] = 1'b1;  addr_rom[10290]='h0000347c;  wr_data_rom[10290]='h00003e51;
    rd_cycle[10291] = 1'b0;  wr_cycle[10291] = 1'b1;  addr_rom[10291]='h00000350;  wr_data_rom[10291]='h00001416;
    rd_cycle[10292] = 1'b1;  wr_cycle[10292] = 1'b0;  addr_rom[10292]='h0000270c;  wr_data_rom[10292]='h00000000;
    rd_cycle[10293] = 1'b1;  wr_cycle[10293] = 1'b0;  addr_rom[10293]='h00002a3c;  wr_data_rom[10293]='h00000000;
    rd_cycle[10294] = 1'b1;  wr_cycle[10294] = 1'b0;  addr_rom[10294]='h00003d98;  wr_data_rom[10294]='h00000000;
    rd_cycle[10295] = 1'b0;  wr_cycle[10295] = 1'b1;  addr_rom[10295]='h00002ed4;  wr_data_rom[10295]='h00000471;
    rd_cycle[10296] = 1'b1;  wr_cycle[10296] = 1'b0;  addr_rom[10296]='h00002f04;  wr_data_rom[10296]='h00000000;
    rd_cycle[10297] = 1'b1;  wr_cycle[10297] = 1'b0;  addr_rom[10297]='h00000658;  wr_data_rom[10297]='h00000000;
    rd_cycle[10298] = 1'b0;  wr_cycle[10298] = 1'b1;  addr_rom[10298]='h00002094;  wr_data_rom[10298]='h00002071;
    rd_cycle[10299] = 1'b0;  wr_cycle[10299] = 1'b1;  addr_rom[10299]='h00003f54;  wr_data_rom[10299]='h0000140d;
    rd_cycle[10300] = 1'b1;  wr_cycle[10300] = 1'b0;  addr_rom[10300]='h00003430;  wr_data_rom[10300]='h00000000;
    rd_cycle[10301] = 1'b0;  wr_cycle[10301] = 1'b1;  addr_rom[10301]='h000020f8;  wr_data_rom[10301]='h00001c6b;
    rd_cycle[10302] = 1'b1;  wr_cycle[10302] = 1'b0;  addr_rom[10302]='h00003374;  wr_data_rom[10302]='h00000000;
    rd_cycle[10303] = 1'b1;  wr_cycle[10303] = 1'b0;  addr_rom[10303]='h00000a70;  wr_data_rom[10303]='h00000000;
    rd_cycle[10304] = 1'b0;  wr_cycle[10304] = 1'b1;  addr_rom[10304]='h000023a0;  wr_data_rom[10304]='h00003a99;
    rd_cycle[10305] = 1'b0;  wr_cycle[10305] = 1'b1;  addr_rom[10305]='h000027d0;  wr_data_rom[10305]='h00003eff;
    rd_cycle[10306] = 1'b1;  wr_cycle[10306] = 1'b0;  addr_rom[10306]='h000030d0;  wr_data_rom[10306]='h00000000;
    rd_cycle[10307] = 1'b0;  wr_cycle[10307] = 1'b1;  addr_rom[10307]='h00001660;  wr_data_rom[10307]='h00003cd6;
    rd_cycle[10308] = 1'b1;  wr_cycle[10308] = 1'b0;  addr_rom[10308]='h00003174;  wr_data_rom[10308]='h00000000;
    rd_cycle[10309] = 1'b1;  wr_cycle[10309] = 1'b0;  addr_rom[10309]='h000023b0;  wr_data_rom[10309]='h00000000;
    rd_cycle[10310] = 1'b0;  wr_cycle[10310] = 1'b1;  addr_rom[10310]='h00002380;  wr_data_rom[10310]='h00001254;
    rd_cycle[10311] = 1'b0;  wr_cycle[10311] = 1'b1;  addr_rom[10311]='h00000860;  wr_data_rom[10311]='h000032bc;
    rd_cycle[10312] = 1'b1;  wr_cycle[10312] = 1'b0;  addr_rom[10312]='h00000a90;  wr_data_rom[10312]='h00000000;
    rd_cycle[10313] = 1'b0;  wr_cycle[10313] = 1'b1;  addr_rom[10313]='h00000714;  wr_data_rom[10313]='h0000109d;
    rd_cycle[10314] = 1'b1;  wr_cycle[10314] = 1'b0;  addr_rom[10314]='h00003464;  wr_data_rom[10314]='h00000000;
    rd_cycle[10315] = 1'b1;  wr_cycle[10315] = 1'b0;  addr_rom[10315]='h000036b8;  wr_data_rom[10315]='h00000000;
    rd_cycle[10316] = 1'b0;  wr_cycle[10316] = 1'b1;  addr_rom[10316]='h000009e8;  wr_data_rom[10316]='h00002cfe;
    rd_cycle[10317] = 1'b1;  wr_cycle[10317] = 1'b0;  addr_rom[10317]='h0000265c;  wr_data_rom[10317]='h00000000;
    rd_cycle[10318] = 1'b1;  wr_cycle[10318] = 1'b0;  addr_rom[10318]='h00003190;  wr_data_rom[10318]='h00000000;
    rd_cycle[10319] = 1'b0;  wr_cycle[10319] = 1'b1;  addr_rom[10319]='h000025dc;  wr_data_rom[10319]='h00002b6b;
    rd_cycle[10320] = 1'b1;  wr_cycle[10320] = 1'b0;  addr_rom[10320]='h00002d98;  wr_data_rom[10320]='h00000000;
    rd_cycle[10321] = 1'b1;  wr_cycle[10321] = 1'b0;  addr_rom[10321]='h00000774;  wr_data_rom[10321]='h00000000;
    rd_cycle[10322] = 1'b1;  wr_cycle[10322] = 1'b0;  addr_rom[10322]='h00000f18;  wr_data_rom[10322]='h00000000;
    rd_cycle[10323] = 1'b1;  wr_cycle[10323] = 1'b0;  addr_rom[10323]='h00000c1c;  wr_data_rom[10323]='h00000000;
    rd_cycle[10324] = 1'b0;  wr_cycle[10324] = 1'b1;  addr_rom[10324]='h00000360;  wr_data_rom[10324]='h0000141e;
    rd_cycle[10325] = 1'b0;  wr_cycle[10325] = 1'b1;  addr_rom[10325]='h00003624;  wr_data_rom[10325]='h0000024f;
    rd_cycle[10326] = 1'b0;  wr_cycle[10326] = 1'b1;  addr_rom[10326]='h00003574;  wr_data_rom[10326]='h00001086;
    rd_cycle[10327] = 1'b1;  wr_cycle[10327] = 1'b0;  addr_rom[10327]='h00002140;  wr_data_rom[10327]='h00000000;
    rd_cycle[10328] = 1'b1;  wr_cycle[10328] = 1'b0;  addr_rom[10328]='h00000068;  wr_data_rom[10328]='h00000000;
    rd_cycle[10329] = 1'b1;  wr_cycle[10329] = 1'b0;  addr_rom[10329]='h0000303c;  wr_data_rom[10329]='h00000000;
    rd_cycle[10330] = 1'b0;  wr_cycle[10330] = 1'b1;  addr_rom[10330]='h0000114c;  wr_data_rom[10330]='h000029e4;
    rd_cycle[10331] = 1'b1;  wr_cycle[10331] = 1'b0;  addr_rom[10331]='h00000b24;  wr_data_rom[10331]='h00000000;
    rd_cycle[10332] = 1'b0;  wr_cycle[10332] = 1'b1;  addr_rom[10332]='h000019e4;  wr_data_rom[10332]='h00003298;
    rd_cycle[10333] = 1'b1;  wr_cycle[10333] = 1'b0;  addr_rom[10333]='h000034f4;  wr_data_rom[10333]='h00000000;
    rd_cycle[10334] = 1'b1;  wr_cycle[10334] = 1'b0;  addr_rom[10334]='h00000898;  wr_data_rom[10334]='h00000000;
    rd_cycle[10335] = 1'b0;  wr_cycle[10335] = 1'b1;  addr_rom[10335]='h0000257c;  wr_data_rom[10335]='h00000aa9;
    rd_cycle[10336] = 1'b1;  wr_cycle[10336] = 1'b0;  addr_rom[10336]='h00001dd8;  wr_data_rom[10336]='h00000000;
    rd_cycle[10337] = 1'b1;  wr_cycle[10337] = 1'b0;  addr_rom[10337]='h00001efc;  wr_data_rom[10337]='h00000000;
    rd_cycle[10338] = 1'b0;  wr_cycle[10338] = 1'b1;  addr_rom[10338]='h0000028c;  wr_data_rom[10338]='h00001a4a;
    rd_cycle[10339] = 1'b0;  wr_cycle[10339] = 1'b1;  addr_rom[10339]='h000021ec;  wr_data_rom[10339]='h00003fbe;
    rd_cycle[10340] = 1'b1;  wr_cycle[10340] = 1'b0;  addr_rom[10340]='h00001398;  wr_data_rom[10340]='h00000000;
    rd_cycle[10341] = 1'b1;  wr_cycle[10341] = 1'b0;  addr_rom[10341]='h00002598;  wr_data_rom[10341]='h00000000;
    rd_cycle[10342] = 1'b1;  wr_cycle[10342] = 1'b0;  addr_rom[10342]='h00002d64;  wr_data_rom[10342]='h00000000;
    rd_cycle[10343] = 1'b0;  wr_cycle[10343] = 1'b1;  addr_rom[10343]='h00001648;  wr_data_rom[10343]='h000013bf;
    rd_cycle[10344] = 1'b1;  wr_cycle[10344] = 1'b0;  addr_rom[10344]='h00003800;  wr_data_rom[10344]='h00000000;
    rd_cycle[10345] = 1'b1;  wr_cycle[10345] = 1'b0;  addr_rom[10345]='h000032b4;  wr_data_rom[10345]='h00000000;
    rd_cycle[10346] = 1'b1;  wr_cycle[10346] = 1'b0;  addr_rom[10346]='h00001118;  wr_data_rom[10346]='h00000000;
    rd_cycle[10347] = 1'b1;  wr_cycle[10347] = 1'b0;  addr_rom[10347]='h00003988;  wr_data_rom[10347]='h00000000;
    rd_cycle[10348] = 1'b1;  wr_cycle[10348] = 1'b0;  addr_rom[10348]='h000027d0;  wr_data_rom[10348]='h00000000;
    rd_cycle[10349] = 1'b0;  wr_cycle[10349] = 1'b1;  addr_rom[10349]='h0000164c;  wr_data_rom[10349]='h00003685;
    rd_cycle[10350] = 1'b0;  wr_cycle[10350] = 1'b1;  addr_rom[10350]='h00001f6c;  wr_data_rom[10350]='h00003961;
    rd_cycle[10351] = 1'b0;  wr_cycle[10351] = 1'b1;  addr_rom[10351]='h00003988;  wr_data_rom[10351]='h00001381;
    rd_cycle[10352] = 1'b0;  wr_cycle[10352] = 1'b1;  addr_rom[10352]='h00002724;  wr_data_rom[10352]='h00002bb9;
    rd_cycle[10353] = 1'b1;  wr_cycle[10353] = 1'b0;  addr_rom[10353]='h000023e4;  wr_data_rom[10353]='h00000000;
    rd_cycle[10354] = 1'b1;  wr_cycle[10354] = 1'b0;  addr_rom[10354]='h00000728;  wr_data_rom[10354]='h00000000;
    rd_cycle[10355] = 1'b0;  wr_cycle[10355] = 1'b1;  addr_rom[10355]='h000037b8;  wr_data_rom[10355]='h00002433;
    rd_cycle[10356] = 1'b0;  wr_cycle[10356] = 1'b1;  addr_rom[10356]='h00001080;  wr_data_rom[10356]='h00003f60;
    rd_cycle[10357] = 1'b1;  wr_cycle[10357] = 1'b0;  addr_rom[10357]='h00001bc4;  wr_data_rom[10357]='h00000000;
    rd_cycle[10358] = 1'b0;  wr_cycle[10358] = 1'b1;  addr_rom[10358]='h000012cc;  wr_data_rom[10358]='h00001135;
    rd_cycle[10359] = 1'b1;  wr_cycle[10359] = 1'b0;  addr_rom[10359]='h00000620;  wr_data_rom[10359]='h00000000;
    rd_cycle[10360] = 1'b1;  wr_cycle[10360] = 1'b0;  addr_rom[10360]='h00002de4;  wr_data_rom[10360]='h00000000;
    rd_cycle[10361] = 1'b1;  wr_cycle[10361] = 1'b0;  addr_rom[10361]='h00001228;  wr_data_rom[10361]='h00000000;
    rd_cycle[10362] = 1'b1;  wr_cycle[10362] = 1'b0;  addr_rom[10362]='h000004fc;  wr_data_rom[10362]='h00000000;
    rd_cycle[10363] = 1'b1;  wr_cycle[10363] = 1'b0;  addr_rom[10363]='h0000272c;  wr_data_rom[10363]='h00000000;
    rd_cycle[10364] = 1'b1;  wr_cycle[10364] = 1'b0;  addr_rom[10364]='h0000322c;  wr_data_rom[10364]='h00000000;
    rd_cycle[10365] = 1'b1;  wr_cycle[10365] = 1'b0;  addr_rom[10365]='h0000119c;  wr_data_rom[10365]='h00000000;
    rd_cycle[10366] = 1'b1;  wr_cycle[10366] = 1'b0;  addr_rom[10366]='h00000cf0;  wr_data_rom[10366]='h00000000;
    rd_cycle[10367] = 1'b0;  wr_cycle[10367] = 1'b1;  addr_rom[10367]='h00000dcc;  wr_data_rom[10367]='h00000327;
    rd_cycle[10368] = 1'b0;  wr_cycle[10368] = 1'b1;  addr_rom[10368]='h000028fc;  wr_data_rom[10368]='h00002186;
    rd_cycle[10369] = 1'b0;  wr_cycle[10369] = 1'b1;  addr_rom[10369]='h0000281c;  wr_data_rom[10369]='h000006e4;
    rd_cycle[10370] = 1'b1;  wr_cycle[10370] = 1'b0;  addr_rom[10370]='h00002b2c;  wr_data_rom[10370]='h00000000;
    rd_cycle[10371] = 1'b1;  wr_cycle[10371] = 1'b0;  addr_rom[10371]='h000023e8;  wr_data_rom[10371]='h00000000;
    rd_cycle[10372] = 1'b1;  wr_cycle[10372] = 1'b0;  addr_rom[10372]='h00003234;  wr_data_rom[10372]='h00000000;
    rd_cycle[10373] = 1'b1;  wr_cycle[10373] = 1'b0;  addr_rom[10373]='h00002a48;  wr_data_rom[10373]='h00000000;
    rd_cycle[10374] = 1'b0;  wr_cycle[10374] = 1'b1;  addr_rom[10374]='h000010e0;  wr_data_rom[10374]='h000018e0;
    rd_cycle[10375] = 1'b0;  wr_cycle[10375] = 1'b1;  addr_rom[10375]='h00001678;  wr_data_rom[10375]='h00002368;
    rd_cycle[10376] = 1'b0;  wr_cycle[10376] = 1'b1;  addr_rom[10376]='h00001fa0;  wr_data_rom[10376]='h00000648;
    rd_cycle[10377] = 1'b0;  wr_cycle[10377] = 1'b1;  addr_rom[10377]='h00000c28;  wr_data_rom[10377]='h0000071c;
    rd_cycle[10378] = 1'b0;  wr_cycle[10378] = 1'b1;  addr_rom[10378]='h00001a64;  wr_data_rom[10378]='h00001ff6;
    rd_cycle[10379] = 1'b0;  wr_cycle[10379] = 1'b1;  addr_rom[10379]='h000017e8;  wr_data_rom[10379]='h00001c31;
    rd_cycle[10380] = 1'b1;  wr_cycle[10380] = 1'b0;  addr_rom[10380]='h00003728;  wr_data_rom[10380]='h00000000;
    rd_cycle[10381] = 1'b1;  wr_cycle[10381] = 1'b0;  addr_rom[10381]='h000007c4;  wr_data_rom[10381]='h00000000;
    rd_cycle[10382] = 1'b0;  wr_cycle[10382] = 1'b1;  addr_rom[10382]='h00001db0;  wr_data_rom[10382]='h000036c9;
    rd_cycle[10383] = 1'b0;  wr_cycle[10383] = 1'b1;  addr_rom[10383]='h00000468;  wr_data_rom[10383]='h00000858;
    rd_cycle[10384] = 1'b0;  wr_cycle[10384] = 1'b1;  addr_rom[10384]='h00001808;  wr_data_rom[10384]='h00003cd4;
    rd_cycle[10385] = 1'b1;  wr_cycle[10385] = 1'b0;  addr_rom[10385]='h00003088;  wr_data_rom[10385]='h00000000;
    rd_cycle[10386] = 1'b1;  wr_cycle[10386] = 1'b0;  addr_rom[10386]='h00000e20;  wr_data_rom[10386]='h00000000;
    rd_cycle[10387] = 1'b0;  wr_cycle[10387] = 1'b1;  addr_rom[10387]='h00001624;  wr_data_rom[10387]='h00003d7d;
    rd_cycle[10388] = 1'b1;  wr_cycle[10388] = 1'b0;  addr_rom[10388]='h00002940;  wr_data_rom[10388]='h00000000;
    rd_cycle[10389] = 1'b0;  wr_cycle[10389] = 1'b1;  addr_rom[10389]='h00002800;  wr_data_rom[10389]='h0000097d;
    rd_cycle[10390] = 1'b0;  wr_cycle[10390] = 1'b1;  addr_rom[10390]='h000025b8;  wr_data_rom[10390]='h000011e4;
    rd_cycle[10391] = 1'b1;  wr_cycle[10391] = 1'b0;  addr_rom[10391]='h00001b4c;  wr_data_rom[10391]='h00000000;
    rd_cycle[10392] = 1'b0;  wr_cycle[10392] = 1'b1;  addr_rom[10392]='h00002124;  wr_data_rom[10392]='h00001bb5;
    rd_cycle[10393] = 1'b0;  wr_cycle[10393] = 1'b1;  addr_rom[10393]='h00002598;  wr_data_rom[10393]='h00003d5a;
    rd_cycle[10394] = 1'b0;  wr_cycle[10394] = 1'b1;  addr_rom[10394]='h000009b0;  wr_data_rom[10394]='h00002f21;
    rd_cycle[10395] = 1'b0;  wr_cycle[10395] = 1'b1;  addr_rom[10395]='h00000010;  wr_data_rom[10395]='h00003c33;
    rd_cycle[10396] = 1'b1;  wr_cycle[10396] = 1'b0;  addr_rom[10396]='h0000036c;  wr_data_rom[10396]='h00000000;
    rd_cycle[10397] = 1'b1;  wr_cycle[10397] = 1'b0;  addr_rom[10397]='h00001510;  wr_data_rom[10397]='h00000000;
    rd_cycle[10398] = 1'b1;  wr_cycle[10398] = 1'b0;  addr_rom[10398]='h00001e44;  wr_data_rom[10398]='h00000000;
    rd_cycle[10399] = 1'b0;  wr_cycle[10399] = 1'b1;  addr_rom[10399]='h00002fcc;  wr_data_rom[10399]='h00002aa5;
    rd_cycle[10400] = 1'b1;  wr_cycle[10400] = 1'b0;  addr_rom[10400]='h00000e54;  wr_data_rom[10400]='h00000000;
    rd_cycle[10401] = 1'b0;  wr_cycle[10401] = 1'b1;  addr_rom[10401]='h000036f8;  wr_data_rom[10401]='h000032fd;
    rd_cycle[10402] = 1'b0;  wr_cycle[10402] = 1'b1;  addr_rom[10402]='h00000598;  wr_data_rom[10402]='h000033e4;
    rd_cycle[10403] = 1'b0;  wr_cycle[10403] = 1'b1;  addr_rom[10403]='h000037ec;  wr_data_rom[10403]='h000017ea;
    rd_cycle[10404] = 1'b1;  wr_cycle[10404] = 1'b0;  addr_rom[10404]='h000011c0;  wr_data_rom[10404]='h00000000;
    rd_cycle[10405] = 1'b0;  wr_cycle[10405] = 1'b1;  addr_rom[10405]='h000006d0;  wr_data_rom[10405]='h00003166;
    rd_cycle[10406] = 1'b0;  wr_cycle[10406] = 1'b1;  addr_rom[10406]='h000007dc;  wr_data_rom[10406]='h00003b15;
    rd_cycle[10407] = 1'b0;  wr_cycle[10407] = 1'b1;  addr_rom[10407]='h000021c4;  wr_data_rom[10407]='h00000ba9;
    rd_cycle[10408] = 1'b0;  wr_cycle[10408] = 1'b1;  addr_rom[10408]='h000039a0;  wr_data_rom[10408]='h000023c7;
    rd_cycle[10409] = 1'b0;  wr_cycle[10409] = 1'b1;  addr_rom[10409]='h000019e4;  wr_data_rom[10409]='h000019ac;
    rd_cycle[10410] = 1'b1;  wr_cycle[10410] = 1'b0;  addr_rom[10410]='h0000346c;  wr_data_rom[10410]='h00000000;
    rd_cycle[10411] = 1'b0;  wr_cycle[10411] = 1'b1;  addr_rom[10411]='h00001cbc;  wr_data_rom[10411]='h00000b54;
    rd_cycle[10412] = 1'b0;  wr_cycle[10412] = 1'b1;  addr_rom[10412]='h0000275c;  wr_data_rom[10412]='h00001f2d;
    rd_cycle[10413] = 1'b0;  wr_cycle[10413] = 1'b1;  addr_rom[10413]='h00001da8;  wr_data_rom[10413]='h00000234;
    rd_cycle[10414] = 1'b1;  wr_cycle[10414] = 1'b0;  addr_rom[10414]='h00003fa8;  wr_data_rom[10414]='h00000000;
    rd_cycle[10415] = 1'b1;  wr_cycle[10415] = 1'b0;  addr_rom[10415]='h00001d2c;  wr_data_rom[10415]='h00000000;
    rd_cycle[10416] = 1'b0;  wr_cycle[10416] = 1'b1;  addr_rom[10416]='h00003c74;  wr_data_rom[10416]='h0000113d;
    rd_cycle[10417] = 1'b0;  wr_cycle[10417] = 1'b1;  addr_rom[10417]='h000001a8;  wr_data_rom[10417]='h00001f10;
    rd_cycle[10418] = 1'b1;  wr_cycle[10418] = 1'b0;  addr_rom[10418]='h000008d8;  wr_data_rom[10418]='h00000000;
    rd_cycle[10419] = 1'b0;  wr_cycle[10419] = 1'b1;  addr_rom[10419]='h000018fc;  wr_data_rom[10419]='h0000024f;
    rd_cycle[10420] = 1'b0;  wr_cycle[10420] = 1'b1;  addr_rom[10420]='h00001010;  wr_data_rom[10420]='h000013ff;
    rd_cycle[10421] = 1'b1;  wr_cycle[10421] = 1'b0;  addr_rom[10421]='h00000f5c;  wr_data_rom[10421]='h00000000;
    rd_cycle[10422] = 1'b1;  wr_cycle[10422] = 1'b0;  addr_rom[10422]='h00002294;  wr_data_rom[10422]='h00000000;
    rd_cycle[10423] = 1'b1;  wr_cycle[10423] = 1'b0;  addr_rom[10423]='h00000d84;  wr_data_rom[10423]='h00000000;
    rd_cycle[10424] = 1'b1;  wr_cycle[10424] = 1'b0;  addr_rom[10424]='h00000c40;  wr_data_rom[10424]='h00000000;
    rd_cycle[10425] = 1'b1;  wr_cycle[10425] = 1'b0;  addr_rom[10425]='h000007fc;  wr_data_rom[10425]='h00000000;
    rd_cycle[10426] = 1'b1;  wr_cycle[10426] = 1'b0;  addr_rom[10426]='h00000d54;  wr_data_rom[10426]='h00000000;
    rd_cycle[10427] = 1'b0;  wr_cycle[10427] = 1'b1;  addr_rom[10427]='h00001e24;  wr_data_rom[10427]='h00000e02;
    rd_cycle[10428] = 1'b1;  wr_cycle[10428] = 1'b0;  addr_rom[10428]='h000010a4;  wr_data_rom[10428]='h00000000;
    rd_cycle[10429] = 1'b0;  wr_cycle[10429] = 1'b1;  addr_rom[10429]='h00000a40;  wr_data_rom[10429]='h000005dc;
    rd_cycle[10430] = 1'b1;  wr_cycle[10430] = 1'b0;  addr_rom[10430]='h00001978;  wr_data_rom[10430]='h00000000;
    rd_cycle[10431] = 1'b0;  wr_cycle[10431] = 1'b1;  addr_rom[10431]='h00000fd8;  wr_data_rom[10431]='h00002f3e;
    rd_cycle[10432] = 1'b0;  wr_cycle[10432] = 1'b1;  addr_rom[10432]='h00001888;  wr_data_rom[10432]='h0000088d;
    rd_cycle[10433] = 1'b1;  wr_cycle[10433] = 1'b0;  addr_rom[10433]='h0000239c;  wr_data_rom[10433]='h00000000;
    rd_cycle[10434] = 1'b1;  wr_cycle[10434] = 1'b0;  addr_rom[10434]='h00002b54;  wr_data_rom[10434]='h00000000;
    rd_cycle[10435] = 1'b0;  wr_cycle[10435] = 1'b1;  addr_rom[10435]='h0000045c;  wr_data_rom[10435]='h00002654;
    rd_cycle[10436] = 1'b1;  wr_cycle[10436] = 1'b0;  addr_rom[10436]='h00002860;  wr_data_rom[10436]='h00000000;
    rd_cycle[10437] = 1'b0;  wr_cycle[10437] = 1'b1;  addr_rom[10437]='h0000388c;  wr_data_rom[10437]='h00001042;
    rd_cycle[10438] = 1'b0;  wr_cycle[10438] = 1'b1;  addr_rom[10438]='h00002774;  wr_data_rom[10438]='h00002e1f;
    rd_cycle[10439] = 1'b0;  wr_cycle[10439] = 1'b1;  addr_rom[10439]='h00003324;  wr_data_rom[10439]='h00000eac;
    rd_cycle[10440] = 1'b0;  wr_cycle[10440] = 1'b1;  addr_rom[10440]='h00001f94;  wr_data_rom[10440]='h0000138e;
    rd_cycle[10441] = 1'b0;  wr_cycle[10441] = 1'b1;  addr_rom[10441]='h00002690;  wr_data_rom[10441]='h0000318d;
    rd_cycle[10442] = 1'b1;  wr_cycle[10442] = 1'b0;  addr_rom[10442]='h000033a8;  wr_data_rom[10442]='h00000000;
    rd_cycle[10443] = 1'b0;  wr_cycle[10443] = 1'b1;  addr_rom[10443]='h00001900;  wr_data_rom[10443]='h000031af;
    rd_cycle[10444] = 1'b0;  wr_cycle[10444] = 1'b1;  addr_rom[10444]='h00003a00;  wr_data_rom[10444]='h00002675;
    rd_cycle[10445] = 1'b0;  wr_cycle[10445] = 1'b1;  addr_rom[10445]='h00002728;  wr_data_rom[10445]='h00003afc;
    rd_cycle[10446] = 1'b1;  wr_cycle[10446] = 1'b0;  addr_rom[10446]='h00003028;  wr_data_rom[10446]='h00000000;
    rd_cycle[10447] = 1'b0;  wr_cycle[10447] = 1'b1;  addr_rom[10447]='h000034bc;  wr_data_rom[10447]='h00003b9c;
    rd_cycle[10448] = 1'b0;  wr_cycle[10448] = 1'b1;  addr_rom[10448]='h000032e0;  wr_data_rom[10448]='h0000336a;
    rd_cycle[10449] = 1'b0;  wr_cycle[10449] = 1'b1;  addr_rom[10449]='h00001bd8;  wr_data_rom[10449]='h000015de;
    rd_cycle[10450] = 1'b0;  wr_cycle[10450] = 1'b1;  addr_rom[10450]='h00003da8;  wr_data_rom[10450]='h00000136;
    rd_cycle[10451] = 1'b0;  wr_cycle[10451] = 1'b1;  addr_rom[10451]='h0000395c;  wr_data_rom[10451]='h000021c7;
    rd_cycle[10452] = 1'b0;  wr_cycle[10452] = 1'b1;  addr_rom[10452]='h00001390;  wr_data_rom[10452]='h000017e2;
    rd_cycle[10453] = 1'b0;  wr_cycle[10453] = 1'b1;  addr_rom[10453]='h000018f4;  wr_data_rom[10453]='h000030f8;
    rd_cycle[10454] = 1'b1;  wr_cycle[10454] = 1'b0;  addr_rom[10454]='h00003be0;  wr_data_rom[10454]='h00000000;
    rd_cycle[10455] = 1'b1;  wr_cycle[10455] = 1'b0;  addr_rom[10455]='h000028c8;  wr_data_rom[10455]='h00000000;
    rd_cycle[10456] = 1'b1;  wr_cycle[10456] = 1'b0;  addr_rom[10456]='h00000234;  wr_data_rom[10456]='h00000000;
    rd_cycle[10457] = 1'b1;  wr_cycle[10457] = 1'b0;  addr_rom[10457]='h00001f9c;  wr_data_rom[10457]='h00000000;
    rd_cycle[10458] = 1'b0;  wr_cycle[10458] = 1'b1;  addr_rom[10458]='h00002560;  wr_data_rom[10458]='h00003188;
    rd_cycle[10459] = 1'b1;  wr_cycle[10459] = 1'b0;  addr_rom[10459]='h000013b8;  wr_data_rom[10459]='h00000000;
    rd_cycle[10460] = 1'b1;  wr_cycle[10460] = 1'b0;  addr_rom[10460]='h000004ec;  wr_data_rom[10460]='h00000000;
    rd_cycle[10461] = 1'b0;  wr_cycle[10461] = 1'b1;  addr_rom[10461]='h00000644;  wr_data_rom[10461]='h000037fb;
    rd_cycle[10462] = 1'b0;  wr_cycle[10462] = 1'b1;  addr_rom[10462]='h00001258;  wr_data_rom[10462]='h000029c0;
    rd_cycle[10463] = 1'b1;  wr_cycle[10463] = 1'b0;  addr_rom[10463]='h000030c0;  wr_data_rom[10463]='h00000000;
    rd_cycle[10464] = 1'b1;  wr_cycle[10464] = 1'b0;  addr_rom[10464]='h0000046c;  wr_data_rom[10464]='h00000000;
    rd_cycle[10465] = 1'b0;  wr_cycle[10465] = 1'b1;  addr_rom[10465]='h000012f0;  wr_data_rom[10465]='h00000e85;
    rd_cycle[10466] = 1'b1;  wr_cycle[10466] = 1'b0;  addr_rom[10466]='h000036d4;  wr_data_rom[10466]='h00000000;
    rd_cycle[10467] = 1'b1;  wr_cycle[10467] = 1'b0;  addr_rom[10467]='h00003ddc;  wr_data_rom[10467]='h00000000;
    rd_cycle[10468] = 1'b0;  wr_cycle[10468] = 1'b1;  addr_rom[10468]='h000016f8;  wr_data_rom[10468]='h00001c3a;
    rd_cycle[10469] = 1'b0;  wr_cycle[10469] = 1'b1;  addr_rom[10469]='h00002d50;  wr_data_rom[10469]='h00001a22;
    rd_cycle[10470] = 1'b0;  wr_cycle[10470] = 1'b1;  addr_rom[10470]='h0000017c;  wr_data_rom[10470]='h000013bc;
    rd_cycle[10471] = 1'b1;  wr_cycle[10471] = 1'b0;  addr_rom[10471]='h000027dc;  wr_data_rom[10471]='h00000000;
    rd_cycle[10472] = 1'b0;  wr_cycle[10472] = 1'b1;  addr_rom[10472]='h00001e68;  wr_data_rom[10472]='h000005aa;
    rd_cycle[10473] = 1'b1;  wr_cycle[10473] = 1'b0;  addr_rom[10473]='h00003644;  wr_data_rom[10473]='h00000000;
    rd_cycle[10474] = 1'b0;  wr_cycle[10474] = 1'b1;  addr_rom[10474]='h00001628;  wr_data_rom[10474]='h00002aa9;
    rd_cycle[10475] = 1'b1;  wr_cycle[10475] = 1'b0;  addr_rom[10475]='h000035b8;  wr_data_rom[10475]='h00000000;
    rd_cycle[10476] = 1'b0;  wr_cycle[10476] = 1'b1;  addr_rom[10476]='h00000c04;  wr_data_rom[10476]='h00002055;
    rd_cycle[10477] = 1'b0;  wr_cycle[10477] = 1'b1;  addr_rom[10477]='h000024a0;  wr_data_rom[10477]='h0000217e;
    rd_cycle[10478] = 1'b0;  wr_cycle[10478] = 1'b1;  addr_rom[10478]='h000016d8;  wr_data_rom[10478]='h00002f86;
    rd_cycle[10479] = 1'b1;  wr_cycle[10479] = 1'b0;  addr_rom[10479]='h00003c0c;  wr_data_rom[10479]='h00000000;
    rd_cycle[10480] = 1'b0;  wr_cycle[10480] = 1'b1;  addr_rom[10480]='h00003120;  wr_data_rom[10480]='h00001ce9;
    rd_cycle[10481] = 1'b1;  wr_cycle[10481] = 1'b0;  addr_rom[10481]='h000037b4;  wr_data_rom[10481]='h00000000;
    rd_cycle[10482] = 1'b1;  wr_cycle[10482] = 1'b0;  addr_rom[10482]='h00003484;  wr_data_rom[10482]='h00000000;
    rd_cycle[10483] = 1'b1;  wr_cycle[10483] = 1'b0;  addr_rom[10483]='h00002b70;  wr_data_rom[10483]='h00000000;
    rd_cycle[10484] = 1'b1;  wr_cycle[10484] = 1'b0;  addr_rom[10484]='h00003a78;  wr_data_rom[10484]='h00000000;
    rd_cycle[10485] = 1'b0;  wr_cycle[10485] = 1'b1;  addr_rom[10485]='h00000210;  wr_data_rom[10485]='h00001358;
    rd_cycle[10486] = 1'b1;  wr_cycle[10486] = 1'b0;  addr_rom[10486]='h0000094c;  wr_data_rom[10486]='h00000000;
    rd_cycle[10487] = 1'b0;  wr_cycle[10487] = 1'b1;  addr_rom[10487]='h000013d4;  wr_data_rom[10487]='h000022ec;
    rd_cycle[10488] = 1'b0;  wr_cycle[10488] = 1'b1;  addr_rom[10488]='h00003d28;  wr_data_rom[10488]='h0000296d;
    rd_cycle[10489] = 1'b1;  wr_cycle[10489] = 1'b0;  addr_rom[10489]='h00001820;  wr_data_rom[10489]='h00000000;
    rd_cycle[10490] = 1'b1;  wr_cycle[10490] = 1'b0;  addr_rom[10490]='h000001b4;  wr_data_rom[10490]='h00000000;
    rd_cycle[10491] = 1'b0;  wr_cycle[10491] = 1'b1;  addr_rom[10491]='h000028a4;  wr_data_rom[10491]='h00001e18;
    rd_cycle[10492] = 1'b1;  wr_cycle[10492] = 1'b0;  addr_rom[10492]='h0000054c;  wr_data_rom[10492]='h00000000;
    rd_cycle[10493] = 1'b0;  wr_cycle[10493] = 1'b1;  addr_rom[10493]='h000000fc;  wr_data_rom[10493]='h00003819;
    rd_cycle[10494] = 1'b0;  wr_cycle[10494] = 1'b1;  addr_rom[10494]='h00000770;  wr_data_rom[10494]='h000024eb;
    rd_cycle[10495] = 1'b1;  wr_cycle[10495] = 1'b0;  addr_rom[10495]='h00003e60;  wr_data_rom[10495]='h00000000;
    rd_cycle[10496] = 1'b0;  wr_cycle[10496] = 1'b1;  addr_rom[10496]='h0000388c;  wr_data_rom[10496]='h0000154d;
    rd_cycle[10497] = 1'b0;  wr_cycle[10497] = 1'b1;  addr_rom[10497]='h00002c24;  wr_data_rom[10497]='h00003ef7;
    rd_cycle[10498] = 1'b1;  wr_cycle[10498] = 1'b0;  addr_rom[10498]='h00001f8c;  wr_data_rom[10498]='h00000000;
    rd_cycle[10499] = 1'b1;  wr_cycle[10499] = 1'b0;  addr_rom[10499]='h000005ec;  wr_data_rom[10499]='h00000000;
    rd_cycle[10500] = 1'b0;  wr_cycle[10500] = 1'b1;  addr_rom[10500]='h00000270;  wr_data_rom[10500]='h000013d7;
    rd_cycle[10501] = 1'b1;  wr_cycle[10501] = 1'b0;  addr_rom[10501]='h00002a7c;  wr_data_rom[10501]='h00000000;
    rd_cycle[10502] = 1'b1;  wr_cycle[10502] = 1'b0;  addr_rom[10502]='h000005cc;  wr_data_rom[10502]='h00000000;
    rd_cycle[10503] = 1'b0;  wr_cycle[10503] = 1'b1;  addr_rom[10503]='h000027f8;  wr_data_rom[10503]='h00003c8b;
    rd_cycle[10504] = 1'b0;  wr_cycle[10504] = 1'b1;  addr_rom[10504]='h00002b20;  wr_data_rom[10504]='h00003aa6;
    rd_cycle[10505] = 1'b1;  wr_cycle[10505] = 1'b0;  addr_rom[10505]='h00003844;  wr_data_rom[10505]='h00000000;
    rd_cycle[10506] = 1'b0;  wr_cycle[10506] = 1'b1;  addr_rom[10506]='h0000159c;  wr_data_rom[10506]='h00000175;
    rd_cycle[10507] = 1'b1;  wr_cycle[10507] = 1'b0;  addr_rom[10507]='h00003a38;  wr_data_rom[10507]='h00000000;
    rd_cycle[10508] = 1'b1;  wr_cycle[10508] = 1'b0;  addr_rom[10508]='h00000ea8;  wr_data_rom[10508]='h00000000;
    rd_cycle[10509] = 1'b0;  wr_cycle[10509] = 1'b1;  addr_rom[10509]='h0000304c;  wr_data_rom[10509]='h00003225;
    rd_cycle[10510] = 1'b1;  wr_cycle[10510] = 1'b0;  addr_rom[10510]='h0000137c;  wr_data_rom[10510]='h00000000;
    rd_cycle[10511] = 1'b0;  wr_cycle[10511] = 1'b1;  addr_rom[10511]='h0000132c;  wr_data_rom[10511]='h00002533;
    rd_cycle[10512] = 1'b1;  wr_cycle[10512] = 1'b0;  addr_rom[10512]='h000026c0;  wr_data_rom[10512]='h00000000;
    rd_cycle[10513] = 1'b0;  wr_cycle[10513] = 1'b1;  addr_rom[10513]='h000014a0;  wr_data_rom[10513]='h00003abc;
    rd_cycle[10514] = 1'b1;  wr_cycle[10514] = 1'b0;  addr_rom[10514]='h00003054;  wr_data_rom[10514]='h00000000;
    rd_cycle[10515] = 1'b0;  wr_cycle[10515] = 1'b1;  addr_rom[10515]='h000009b4;  wr_data_rom[10515]='h00000678;
    rd_cycle[10516] = 1'b0;  wr_cycle[10516] = 1'b1;  addr_rom[10516]='h00000de0;  wr_data_rom[10516]='h000028f9;
    rd_cycle[10517] = 1'b0;  wr_cycle[10517] = 1'b1;  addr_rom[10517]='h00000e44;  wr_data_rom[10517]='h00002506;
    rd_cycle[10518] = 1'b1;  wr_cycle[10518] = 1'b0;  addr_rom[10518]='h00002110;  wr_data_rom[10518]='h00000000;
    rd_cycle[10519] = 1'b1;  wr_cycle[10519] = 1'b0;  addr_rom[10519]='h00000f0c;  wr_data_rom[10519]='h00000000;
    rd_cycle[10520] = 1'b1;  wr_cycle[10520] = 1'b0;  addr_rom[10520]='h00001cac;  wr_data_rom[10520]='h00000000;
    rd_cycle[10521] = 1'b1;  wr_cycle[10521] = 1'b0;  addr_rom[10521]='h0000142c;  wr_data_rom[10521]='h00000000;
    rd_cycle[10522] = 1'b0;  wr_cycle[10522] = 1'b1;  addr_rom[10522]='h00001c5c;  wr_data_rom[10522]='h00003556;
    rd_cycle[10523] = 1'b1;  wr_cycle[10523] = 1'b0;  addr_rom[10523]='h00003fd8;  wr_data_rom[10523]='h00000000;
    rd_cycle[10524] = 1'b0;  wr_cycle[10524] = 1'b1;  addr_rom[10524]='h00001eb8;  wr_data_rom[10524]='h00001995;
    rd_cycle[10525] = 1'b0;  wr_cycle[10525] = 1'b1;  addr_rom[10525]='h000027e8;  wr_data_rom[10525]='h00001fc5;
    rd_cycle[10526] = 1'b0;  wr_cycle[10526] = 1'b1;  addr_rom[10526]='h000035d8;  wr_data_rom[10526]='h00000597;
    rd_cycle[10527] = 1'b0;  wr_cycle[10527] = 1'b1;  addr_rom[10527]='h00001064;  wr_data_rom[10527]='h0000306f;
    rd_cycle[10528] = 1'b1;  wr_cycle[10528] = 1'b0;  addr_rom[10528]='h00000988;  wr_data_rom[10528]='h00000000;
    rd_cycle[10529] = 1'b0;  wr_cycle[10529] = 1'b1;  addr_rom[10529]='h000015c8;  wr_data_rom[10529]='h000026c0;
    rd_cycle[10530] = 1'b1;  wr_cycle[10530] = 1'b0;  addr_rom[10530]='h00002a3c;  wr_data_rom[10530]='h00000000;
    rd_cycle[10531] = 1'b1;  wr_cycle[10531] = 1'b0;  addr_rom[10531]='h0000009c;  wr_data_rom[10531]='h00000000;
    rd_cycle[10532] = 1'b0;  wr_cycle[10532] = 1'b1;  addr_rom[10532]='h00001f28;  wr_data_rom[10532]='h000029db;
    rd_cycle[10533] = 1'b0;  wr_cycle[10533] = 1'b1;  addr_rom[10533]='h00000f5c;  wr_data_rom[10533]='h00000a67;
    rd_cycle[10534] = 1'b1;  wr_cycle[10534] = 1'b0;  addr_rom[10534]='h00001ef0;  wr_data_rom[10534]='h00000000;
    rd_cycle[10535] = 1'b1;  wr_cycle[10535] = 1'b0;  addr_rom[10535]='h00003c4c;  wr_data_rom[10535]='h00000000;
    rd_cycle[10536] = 1'b0;  wr_cycle[10536] = 1'b1;  addr_rom[10536]='h0000151c;  wr_data_rom[10536]='h00003812;
    rd_cycle[10537] = 1'b0;  wr_cycle[10537] = 1'b1;  addr_rom[10537]='h00000e20;  wr_data_rom[10537]='h00002d01;
    rd_cycle[10538] = 1'b0;  wr_cycle[10538] = 1'b1;  addr_rom[10538]='h000034ac;  wr_data_rom[10538]='h00000cb4;
    rd_cycle[10539] = 1'b1;  wr_cycle[10539] = 1'b0;  addr_rom[10539]='h00000138;  wr_data_rom[10539]='h00000000;
    rd_cycle[10540] = 1'b0;  wr_cycle[10540] = 1'b1;  addr_rom[10540]='h00000274;  wr_data_rom[10540]='h00000962;
    rd_cycle[10541] = 1'b1;  wr_cycle[10541] = 1'b0;  addr_rom[10541]='h00000904;  wr_data_rom[10541]='h00000000;
    rd_cycle[10542] = 1'b1;  wr_cycle[10542] = 1'b0;  addr_rom[10542]='h000011d4;  wr_data_rom[10542]='h00000000;
    rd_cycle[10543] = 1'b0;  wr_cycle[10543] = 1'b1;  addr_rom[10543]='h0000251c;  wr_data_rom[10543]='h0000143d;
    rd_cycle[10544] = 1'b0;  wr_cycle[10544] = 1'b1;  addr_rom[10544]='h000025a8;  wr_data_rom[10544]='h00000e11;
    rd_cycle[10545] = 1'b1;  wr_cycle[10545] = 1'b0;  addr_rom[10545]='h000000f0;  wr_data_rom[10545]='h00000000;
    rd_cycle[10546] = 1'b0;  wr_cycle[10546] = 1'b1;  addr_rom[10546]='h00002468;  wr_data_rom[10546]='h00002a55;
    rd_cycle[10547] = 1'b0;  wr_cycle[10547] = 1'b1;  addr_rom[10547]='h00002680;  wr_data_rom[10547]='h0000120e;
    rd_cycle[10548] = 1'b0;  wr_cycle[10548] = 1'b1;  addr_rom[10548]='h000015ec;  wr_data_rom[10548]='h00000a7d;
    rd_cycle[10549] = 1'b0;  wr_cycle[10549] = 1'b1;  addr_rom[10549]='h00003838;  wr_data_rom[10549]='h000034ab;
    rd_cycle[10550] = 1'b0;  wr_cycle[10550] = 1'b1;  addr_rom[10550]='h000028bc;  wr_data_rom[10550]='h00000486;
    rd_cycle[10551] = 1'b0;  wr_cycle[10551] = 1'b1;  addr_rom[10551]='h00002a2c;  wr_data_rom[10551]='h000024bb;
    rd_cycle[10552] = 1'b0;  wr_cycle[10552] = 1'b1;  addr_rom[10552]='h00001c40;  wr_data_rom[10552]='h00002ded;
    rd_cycle[10553] = 1'b0;  wr_cycle[10553] = 1'b1;  addr_rom[10553]='h000006e0;  wr_data_rom[10553]='h00000d82;
    rd_cycle[10554] = 1'b1;  wr_cycle[10554] = 1'b0;  addr_rom[10554]='h00001fa8;  wr_data_rom[10554]='h00000000;
    rd_cycle[10555] = 1'b0;  wr_cycle[10555] = 1'b1;  addr_rom[10555]='h0000108c;  wr_data_rom[10555]='h000016d4;
    rd_cycle[10556] = 1'b1;  wr_cycle[10556] = 1'b0;  addr_rom[10556]='h0000328c;  wr_data_rom[10556]='h00000000;
    rd_cycle[10557] = 1'b1;  wr_cycle[10557] = 1'b0;  addr_rom[10557]='h00002834;  wr_data_rom[10557]='h00000000;
    rd_cycle[10558] = 1'b0;  wr_cycle[10558] = 1'b1;  addr_rom[10558]='h00002770;  wr_data_rom[10558]='h000035c9;
    rd_cycle[10559] = 1'b0;  wr_cycle[10559] = 1'b1;  addr_rom[10559]='h00000cac;  wr_data_rom[10559]='h00000fe1;
    rd_cycle[10560] = 1'b0;  wr_cycle[10560] = 1'b1;  addr_rom[10560]='h00001bd0;  wr_data_rom[10560]='h000036f0;
    rd_cycle[10561] = 1'b1;  wr_cycle[10561] = 1'b0;  addr_rom[10561]='h000038fc;  wr_data_rom[10561]='h00000000;
    rd_cycle[10562] = 1'b0;  wr_cycle[10562] = 1'b1;  addr_rom[10562]='h00002150;  wr_data_rom[10562]='h000013a5;
    rd_cycle[10563] = 1'b1;  wr_cycle[10563] = 1'b0;  addr_rom[10563]='h00003d28;  wr_data_rom[10563]='h00000000;
    rd_cycle[10564] = 1'b0;  wr_cycle[10564] = 1'b1;  addr_rom[10564]='h0000325c;  wr_data_rom[10564]='h00003c12;
    rd_cycle[10565] = 1'b1;  wr_cycle[10565] = 1'b0;  addr_rom[10565]='h00002a5c;  wr_data_rom[10565]='h00000000;
    rd_cycle[10566] = 1'b1;  wr_cycle[10566] = 1'b0;  addr_rom[10566]='h00002e78;  wr_data_rom[10566]='h00000000;
    rd_cycle[10567] = 1'b0;  wr_cycle[10567] = 1'b1;  addr_rom[10567]='h00000498;  wr_data_rom[10567]='h00002fb9;
    rd_cycle[10568] = 1'b1;  wr_cycle[10568] = 1'b0;  addr_rom[10568]='h00000340;  wr_data_rom[10568]='h00000000;
    rd_cycle[10569] = 1'b1;  wr_cycle[10569] = 1'b0;  addr_rom[10569]='h00002398;  wr_data_rom[10569]='h00000000;
    rd_cycle[10570] = 1'b1;  wr_cycle[10570] = 1'b0;  addr_rom[10570]='h0000250c;  wr_data_rom[10570]='h00000000;
    rd_cycle[10571] = 1'b0;  wr_cycle[10571] = 1'b1;  addr_rom[10571]='h000031c8;  wr_data_rom[10571]='h0000214d;
    rd_cycle[10572] = 1'b1;  wr_cycle[10572] = 1'b0;  addr_rom[10572]='h00002b44;  wr_data_rom[10572]='h00000000;
    rd_cycle[10573] = 1'b1;  wr_cycle[10573] = 1'b0;  addr_rom[10573]='h0000086c;  wr_data_rom[10573]='h00000000;
    rd_cycle[10574] = 1'b0;  wr_cycle[10574] = 1'b1;  addr_rom[10574]='h00003eac;  wr_data_rom[10574]='h00002ce3;
    rd_cycle[10575] = 1'b0;  wr_cycle[10575] = 1'b1;  addr_rom[10575]='h000033b4;  wr_data_rom[10575]='h00000f6d;
    rd_cycle[10576] = 1'b0;  wr_cycle[10576] = 1'b1;  addr_rom[10576]='h00001678;  wr_data_rom[10576]='h00000b47;
    rd_cycle[10577] = 1'b0;  wr_cycle[10577] = 1'b1;  addr_rom[10577]='h000027fc;  wr_data_rom[10577]='h0000109b;
    rd_cycle[10578] = 1'b1;  wr_cycle[10578] = 1'b0;  addr_rom[10578]='h00001b64;  wr_data_rom[10578]='h00000000;
    rd_cycle[10579] = 1'b1;  wr_cycle[10579] = 1'b0;  addr_rom[10579]='h00002484;  wr_data_rom[10579]='h00000000;
    rd_cycle[10580] = 1'b0;  wr_cycle[10580] = 1'b1;  addr_rom[10580]='h00003fb0;  wr_data_rom[10580]='h00002461;
    rd_cycle[10581] = 1'b0;  wr_cycle[10581] = 1'b1;  addr_rom[10581]='h00000dc0;  wr_data_rom[10581]='h00003d3b;
    rd_cycle[10582] = 1'b0;  wr_cycle[10582] = 1'b1;  addr_rom[10582]='h00003f98;  wr_data_rom[10582]='h00002cbd;
    rd_cycle[10583] = 1'b0;  wr_cycle[10583] = 1'b1;  addr_rom[10583]='h00002204;  wr_data_rom[10583]='h00001eaf;
    rd_cycle[10584] = 1'b1;  wr_cycle[10584] = 1'b0;  addr_rom[10584]='h000033c8;  wr_data_rom[10584]='h00000000;
    rd_cycle[10585] = 1'b0;  wr_cycle[10585] = 1'b1;  addr_rom[10585]='h000009a0;  wr_data_rom[10585]='h00000706;
    rd_cycle[10586] = 1'b1;  wr_cycle[10586] = 1'b0;  addr_rom[10586]='h00001aa0;  wr_data_rom[10586]='h00000000;
    rd_cycle[10587] = 1'b1;  wr_cycle[10587] = 1'b0;  addr_rom[10587]='h00001b34;  wr_data_rom[10587]='h00000000;
    rd_cycle[10588] = 1'b0;  wr_cycle[10588] = 1'b1;  addr_rom[10588]='h000034e8;  wr_data_rom[10588]='h000013cb;
    rd_cycle[10589] = 1'b1;  wr_cycle[10589] = 1'b0;  addr_rom[10589]='h00002370;  wr_data_rom[10589]='h00000000;
    rd_cycle[10590] = 1'b0;  wr_cycle[10590] = 1'b1;  addr_rom[10590]='h000033c8;  wr_data_rom[10590]='h000005e1;
    rd_cycle[10591] = 1'b1;  wr_cycle[10591] = 1'b0;  addr_rom[10591]='h0000078c;  wr_data_rom[10591]='h00000000;
    rd_cycle[10592] = 1'b0;  wr_cycle[10592] = 1'b1;  addr_rom[10592]='h00000984;  wr_data_rom[10592]='h00003693;
    rd_cycle[10593] = 1'b0;  wr_cycle[10593] = 1'b1;  addr_rom[10593]='h000002f8;  wr_data_rom[10593]='h00000ce6;
    rd_cycle[10594] = 1'b1;  wr_cycle[10594] = 1'b0;  addr_rom[10594]='h00002f00;  wr_data_rom[10594]='h00000000;
    rd_cycle[10595] = 1'b0;  wr_cycle[10595] = 1'b1;  addr_rom[10595]='h00000d4c;  wr_data_rom[10595]='h00000a3b;
    rd_cycle[10596] = 1'b0;  wr_cycle[10596] = 1'b1;  addr_rom[10596]='h000033c4;  wr_data_rom[10596]='h000013ff;
    rd_cycle[10597] = 1'b0;  wr_cycle[10597] = 1'b1;  addr_rom[10597]='h00002d54;  wr_data_rom[10597]='h00003d61;
    rd_cycle[10598] = 1'b0;  wr_cycle[10598] = 1'b1;  addr_rom[10598]='h000004f8;  wr_data_rom[10598]='h00000495;
    rd_cycle[10599] = 1'b1;  wr_cycle[10599] = 1'b0;  addr_rom[10599]='h00003264;  wr_data_rom[10599]='h00000000;
    rd_cycle[10600] = 1'b0;  wr_cycle[10600] = 1'b1;  addr_rom[10600]='h00003ff4;  wr_data_rom[10600]='h00000d7b;
    rd_cycle[10601] = 1'b0;  wr_cycle[10601] = 1'b1;  addr_rom[10601]='h00002978;  wr_data_rom[10601]='h00002e57;
    rd_cycle[10602] = 1'b1;  wr_cycle[10602] = 1'b0;  addr_rom[10602]='h00002f00;  wr_data_rom[10602]='h00000000;
    rd_cycle[10603] = 1'b0;  wr_cycle[10603] = 1'b1;  addr_rom[10603]='h00001000;  wr_data_rom[10603]='h00001ded;
    rd_cycle[10604] = 1'b0;  wr_cycle[10604] = 1'b1;  addr_rom[10604]='h00003474;  wr_data_rom[10604]='h00002c4e;
    rd_cycle[10605] = 1'b1;  wr_cycle[10605] = 1'b0;  addr_rom[10605]='h00002388;  wr_data_rom[10605]='h00000000;
    rd_cycle[10606] = 1'b0;  wr_cycle[10606] = 1'b1;  addr_rom[10606]='h00000c60;  wr_data_rom[10606]='h000007f9;
    rd_cycle[10607] = 1'b1;  wr_cycle[10607] = 1'b0;  addr_rom[10607]='h00001ad8;  wr_data_rom[10607]='h00000000;
    rd_cycle[10608] = 1'b1;  wr_cycle[10608] = 1'b0;  addr_rom[10608]='h0000098c;  wr_data_rom[10608]='h00000000;
    rd_cycle[10609] = 1'b0;  wr_cycle[10609] = 1'b1;  addr_rom[10609]='h00001dec;  wr_data_rom[10609]='h000024ed;
    rd_cycle[10610] = 1'b1;  wr_cycle[10610] = 1'b0;  addr_rom[10610]='h00003eec;  wr_data_rom[10610]='h00000000;
    rd_cycle[10611] = 1'b0;  wr_cycle[10611] = 1'b1;  addr_rom[10611]='h00001478;  wr_data_rom[10611]='h00001be9;
    rd_cycle[10612] = 1'b1;  wr_cycle[10612] = 1'b0;  addr_rom[10612]='h000031dc;  wr_data_rom[10612]='h00000000;
    rd_cycle[10613] = 1'b1;  wr_cycle[10613] = 1'b0;  addr_rom[10613]='h000001e0;  wr_data_rom[10613]='h00000000;
    rd_cycle[10614] = 1'b0;  wr_cycle[10614] = 1'b1;  addr_rom[10614]='h000032ac;  wr_data_rom[10614]='h000020bd;
    rd_cycle[10615] = 1'b0;  wr_cycle[10615] = 1'b1;  addr_rom[10615]='h00002224;  wr_data_rom[10615]='h00002acb;
    rd_cycle[10616] = 1'b0;  wr_cycle[10616] = 1'b1;  addr_rom[10616]='h000027c0;  wr_data_rom[10616]='h0000073f;
    rd_cycle[10617] = 1'b1;  wr_cycle[10617] = 1'b0;  addr_rom[10617]='h000028c4;  wr_data_rom[10617]='h00000000;
    rd_cycle[10618] = 1'b0;  wr_cycle[10618] = 1'b1;  addr_rom[10618]='h00000e90;  wr_data_rom[10618]='h0000121e;
    rd_cycle[10619] = 1'b0;  wr_cycle[10619] = 1'b1;  addr_rom[10619]='h00001bac;  wr_data_rom[10619]='h00002f42;
    rd_cycle[10620] = 1'b1;  wr_cycle[10620] = 1'b0;  addr_rom[10620]='h000014fc;  wr_data_rom[10620]='h00000000;
    rd_cycle[10621] = 1'b1;  wr_cycle[10621] = 1'b0;  addr_rom[10621]='h00000f20;  wr_data_rom[10621]='h00000000;
    rd_cycle[10622] = 1'b0;  wr_cycle[10622] = 1'b1;  addr_rom[10622]='h000005ec;  wr_data_rom[10622]='h00000276;
    rd_cycle[10623] = 1'b0;  wr_cycle[10623] = 1'b1;  addr_rom[10623]='h0000242c;  wr_data_rom[10623]='h00000638;
    rd_cycle[10624] = 1'b1;  wr_cycle[10624] = 1'b0;  addr_rom[10624]='h00003100;  wr_data_rom[10624]='h00000000;
    rd_cycle[10625] = 1'b1;  wr_cycle[10625] = 1'b0;  addr_rom[10625]='h00000ad4;  wr_data_rom[10625]='h00000000;
    rd_cycle[10626] = 1'b0;  wr_cycle[10626] = 1'b1;  addr_rom[10626]='h00000988;  wr_data_rom[10626]='h00003fcb;
    rd_cycle[10627] = 1'b0;  wr_cycle[10627] = 1'b1;  addr_rom[10627]='h000021cc;  wr_data_rom[10627]='h00001d6c;
    rd_cycle[10628] = 1'b0;  wr_cycle[10628] = 1'b1;  addr_rom[10628]='h000025e8;  wr_data_rom[10628]='h00002316;
    rd_cycle[10629] = 1'b1;  wr_cycle[10629] = 1'b0;  addr_rom[10629]='h00000b44;  wr_data_rom[10629]='h00000000;
    rd_cycle[10630] = 1'b0;  wr_cycle[10630] = 1'b1;  addr_rom[10630]='h00003d60;  wr_data_rom[10630]='h000027de;
    rd_cycle[10631] = 1'b1;  wr_cycle[10631] = 1'b0;  addr_rom[10631]='h00002fc4;  wr_data_rom[10631]='h00000000;
    rd_cycle[10632] = 1'b0;  wr_cycle[10632] = 1'b1;  addr_rom[10632]='h00001300;  wr_data_rom[10632]='h00000e48;
    rd_cycle[10633] = 1'b1;  wr_cycle[10633] = 1'b0;  addr_rom[10633]='h00003754;  wr_data_rom[10633]='h00000000;
    rd_cycle[10634] = 1'b1;  wr_cycle[10634] = 1'b0;  addr_rom[10634]='h000028d4;  wr_data_rom[10634]='h00000000;
    rd_cycle[10635] = 1'b0;  wr_cycle[10635] = 1'b1;  addr_rom[10635]='h0000061c;  wr_data_rom[10635]='h00003266;
    rd_cycle[10636] = 1'b0;  wr_cycle[10636] = 1'b1;  addr_rom[10636]='h00001008;  wr_data_rom[10636]='h00001c9f;
    rd_cycle[10637] = 1'b1;  wr_cycle[10637] = 1'b0;  addr_rom[10637]='h00000130;  wr_data_rom[10637]='h00000000;
    rd_cycle[10638] = 1'b0;  wr_cycle[10638] = 1'b1;  addr_rom[10638]='h000024cc;  wr_data_rom[10638]='h0000050e;
    rd_cycle[10639] = 1'b0;  wr_cycle[10639] = 1'b1;  addr_rom[10639]='h00000d0c;  wr_data_rom[10639]='h00000a6b;
    rd_cycle[10640] = 1'b1;  wr_cycle[10640] = 1'b0;  addr_rom[10640]='h00001334;  wr_data_rom[10640]='h00000000;
    rd_cycle[10641] = 1'b1;  wr_cycle[10641] = 1'b0;  addr_rom[10641]='h00001058;  wr_data_rom[10641]='h00000000;
    rd_cycle[10642] = 1'b1;  wr_cycle[10642] = 1'b0;  addr_rom[10642]='h000021b0;  wr_data_rom[10642]='h00000000;
    rd_cycle[10643] = 1'b1;  wr_cycle[10643] = 1'b0;  addr_rom[10643]='h00000058;  wr_data_rom[10643]='h00000000;
    rd_cycle[10644] = 1'b1;  wr_cycle[10644] = 1'b0;  addr_rom[10644]='h00000214;  wr_data_rom[10644]='h00000000;
    rd_cycle[10645] = 1'b0;  wr_cycle[10645] = 1'b1;  addr_rom[10645]='h00000b14;  wr_data_rom[10645]='h00002075;
    rd_cycle[10646] = 1'b1;  wr_cycle[10646] = 1'b0;  addr_rom[10646]='h00000a50;  wr_data_rom[10646]='h00000000;
    rd_cycle[10647] = 1'b1;  wr_cycle[10647] = 1'b0;  addr_rom[10647]='h0000218c;  wr_data_rom[10647]='h00000000;
    rd_cycle[10648] = 1'b1;  wr_cycle[10648] = 1'b0;  addr_rom[10648]='h00003d04;  wr_data_rom[10648]='h00000000;
    rd_cycle[10649] = 1'b1;  wr_cycle[10649] = 1'b0;  addr_rom[10649]='h00002e24;  wr_data_rom[10649]='h00000000;
    rd_cycle[10650] = 1'b1;  wr_cycle[10650] = 1'b0;  addr_rom[10650]='h000025e4;  wr_data_rom[10650]='h00000000;
    rd_cycle[10651] = 1'b1;  wr_cycle[10651] = 1'b0;  addr_rom[10651]='h00000798;  wr_data_rom[10651]='h00000000;
    rd_cycle[10652] = 1'b1;  wr_cycle[10652] = 1'b0;  addr_rom[10652]='h000005f0;  wr_data_rom[10652]='h00000000;
    rd_cycle[10653] = 1'b0;  wr_cycle[10653] = 1'b1;  addr_rom[10653]='h00002404;  wr_data_rom[10653]='h00003ee7;
    rd_cycle[10654] = 1'b1;  wr_cycle[10654] = 1'b0;  addr_rom[10654]='h000017a4;  wr_data_rom[10654]='h00000000;
    rd_cycle[10655] = 1'b1;  wr_cycle[10655] = 1'b0;  addr_rom[10655]='h0000197c;  wr_data_rom[10655]='h00000000;
    rd_cycle[10656] = 1'b1;  wr_cycle[10656] = 1'b0;  addr_rom[10656]='h0000343c;  wr_data_rom[10656]='h00000000;
    rd_cycle[10657] = 1'b0;  wr_cycle[10657] = 1'b1;  addr_rom[10657]='h00002a0c;  wr_data_rom[10657]='h000010e8;
    rd_cycle[10658] = 1'b0;  wr_cycle[10658] = 1'b1;  addr_rom[10658]='h00000434;  wr_data_rom[10658]='h0000090e;
    rd_cycle[10659] = 1'b1;  wr_cycle[10659] = 1'b0;  addr_rom[10659]='h00002500;  wr_data_rom[10659]='h00000000;
    rd_cycle[10660] = 1'b0;  wr_cycle[10660] = 1'b1;  addr_rom[10660]='h00002d20;  wr_data_rom[10660]='h000014bf;
    rd_cycle[10661] = 1'b0;  wr_cycle[10661] = 1'b1;  addr_rom[10661]='h00001524;  wr_data_rom[10661]='h00000e09;
    rd_cycle[10662] = 1'b1;  wr_cycle[10662] = 1'b0;  addr_rom[10662]='h00000be0;  wr_data_rom[10662]='h00000000;
    rd_cycle[10663] = 1'b0;  wr_cycle[10663] = 1'b1;  addr_rom[10663]='h00000d00;  wr_data_rom[10663]='h000031d9;
    rd_cycle[10664] = 1'b0;  wr_cycle[10664] = 1'b1;  addr_rom[10664]='h000027bc;  wr_data_rom[10664]='h000017cf;
    rd_cycle[10665] = 1'b0;  wr_cycle[10665] = 1'b1;  addr_rom[10665]='h00002120;  wr_data_rom[10665]='h0000148f;
    rd_cycle[10666] = 1'b0;  wr_cycle[10666] = 1'b1;  addr_rom[10666]='h00001228;  wr_data_rom[10666]='h00002d54;
    rd_cycle[10667] = 1'b1;  wr_cycle[10667] = 1'b0;  addr_rom[10667]='h00003c10;  wr_data_rom[10667]='h00000000;
    rd_cycle[10668] = 1'b1;  wr_cycle[10668] = 1'b0;  addr_rom[10668]='h00001aa4;  wr_data_rom[10668]='h00000000;
    rd_cycle[10669] = 1'b1;  wr_cycle[10669] = 1'b0;  addr_rom[10669]='h000007b0;  wr_data_rom[10669]='h00000000;
    rd_cycle[10670] = 1'b0;  wr_cycle[10670] = 1'b1;  addr_rom[10670]='h000007d0;  wr_data_rom[10670]='h0000289c;
    rd_cycle[10671] = 1'b0;  wr_cycle[10671] = 1'b1;  addr_rom[10671]='h000038e8;  wr_data_rom[10671]='h000037d3;
    rd_cycle[10672] = 1'b0;  wr_cycle[10672] = 1'b1;  addr_rom[10672]='h00001d34;  wr_data_rom[10672]='h00000607;
    rd_cycle[10673] = 1'b1;  wr_cycle[10673] = 1'b0;  addr_rom[10673]='h00002a9c;  wr_data_rom[10673]='h00000000;
    rd_cycle[10674] = 1'b1;  wr_cycle[10674] = 1'b0;  addr_rom[10674]='h00002ca0;  wr_data_rom[10674]='h00000000;
    rd_cycle[10675] = 1'b1;  wr_cycle[10675] = 1'b0;  addr_rom[10675]='h00003960;  wr_data_rom[10675]='h00000000;
    rd_cycle[10676] = 1'b1;  wr_cycle[10676] = 1'b0;  addr_rom[10676]='h000026f0;  wr_data_rom[10676]='h00000000;
    rd_cycle[10677] = 1'b1;  wr_cycle[10677] = 1'b0;  addr_rom[10677]='h000031fc;  wr_data_rom[10677]='h00000000;
    rd_cycle[10678] = 1'b0;  wr_cycle[10678] = 1'b1;  addr_rom[10678]='h0000091c;  wr_data_rom[10678]='h000008e2;
    rd_cycle[10679] = 1'b0;  wr_cycle[10679] = 1'b1;  addr_rom[10679]='h00003c6c;  wr_data_rom[10679]='h000003aa;
    rd_cycle[10680] = 1'b0;  wr_cycle[10680] = 1'b1;  addr_rom[10680]='h00001aa8;  wr_data_rom[10680]='h00002d72;
    rd_cycle[10681] = 1'b1;  wr_cycle[10681] = 1'b0;  addr_rom[10681]='h00001f04;  wr_data_rom[10681]='h00000000;
    rd_cycle[10682] = 1'b0;  wr_cycle[10682] = 1'b1;  addr_rom[10682]='h00002ac8;  wr_data_rom[10682]='h00001761;
    rd_cycle[10683] = 1'b1;  wr_cycle[10683] = 1'b0;  addr_rom[10683]='h00000c4c;  wr_data_rom[10683]='h00000000;
    rd_cycle[10684] = 1'b0;  wr_cycle[10684] = 1'b1;  addr_rom[10684]='h00000c54;  wr_data_rom[10684]='h00002ae9;
    rd_cycle[10685] = 1'b0;  wr_cycle[10685] = 1'b1;  addr_rom[10685]='h00003e9c;  wr_data_rom[10685]='h0000339f;
    rd_cycle[10686] = 1'b1;  wr_cycle[10686] = 1'b0;  addr_rom[10686]='h00000768;  wr_data_rom[10686]='h00000000;
    rd_cycle[10687] = 1'b0;  wr_cycle[10687] = 1'b1;  addr_rom[10687]='h00003124;  wr_data_rom[10687]='h0000117b;
    rd_cycle[10688] = 1'b0;  wr_cycle[10688] = 1'b1;  addr_rom[10688]='h00002700;  wr_data_rom[10688]='h0000107f;
    rd_cycle[10689] = 1'b0;  wr_cycle[10689] = 1'b1;  addr_rom[10689]='h00000e44;  wr_data_rom[10689]='h000008a5;
    rd_cycle[10690] = 1'b0;  wr_cycle[10690] = 1'b1;  addr_rom[10690]='h00002ca8;  wr_data_rom[10690]='h000017f9;
    rd_cycle[10691] = 1'b0;  wr_cycle[10691] = 1'b1;  addr_rom[10691]='h000014ac;  wr_data_rom[10691]='h000007de;
    rd_cycle[10692] = 1'b1;  wr_cycle[10692] = 1'b0;  addr_rom[10692]='h00000c50;  wr_data_rom[10692]='h00000000;
    rd_cycle[10693] = 1'b1;  wr_cycle[10693] = 1'b0;  addr_rom[10693]='h000003d4;  wr_data_rom[10693]='h00000000;
    rd_cycle[10694] = 1'b0;  wr_cycle[10694] = 1'b1;  addr_rom[10694]='h000015ac;  wr_data_rom[10694]='h0000173b;
    rd_cycle[10695] = 1'b1;  wr_cycle[10695] = 1'b0;  addr_rom[10695]='h000013b8;  wr_data_rom[10695]='h00000000;
    rd_cycle[10696] = 1'b0;  wr_cycle[10696] = 1'b1;  addr_rom[10696]='h000030d4;  wr_data_rom[10696]='h00001cd2;
    rd_cycle[10697] = 1'b1;  wr_cycle[10697] = 1'b0;  addr_rom[10697]='h0000374c;  wr_data_rom[10697]='h00000000;
    rd_cycle[10698] = 1'b0;  wr_cycle[10698] = 1'b1;  addr_rom[10698]='h00002dec;  wr_data_rom[10698]='h000035d7;
    rd_cycle[10699] = 1'b0;  wr_cycle[10699] = 1'b1;  addr_rom[10699]='h00003e40;  wr_data_rom[10699]='h000011c4;
    rd_cycle[10700] = 1'b0;  wr_cycle[10700] = 1'b1;  addr_rom[10700]='h00001150;  wr_data_rom[10700]='h00001466;
    rd_cycle[10701] = 1'b1;  wr_cycle[10701] = 1'b0;  addr_rom[10701]='h000030d0;  wr_data_rom[10701]='h00000000;
    rd_cycle[10702] = 1'b0;  wr_cycle[10702] = 1'b1;  addr_rom[10702]='h0000160c;  wr_data_rom[10702]='h00002bd3;
    rd_cycle[10703] = 1'b1;  wr_cycle[10703] = 1'b0;  addr_rom[10703]='h0000152c;  wr_data_rom[10703]='h00000000;
    rd_cycle[10704] = 1'b1;  wr_cycle[10704] = 1'b0;  addr_rom[10704]='h00001d5c;  wr_data_rom[10704]='h00000000;
    rd_cycle[10705] = 1'b0;  wr_cycle[10705] = 1'b1;  addr_rom[10705]='h00000afc;  wr_data_rom[10705]='h00001a39;
    rd_cycle[10706] = 1'b0;  wr_cycle[10706] = 1'b1;  addr_rom[10706]='h00001548;  wr_data_rom[10706]='h0000011f;
    rd_cycle[10707] = 1'b0;  wr_cycle[10707] = 1'b1;  addr_rom[10707]='h000001c4;  wr_data_rom[10707]='h00003fe7;
    rd_cycle[10708] = 1'b0;  wr_cycle[10708] = 1'b1;  addr_rom[10708]='h000025d8;  wr_data_rom[10708]='h0000388a;
    rd_cycle[10709] = 1'b0;  wr_cycle[10709] = 1'b1;  addr_rom[10709]='h0000186c;  wr_data_rom[10709]='h000033d1;
    rd_cycle[10710] = 1'b0;  wr_cycle[10710] = 1'b1;  addr_rom[10710]='h00001594;  wr_data_rom[10710]='h00001d4c;
    rd_cycle[10711] = 1'b0;  wr_cycle[10711] = 1'b1;  addr_rom[10711]='h00001380;  wr_data_rom[10711]='h00002a93;
    rd_cycle[10712] = 1'b1;  wr_cycle[10712] = 1'b0;  addr_rom[10712]='h00003e70;  wr_data_rom[10712]='h00000000;
    rd_cycle[10713] = 1'b1;  wr_cycle[10713] = 1'b0;  addr_rom[10713]='h0000160c;  wr_data_rom[10713]='h00000000;
    rd_cycle[10714] = 1'b0;  wr_cycle[10714] = 1'b1;  addr_rom[10714]='h00003e78;  wr_data_rom[10714]='h00001520;
    rd_cycle[10715] = 1'b0;  wr_cycle[10715] = 1'b1;  addr_rom[10715]='h000020d0;  wr_data_rom[10715]='h0000112e;
    rd_cycle[10716] = 1'b0;  wr_cycle[10716] = 1'b1;  addr_rom[10716]='h000015ac;  wr_data_rom[10716]='h00000799;
    rd_cycle[10717] = 1'b0;  wr_cycle[10717] = 1'b1;  addr_rom[10717]='h00002b84;  wr_data_rom[10717]='h00002f56;
    rd_cycle[10718] = 1'b1;  wr_cycle[10718] = 1'b0;  addr_rom[10718]='h000028cc;  wr_data_rom[10718]='h00000000;
    rd_cycle[10719] = 1'b0;  wr_cycle[10719] = 1'b1;  addr_rom[10719]='h00002c54;  wr_data_rom[10719]='h000023fb;
    rd_cycle[10720] = 1'b0;  wr_cycle[10720] = 1'b1;  addr_rom[10720]='h00002218;  wr_data_rom[10720]='h000032d1;
    rd_cycle[10721] = 1'b0;  wr_cycle[10721] = 1'b1;  addr_rom[10721]='h000000c8;  wr_data_rom[10721]='h0000092e;
    rd_cycle[10722] = 1'b0;  wr_cycle[10722] = 1'b1;  addr_rom[10722]='h00000fc0;  wr_data_rom[10722]='h00003ec4;
    rd_cycle[10723] = 1'b0;  wr_cycle[10723] = 1'b1;  addr_rom[10723]='h000009c8;  wr_data_rom[10723]='h00003ed6;
    rd_cycle[10724] = 1'b1;  wr_cycle[10724] = 1'b0;  addr_rom[10724]='h00002564;  wr_data_rom[10724]='h00000000;
    rd_cycle[10725] = 1'b0;  wr_cycle[10725] = 1'b1;  addr_rom[10725]='h00003a3c;  wr_data_rom[10725]='h0000097b;
    rd_cycle[10726] = 1'b1;  wr_cycle[10726] = 1'b0;  addr_rom[10726]='h00002a58;  wr_data_rom[10726]='h00000000;
    rd_cycle[10727] = 1'b0;  wr_cycle[10727] = 1'b1;  addr_rom[10727]='h00000ad4;  wr_data_rom[10727]='h000024ca;
    rd_cycle[10728] = 1'b0;  wr_cycle[10728] = 1'b1;  addr_rom[10728]='h00000e98;  wr_data_rom[10728]='h0000021f;
    rd_cycle[10729] = 1'b1;  wr_cycle[10729] = 1'b0;  addr_rom[10729]='h0000247c;  wr_data_rom[10729]='h00000000;
    rd_cycle[10730] = 1'b0;  wr_cycle[10730] = 1'b1;  addr_rom[10730]='h000012d0;  wr_data_rom[10730]='h000003c6;
    rd_cycle[10731] = 1'b1;  wr_cycle[10731] = 1'b0;  addr_rom[10731]='h00002148;  wr_data_rom[10731]='h00000000;
    rd_cycle[10732] = 1'b1;  wr_cycle[10732] = 1'b0;  addr_rom[10732]='h00002f54;  wr_data_rom[10732]='h00000000;
    rd_cycle[10733] = 1'b0;  wr_cycle[10733] = 1'b1;  addr_rom[10733]='h00002608;  wr_data_rom[10733]='h00003742;
    rd_cycle[10734] = 1'b0;  wr_cycle[10734] = 1'b1;  addr_rom[10734]='h00001d88;  wr_data_rom[10734]='h000021fd;
    rd_cycle[10735] = 1'b0;  wr_cycle[10735] = 1'b1;  addr_rom[10735]='h00001acc;  wr_data_rom[10735]='h00003b7a;
    rd_cycle[10736] = 1'b1;  wr_cycle[10736] = 1'b0;  addr_rom[10736]='h00001c80;  wr_data_rom[10736]='h00000000;
    rd_cycle[10737] = 1'b1;  wr_cycle[10737] = 1'b0;  addr_rom[10737]='h00002b1c;  wr_data_rom[10737]='h00000000;
    rd_cycle[10738] = 1'b1;  wr_cycle[10738] = 1'b0;  addr_rom[10738]='h00000eb4;  wr_data_rom[10738]='h00000000;
    rd_cycle[10739] = 1'b1;  wr_cycle[10739] = 1'b0;  addr_rom[10739]='h00001620;  wr_data_rom[10739]='h00000000;
    rd_cycle[10740] = 1'b0;  wr_cycle[10740] = 1'b1;  addr_rom[10740]='h000000f0;  wr_data_rom[10740]='h00000e8c;
    rd_cycle[10741] = 1'b0;  wr_cycle[10741] = 1'b1;  addr_rom[10741]='h00003e90;  wr_data_rom[10741]='h00001030;
    rd_cycle[10742] = 1'b1;  wr_cycle[10742] = 1'b0;  addr_rom[10742]='h000003f4;  wr_data_rom[10742]='h00000000;
    rd_cycle[10743] = 1'b1;  wr_cycle[10743] = 1'b0;  addr_rom[10743]='h000024ac;  wr_data_rom[10743]='h00000000;
    rd_cycle[10744] = 1'b0;  wr_cycle[10744] = 1'b1;  addr_rom[10744]='h00000fec;  wr_data_rom[10744]='h00002845;
    rd_cycle[10745] = 1'b0;  wr_cycle[10745] = 1'b1;  addr_rom[10745]='h00002f8c;  wr_data_rom[10745]='h00000505;
    rd_cycle[10746] = 1'b1;  wr_cycle[10746] = 1'b0;  addr_rom[10746]='h00002c1c;  wr_data_rom[10746]='h00000000;
    rd_cycle[10747] = 1'b0;  wr_cycle[10747] = 1'b1;  addr_rom[10747]='h00000f28;  wr_data_rom[10747]='h00001ce0;
    rd_cycle[10748] = 1'b1;  wr_cycle[10748] = 1'b0;  addr_rom[10748]='h00002400;  wr_data_rom[10748]='h00000000;
    rd_cycle[10749] = 1'b0;  wr_cycle[10749] = 1'b1;  addr_rom[10749]='h00000b1c;  wr_data_rom[10749]='h00003ade;
    rd_cycle[10750] = 1'b1;  wr_cycle[10750] = 1'b0;  addr_rom[10750]='h00002cb8;  wr_data_rom[10750]='h00000000;
    rd_cycle[10751] = 1'b0;  wr_cycle[10751] = 1'b1;  addr_rom[10751]='h00001f18;  wr_data_rom[10751]='h00001980;
    rd_cycle[10752] = 1'b0;  wr_cycle[10752] = 1'b1;  addr_rom[10752]='h00000400;  wr_data_rom[10752]='h0000177b;
    rd_cycle[10753] = 1'b1;  wr_cycle[10753] = 1'b0;  addr_rom[10753]='h00000794;  wr_data_rom[10753]='h00000000;
    rd_cycle[10754] = 1'b0;  wr_cycle[10754] = 1'b1;  addr_rom[10754]='h00002cb4;  wr_data_rom[10754]='h00000526;
    rd_cycle[10755] = 1'b0;  wr_cycle[10755] = 1'b1;  addr_rom[10755]='h00001e1c;  wr_data_rom[10755]='h0000108e;
    rd_cycle[10756] = 1'b1;  wr_cycle[10756] = 1'b0;  addr_rom[10756]='h00002060;  wr_data_rom[10756]='h00000000;
    rd_cycle[10757] = 1'b1;  wr_cycle[10757] = 1'b0;  addr_rom[10757]='h0000133c;  wr_data_rom[10757]='h00000000;
    rd_cycle[10758] = 1'b0;  wr_cycle[10758] = 1'b1;  addr_rom[10758]='h00003db8;  wr_data_rom[10758]='h0000354c;
    rd_cycle[10759] = 1'b0;  wr_cycle[10759] = 1'b1;  addr_rom[10759]='h000028f0;  wr_data_rom[10759]='h00001ad5;
    rd_cycle[10760] = 1'b0;  wr_cycle[10760] = 1'b1;  addr_rom[10760]='h00002220;  wr_data_rom[10760]='h00003a6f;
    rd_cycle[10761] = 1'b1;  wr_cycle[10761] = 1'b0;  addr_rom[10761]='h000013b4;  wr_data_rom[10761]='h00000000;
    rd_cycle[10762] = 1'b0;  wr_cycle[10762] = 1'b1;  addr_rom[10762]='h000034c4;  wr_data_rom[10762]='h00003a8d;
    rd_cycle[10763] = 1'b1;  wr_cycle[10763] = 1'b0;  addr_rom[10763]='h00001c68;  wr_data_rom[10763]='h00000000;
    rd_cycle[10764] = 1'b0;  wr_cycle[10764] = 1'b1;  addr_rom[10764]='h00003a88;  wr_data_rom[10764]='h00003a1b;
    rd_cycle[10765] = 1'b0;  wr_cycle[10765] = 1'b1;  addr_rom[10765]='h0000052c;  wr_data_rom[10765]='h000018dc;
    rd_cycle[10766] = 1'b1;  wr_cycle[10766] = 1'b0;  addr_rom[10766]='h00002ce8;  wr_data_rom[10766]='h00000000;
    rd_cycle[10767] = 1'b0;  wr_cycle[10767] = 1'b1;  addr_rom[10767]='h000033a4;  wr_data_rom[10767]='h00001b64;
    rd_cycle[10768] = 1'b0;  wr_cycle[10768] = 1'b1;  addr_rom[10768]='h00000518;  wr_data_rom[10768]='h00003978;
    rd_cycle[10769] = 1'b0;  wr_cycle[10769] = 1'b1;  addr_rom[10769]='h000031b0;  wr_data_rom[10769]='h00002fb4;
    rd_cycle[10770] = 1'b0;  wr_cycle[10770] = 1'b1;  addr_rom[10770]='h00000ca8;  wr_data_rom[10770]='h00001149;
    rd_cycle[10771] = 1'b0;  wr_cycle[10771] = 1'b1;  addr_rom[10771]='h00003648;  wr_data_rom[10771]='h00001520;
    rd_cycle[10772] = 1'b0;  wr_cycle[10772] = 1'b1;  addr_rom[10772]='h00003f1c;  wr_data_rom[10772]='h0000292a;
    rd_cycle[10773] = 1'b0;  wr_cycle[10773] = 1'b1;  addr_rom[10773]='h000010f4;  wr_data_rom[10773]='h00003552;
    rd_cycle[10774] = 1'b0;  wr_cycle[10774] = 1'b1;  addr_rom[10774]='h00002eb4;  wr_data_rom[10774]='h000001af;
    rd_cycle[10775] = 1'b1;  wr_cycle[10775] = 1'b0;  addr_rom[10775]='h00003900;  wr_data_rom[10775]='h00000000;
    rd_cycle[10776] = 1'b0;  wr_cycle[10776] = 1'b1;  addr_rom[10776]='h00000b08;  wr_data_rom[10776]='h000010a1;
    rd_cycle[10777] = 1'b0;  wr_cycle[10777] = 1'b1;  addr_rom[10777]='h00002288;  wr_data_rom[10777]='h00000796;
    rd_cycle[10778] = 1'b1;  wr_cycle[10778] = 1'b0;  addr_rom[10778]='h000038b4;  wr_data_rom[10778]='h00000000;
    rd_cycle[10779] = 1'b0;  wr_cycle[10779] = 1'b1;  addr_rom[10779]='h000007b0;  wr_data_rom[10779]='h00003949;
    rd_cycle[10780] = 1'b1;  wr_cycle[10780] = 1'b0;  addr_rom[10780]='h000022fc;  wr_data_rom[10780]='h00000000;
    rd_cycle[10781] = 1'b0;  wr_cycle[10781] = 1'b1;  addr_rom[10781]='h00003be4;  wr_data_rom[10781]='h000028f2;
    rd_cycle[10782] = 1'b0;  wr_cycle[10782] = 1'b1;  addr_rom[10782]='h000019dc;  wr_data_rom[10782]='h00003382;
    rd_cycle[10783] = 1'b1;  wr_cycle[10783] = 1'b0;  addr_rom[10783]='h00003a50;  wr_data_rom[10783]='h00000000;
    rd_cycle[10784] = 1'b0;  wr_cycle[10784] = 1'b1;  addr_rom[10784]='h00002374;  wr_data_rom[10784]='h0000190c;
    rd_cycle[10785] = 1'b1;  wr_cycle[10785] = 1'b0;  addr_rom[10785]='h0000334c;  wr_data_rom[10785]='h00000000;
    rd_cycle[10786] = 1'b1;  wr_cycle[10786] = 1'b0;  addr_rom[10786]='h00002fa4;  wr_data_rom[10786]='h00000000;
    rd_cycle[10787] = 1'b1;  wr_cycle[10787] = 1'b0;  addr_rom[10787]='h000019bc;  wr_data_rom[10787]='h00000000;
    rd_cycle[10788] = 1'b1;  wr_cycle[10788] = 1'b0;  addr_rom[10788]='h00003094;  wr_data_rom[10788]='h00000000;
    rd_cycle[10789] = 1'b1;  wr_cycle[10789] = 1'b0;  addr_rom[10789]='h000029f4;  wr_data_rom[10789]='h00000000;
    rd_cycle[10790] = 1'b0;  wr_cycle[10790] = 1'b1;  addr_rom[10790]='h00003528;  wr_data_rom[10790]='h00001fb8;
    rd_cycle[10791] = 1'b0;  wr_cycle[10791] = 1'b1;  addr_rom[10791]='h00000480;  wr_data_rom[10791]='h000008ae;
    rd_cycle[10792] = 1'b0;  wr_cycle[10792] = 1'b1;  addr_rom[10792]='h00000bfc;  wr_data_rom[10792]='h000018f5;
    rd_cycle[10793] = 1'b0;  wr_cycle[10793] = 1'b1;  addr_rom[10793]='h0000113c;  wr_data_rom[10793]='h0000109a;
    rd_cycle[10794] = 1'b0;  wr_cycle[10794] = 1'b1;  addr_rom[10794]='h000035c8;  wr_data_rom[10794]='h0000236d;
    rd_cycle[10795] = 1'b1;  wr_cycle[10795] = 1'b0;  addr_rom[10795]='h00001794;  wr_data_rom[10795]='h00000000;
    rd_cycle[10796] = 1'b1;  wr_cycle[10796] = 1'b0;  addr_rom[10796]='h00000be4;  wr_data_rom[10796]='h00000000;
    rd_cycle[10797] = 1'b0;  wr_cycle[10797] = 1'b1;  addr_rom[10797]='h00001bc4;  wr_data_rom[10797]='h00001318;
    rd_cycle[10798] = 1'b1;  wr_cycle[10798] = 1'b0;  addr_rom[10798]='h00001128;  wr_data_rom[10798]='h00000000;
    rd_cycle[10799] = 1'b1;  wr_cycle[10799] = 1'b0;  addr_rom[10799]='h00003c04;  wr_data_rom[10799]='h00000000;
    rd_cycle[10800] = 1'b1;  wr_cycle[10800] = 1'b0;  addr_rom[10800]='h00001274;  wr_data_rom[10800]='h00000000;
    rd_cycle[10801] = 1'b1;  wr_cycle[10801] = 1'b0;  addr_rom[10801]='h00002110;  wr_data_rom[10801]='h00000000;
    rd_cycle[10802] = 1'b0;  wr_cycle[10802] = 1'b1;  addr_rom[10802]='h000027e8;  wr_data_rom[10802]='h000014f1;
    rd_cycle[10803] = 1'b1;  wr_cycle[10803] = 1'b0;  addr_rom[10803]='h00001ccc;  wr_data_rom[10803]='h00000000;
    rd_cycle[10804] = 1'b0;  wr_cycle[10804] = 1'b1;  addr_rom[10804]='h00001540;  wr_data_rom[10804]='h0000325e;
    rd_cycle[10805] = 1'b0;  wr_cycle[10805] = 1'b1;  addr_rom[10805]='h00000674;  wr_data_rom[10805]='h000035b4;
    rd_cycle[10806] = 1'b1;  wr_cycle[10806] = 1'b0;  addr_rom[10806]='h00003a40;  wr_data_rom[10806]='h00000000;
    rd_cycle[10807] = 1'b1;  wr_cycle[10807] = 1'b0;  addr_rom[10807]='h000033e4;  wr_data_rom[10807]='h00000000;
    rd_cycle[10808] = 1'b1;  wr_cycle[10808] = 1'b0;  addr_rom[10808]='h00002cfc;  wr_data_rom[10808]='h00000000;
    rd_cycle[10809] = 1'b0;  wr_cycle[10809] = 1'b1;  addr_rom[10809]='h00001024;  wr_data_rom[10809]='h00000dac;
    rd_cycle[10810] = 1'b0;  wr_cycle[10810] = 1'b1;  addr_rom[10810]='h00002174;  wr_data_rom[10810]='h00001f69;
    rd_cycle[10811] = 1'b1;  wr_cycle[10811] = 1'b0;  addr_rom[10811]='h0000156c;  wr_data_rom[10811]='h00000000;
    rd_cycle[10812] = 1'b0;  wr_cycle[10812] = 1'b1;  addr_rom[10812]='h00003574;  wr_data_rom[10812]='h00001704;
    rd_cycle[10813] = 1'b0;  wr_cycle[10813] = 1'b1;  addr_rom[10813]='h000032f0;  wr_data_rom[10813]='h000032a8;
    rd_cycle[10814] = 1'b1;  wr_cycle[10814] = 1'b0;  addr_rom[10814]='h00002ab8;  wr_data_rom[10814]='h00000000;
    rd_cycle[10815] = 1'b0;  wr_cycle[10815] = 1'b1;  addr_rom[10815]='h0000007c;  wr_data_rom[10815]='h00003d8c;
    rd_cycle[10816] = 1'b1;  wr_cycle[10816] = 1'b0;  addr_rom[10816]='h00003118;  wr_data_rom[10816]='h00000000;
    rd_cycle[10817] = 1'b1;  wr_cycle[10817] = 1'b0;  addr_rom[10817]='h0000323c;  wr_data_rom[10817]='h00000000;
    rd_cycle[10818] = 1'b0;  wr_cycle[10818] = 1'b1;  addr_rom[10818]='h000028e8;  wr_data_rom[10818]='h00001ed0;
    rd_cycle[10819] = 1'b0;  wr_cycle[10819] = 1'b1;  addr_rom[10819]='h00003b2c;  wr_data_rom[10819]='h00003ee3;
    rd_cycle[10820] = 1'b1;  wr_cycle[10820] = 1'b0;  addr_rom[10820]='h00001f50;  wr_data_rom[10820]='h00000000;
    rd_cycle[10821] = 1'b0;  wr_cycle[10821] = 1'b1;  addr_rom[10821]='h0000167c;  wr_data_rom[10821]='h0000040e;
    rd_cycle[10822] = 1'b1;  wr_cycle[10822] = 1'b0;  addr_rom[10822]='h00001cc4;  wr_data_rom[10822]='h00000000;
    rd_cycle[10823] = 1'b0;  wr_cycle[10823] = 1'b1;  addr_rom[10823]='h00003180;  wr_data_rom[10823]='h00003da0;
    rd_cycle[10824] = 1'b0;  wr_cycle[10824] = 1'b1;  addr_rom[10824]='h00003604;  wr_data_rom[10824]='h000020ea;
    rd_cycle[10825] = 1'b0;  wr_cycle[10825] = 1'b1;  addr_rom[10825]='h00001160;  wr_data_rom[10825]='h00001d76;
    rd_cycle[10826] = 1'b1;  wr_cycle[10826] = 1'b0;  addr_rom[10826]='h00000d34;  wr_data_rom[10826]='h00000000;
    rd_cycle[10827] = 1'b1;  wr_cycle[10827] = 1'b0;  addr_rom[10827]='h00002bc4;  wr_data_rom[10827]='h00000000;
    rd_cycle[10828] = 1'b0;  wr_cycle[10828] = 1'b1;  addr_rom[10828]='h00001da4;  wr_data_rom[10828]='h00001121;
    rd_cycle[10829] = 1'b0;  wr_cycle[10829] = 1'b1;  addr_rom[10829]='h00003c30;  wr_data_rom[10829]='h000023aa;
    rd_cycle[10830] = 1'b0;  wr_cycle[10830] = 1'b1;  addr_rom[10830]='h00002718;  wr_data_rom[10830]='h000023fe;
    rd_cycle[10831] = 1'b0;  wr_cycle[10831] = 1'b1;  addr_rom[10831]='h000039ac;  wr_data_rom[10831]='h00003ac3;
    rd_cycle[10832] = 1'b0;  wr_cycle[10832] = 1'b1;  addr_rom[10832]='h0000193c;  wr_data_rom[10832]='h00002fb0;
    rd_cycle[10833] = 1'b1;  wr_cycle[10833] = 1'b0;  addr_rom[10833]='h000000ec;  wr_data_rom[10833]='h00000000;
    rd_cycle[10834] = 1'b1;  wr_cycle[10834] = 1'b0;  addr_rom[10834]='h00002e80;  wr_data_rom[10834]='h00000000;
    rd_cycle[10835] = 1'b0;  wr_cycle[10835] = 1'b1;  addr_rom[10835]='h00000b04;  wr_data_rom[10835]='h00003d38;
    rd_cycle[10836] = 1'b0;  wr_cycle[10836] = 1'b1;  addr_rom[10836]='h00003ea8;  wr_data_rom[10836]='h00000389;
    rd_cycle[10837] = 1'b1;  wr_cycle[10837] = 1'b0;  addr_rom[10837]='h000001a8;  wr_data_rom[10837]='h00000000;
    rd_cycle[10838] = 1'b1;  wr_cycle[10838] = 1'b0;  addr_rom[10838]='h000014c0;  wr_data_rom[10838]='h00000000;
    rd_cycle[10839] = 1'b0;  wr_cycle[10839] = 1'b1;  addr_rom[10839]='h00000778;  wr_data_rom[10839]='h00001597;
    rd_cycle[10840] = 1'b0;  wr_cycle[10840] = 1'b1;  addr_rom[10840]='h00002594;  wr_data_rom[10840]='h0000349d;
    rd_cycle[10841] = 1'b1;  wr_cycle[10841] = 1'b0;  addr_rom[10841]='h00001cbc;  wr_data_rom[10841]='h00000000;
    rd_cycle[10842] = 1'b1;  wr_cycle[10842] = 1'b0;  addr_rom[10842]='h000039bc;  wr_data_rom[10842]='h00000000;
    rd_cycle[10843] = 1'b0;  wr_cycle[10843] = 1'b1;  addr_rom[10843]='h00000868;  wr_data_rom[10843]='h00002958;
    rd_cycle[10844] = 1'b0;  wr_cycle[10844] = 1'b1;  addr_rom[10844]='h00001fa0;  wr_data_rom[10844]='h000034c4;
    rd_cycle[10845] = 1'b1;  wr_cycle[10845] = 1'b0;  addr_rom[10845]='h000006c4;  wr_data_rom[10845]='h00000000;
    rd_cycle[10846] = 1'b0;  wr_cycle[10846] = 1'b1;  addr_rom[10846]='h000004b0;  wr_data_rom[10846]='h00000e21;
    rd_cycle[10847] = 1'b1;  wr_cycle[10847] = 1'b0;  addr_rom[10847]='h000020a8;  wr_data_rom[10847]='h00000000;
    rd_cycle[10848] = 1'b1;  wr_cycle[10848] = 1'b0;  addr_rom[10848]='h000010c8;  wr_data_rom[10848]='h00000000;
    rd_cycle[10849] = 1'b1;  wr_cycle[10849] = 1'b0;  addr_rom[10849]='h0000208c;  wr_data_rom[10849]='h00000000;
    rd_cycle[10850] = 1'b1;  wr_cycle[10850] = 1'b0;  addr_rom[10850]='h0000313c;  wr_data_rom[10850]='h00000000;
    rd_cycle[10851] = 1'b0;  wr_cycle[10851] = 1'b1;  addr_rom[10851]='h0000090c;  wr_data_rom[10851]='h00003452;
    rd_cycle[10852] = 1'b1;  wr_cycle[10852] = 1'b0;  addr_rom[10852]='h0000150c;  wr_data_rom[10852]='h00000000;
    rd_cycle[10853] = 1'b1;  wr_cycle[10853] = 1'b0;  addr_rom[10853]='h0000370c;  wr_data_rom[10853]='h00000000;
    rd_cycle[10854] = 1'b1;  wr_cycle[10854] = 1'b0;  addr_rom[10854]='h00002964;  wr_data_rom[10854]='h00000000;
    rd_cycle[10855] = 1'b1;  wr_cycle[10855] = 1'b0;  addr_rom[10855]='h00002818;  wr_data_rom[10855]='h00000000;
    rd_cycle[10856] = 1'b0;  wr_cycle[10856] = 1'b1;  addr_rom[10856]='h00000b0c;  wr_data_rom[10856]='h000030e2;
    rd_cycle[10857] = 1'b1;  wr_cycle[10857] = 1'b0;  addr_rom[10857]='h000023e0;  wr_data_rom[10857]='h00000000;
    rd_cycle[10858] = 1'b1;  wr_cycle[10858] = 1'b0;  addr_rom[10858]='h00002310;  wr_data_rom[10858]='h00000000;
    rd_cycle[10859] = 1'b1;  wr_cycle[10859] = 1'b0;  addr_rom[10859]='h000021f0;  wr_data_rom[10859]='h00000000;
    rd_cycle[10860] = 1'b1;  wr_cycle[10860] = 1'b0;  addr_rom[10860]='h00003930;  wr_data_rom[10860]='h00000000;
    rd_cycle[10861] = 1'b1;  wr_cycle[10861] = 1'b0;  addr_rom[10861]='h00003bb0;  wr_data_rom[10861]='h00000000;
    rd_cycle[10862] = 1'b1;  wr_cycle[10862] = 1'b0;  addr_rom[10862]='h00002be0;  wr_data_rom[10862]='h00000000;
    rd_cycle[10863] = 1'b0;  wr_cycle[10863] = 1'b1;  addr_rom[10863]='h0000341c;  wr_data_rom[10863]='h00003c29;
    rd_cycle[10864] = 1'b1;  wr_cycle[10864] = 1'b0;  addr_rom[10864]='h00002fc4;  wr_data_rom[10864]='h00000000;
    rd_cycle[10865] = 1'b1;  wr_cycle[10865] = 1'b0;  addr_rom[10865]='h000024ec;  wr_data_rom[10865]='h00000000;
    rd_cycle[10866] = 1'b1;  wr_cycle[10866] = 1'b0;  addr_rom[10866]='h000007bc;  wr_data_rom[10866]='h00000000;
    rd_cycle[10867] = 1'b1;  wr_cycle[10867] = 1'b0;  addr_rom[10867]='h00003eec;  wr_data_rom[10867]='h00000000;
    rd_cycle[10868] = 1'b0;  wr_cycle[10868] = 1'b1;  addr_rom[10868]='h00001dbc;  wr_data_rom[10868]='h00003aab;
    rd_cycle[10869] = 1'b0;  wr_cycle[10869] = 1'b1;  addr_rom[10869]='h000032b0;  wr_data_rom[10869]='h00003cde;
    rd_cycle[10870] = 1'b0;  wr_cycle[10870] = 1'b1;  addr_rom[10870]='h00003dc4;  wr_data_rom[10870]='h000025fc;
    rd_cycle[10871] = 1'b0;  wr_cycle[10871] = 1'b1;  addr_rom[10871]='h000004fc;  wr_data_rom[10871]='h000030c9;
    rd_cycle[10872] = 1'b0;  wr_cycle[10872] = 1'b1;  addr_rom[10872]='h00001a94;  wr_data_rom[10872]='h00000b97;
    rd_cycle[10873] = 1'b0;  wr_cycle[10873] = 1'b1;  addr_rom[10873]='h00002bcc;  wr_data_rom[10873]='h0000343c;
    rd_cycle[10874] = 1'b1;  wr_cycle[10874] = 1'b0;  addr_rom[10874]='h00002160;  wr_data_rom[10874]='h00000000;
    rd_cycle[10875] = 1'b1;  wr_cycle[10875] = 1'b0;  addr_rom[10875]='h00001ec0;  wr_data_rom[10875]='h00000000;
    rd_cycle[10876] = 1'b1;  wr_cycle[10876] = 1'b0;  addr_rom[10876]='h00002de4;  wr_data_rom[10876]='h00000000;
    rd_cycle[10877] = 1'b1;  wr_cycle[10877] = 1'b0;  addr_rom[10877]='h00003408;  wr_data_rom[10877]='h00000000;
    rd_cycle[10878] = 1'b1;  wr_cycle[10878] = 1'b0;  addr_rom[10878]='h00000738;  wr_data_rom[10878]='h00000000;
    rd_cycle[10879] = 1'b1;  wr_cycle[10879] = 1'b0;  addr_rom[10879]='h00003994;  wr_data_rom[10879]='h00000000;
    rd_cycle[10880] = 1'b1;  wr_cycle[10880] = 1'b0;  addr_rom[10880]='h00000598;  wr_data_rom[10880]='h00000000;
    rd_cycle[10881] = 1'b1;  wr_cycle[10881] = 1'b0;  addr_rom[10881]='h00001db8;  wr_data_rom[10881]='h00000000;
    rd_cycle[10882] = 1'b0;  wr_cycle[10882] = 1'b1;  addr_rom[10882]='h00002d40;  wr_data_rom[10882]='h00001193;
    rd_cycle[10883] = 1'b1;  wr_cycle[10883] = 1'b0;  addr_rom[10883]='h00001fe8;  wr_data_rom[10883]='h00000000;
    rd_cycle[10884] = 1'b0;  wr_cycle[10884] = 1'b1;  addr_rom[10884]='h00001c8c;  wr_data_rom[10884]='h00000b79;
    rd_cycle[10885] = 1'b0;  wr_cycle[10885] = 1'b1;  addr_rom[10885]='h00002528;  wr_data_rom[10885]='h00001645;
    rd_cycle[10886] = 1'b1;  wr_cycle[10886] = 1'b0;  addr_rom[10886]='h00002274;  wr_data_rom[10886]='h00000000;
    rd_cycle[10887] = 1'b0;  wr_cycle[10887] = 1'b1;  addr_rom[10887]='h00002800;  wr_data_rom[10887]='h00001727;
    rd_cycle[10888] = 1'b1;  wr_cycle[10888] = 1'b0;  addr_rom[10888]='h00003660;  wr_data_rom[10888]='h00000000;
    rd_cycle[10889] = 1'b0;  wr_cycle[10889] = 1'b1;  addr_rom[10889]='h00001370;  wr_data_rom[10889]='h00001e39;
    rd_cycle[10890] = 1'b1;  wr_cycle[10890] = 1'b0;  addr_rom[10890]='h00002600;  wr_data_rom[10890]='h00000000;
    rd_cycle[10891] = 1'b1;  wr_cycle[10891] = 1'b0;  addr_rom[10891]='h000028a8;  wr_data_rom[10891]='h00000000;
    rd_cycle[10892] = 1'b0;  wr_cycle[10892] = 1'b1;  addr_rom[10892]='h00001f40;  wr_data_rom[10892]='h00000dbd;
    rd_cycle[10893] = 1'b1;  wr_cycle[10893] = 1'b0;  addr_rom[10893]='h00001de0;  wr_data_rom[10893]='h00000000;
    rd_cycle[10894] = 1'b0;  wr_cycle[10894] = 1'b1;  addr_rom[10894]='h00001ea0;  wr_data_rom[10894]='h000034a4;
    rd_cycle[10895] = 1'b1;  wr_cycle[10895] = 1'b0;  addr_rom[10895]='h00001874;  wr_data_rom[10895]='h00000000;
    rd_cycle[10896] = 1'b1;  wr_cycle[10896] = 1'b0;  addr_rom[10896]='h00002150;  wr_data_rom[10896]='h00000000;
    rd_cycle[10897] = 1'b1;  wr_cycle[10897] = 1'b0;  addr_rom[10897]='h00001720;  wr_data_rom[10897]='h00000000;
    rd_cycle[10898] = 1'b0;  wr_cycle[10898] = 1'b1;  addr_rom[10898]='h0000133c;  wr_data_rom[10898]='h000033c2;
    rd_cycle[10899] = 1'b0;  wr_cycle[10899] = 1'b1;  addr_rom[10899]='h000023d8;  wr_data_rom[10899]='h00003ee3;
    rd_cycle[10900] = 1'b0;  wr_cycle[10900] = 1'b1;  addr_rom[10900]='h00002b0c;  wr_data_rom[10900]='h00003a38;
    rd_cycle[10901] = 1'b0;  wr_cycle[10901] = 1'b1;  addr_rom[10901]='h00000b70;  wr_data_rom[10901]='h0000104a;
    rd_cycle[10902] = 1'b1;  wr_cycle[10902] = 1'b0;  addr_rom[10902]='h00002d34;  wr_data_rom[10902]='h00000000;
    rd_cycle[10903] = 1'b1;  wr_cycle[10903] = 1'b0;  addr_rom[10903]='h00001724;  wr_data_rom[10903]='h00000000;
    rd_cycle[10904] = 1'b1;  wr_cycle[10904] = 1'b0;  addr_rom[10904]='h0000301c;  wr_data_rom[10904]='h00000000;
    rd_cycle[10905] = 1'b0;  wr_cycle[10905] = 1'b1;  addr_rom[10905]='h0000316c;  wr_data_rom[10905]='h00000a4b;
    rd_cycle[10906] = 1'b0;  wr_cycle[10906] = 1'b1;  addr_rom[10906]='h000035b0;  wr_data_rom[10906]='h00003886;
    rd_cycle[10907] = 1'b1;  wr_cycle[10907] = 1'b0;  addr_rom[10907]='h00000f34;  wr_data_rom[10907]='h00000000;
    rd_cycle[10908] = 1'b1;  wr_cycle[10908] = 1'b0;  addr_rom[10908]='h000010d0;  wr_data_rom[10908]='h00000000;
    rd_cycle[10909] = 1'b1;  wr_cycle[10909] = 1'b0;  addr_rom[10909]='h00001040;  wr_data_rom[10909]='h00000000;
    rd_cycle[10910] = 1'b1;  wr_cycle[10910] = 1'b0;  addr_rom[10910]='h00001b48;  wr_data_rom[10910]='h00000000;
    rd_cycle[10911] = 1'b0;  wr_cycle[10911] = 1'b1;  addr_rom[10911]='h00000270;  wr_data_rom[10911]='h0000327b;
    rd_cycle[10912] = 1'b0;  wr_cycle[10912] = 1'b1;  addr_rom[10912]='h00000034;  wr_data_rom[10912]='h00003fdb;
    rd_cycle[10913] = 1'b1;  wr_cycle[10913] = 1'b0;  addr_rom[10913]='h00000da4;  wr_data_rom[10913]='h00000000;
    rd_cycle[10914] = 1'b1;  wr_cycle[10914] = 1'b0;  addr_rom[10914]='h000020f8;  wr_data_rom[10914]='h00000000;
    rd_cycle[10915] = 1'b1;  wr_cycle[10915] = 1'b0;  addr_rom[10915]='h0000330c;  wr_data_rom[10915]='h00000000;
    rd_cycle[10916] = 1'b1;  wr_cycle[10916] = 1'b0;  addr_rom[10916]='h00002624;  wr_data_rom[10916]='h00000000;
    rd_cycle[10917] = 1'b0;  wr_cycle[10917] = 1'b1;  addr_rom[10917]='h000039a0;  wr_data_rom[10917]='h0000094d;
    rd_cycle[10918] = 1'b1;  wr_cycle[10918] = 1'b0;  addr_rom[10918]='h0000269c;  wr_data_rom[10918]='h00000000;
    rd_cycle[10919] = 1'b0;  wr_cycle[10919] = 1'b1;  addr_rom[10919]='h00001d40;  wr_data_rom[10919]='h00001663;
    rd_cycle[10920] = 1'b0;  wr_cycle[10920] = 1'b1;  addr_rom[10920]='h00000f08;  wr_data_rom[10920]='h00002f14;
    rd_cycle[10921] = 1'b0;  wr_cycle[10921] = 1'b1;  addr_rom[10921]='h000011c0;  wr_data_rom[10921]='h00003f5d;
    rd_cycle[10922] = 1'b0;  wr_cycle[10922] = 1'b1;  addr_rom[10922]='h00003094;  wr_data_rom[10922]='h0000114a;
    rd_cycle[10923] = 1'b1;  wr_cycle[10923] = 1'b0;  addr_rom[10923]='h000021b4;  wr_data_rom[10923]='h00000000;
    rd_cycle[10924] = 1'b1;  wr_cycle[10924] = 1'b0;  addr_rom[10924]='h00001304;  wr_data_rom[10924]='h00000000;
    rd_cycle[10925] = 1'b0;  wr_cycle[10925] = 1'b1;  addr_rom[10925]='h00000870;  wr_data_rom[10925]='h00001874;
    rd_cycle[10926] = 1'b1;  wr_cycle[10926] = 1'b0;  addr_rom[10926]='h0000218c;  wr_data_rom[10926]='h00000000;
    rd_cycle[10927] = 1'b1;  wr_cycle[10927] = 1'b0;  addr_rom[10927]='h00003968;  wr_data_rom[10927]='h00000000;
    rd_cycle[10928] = 1'b1;  wr_cycle[10928] = 1'b0;  addr_rom[10928]='h000002b0;  wr_data_rom[10928]='h00000000;
    rd_cycle[10929] = 1'b1;  wr_cycle[10929] = 1'b0;  addr_rom[10929]='h0000218c;  wr_data_rom[10929]='h00000000;
    rd_cycle[10930] = 1'b0;  wr_cycle[10930] = 1'b1;  addr_rom[10930]='h00003518;  wr_data_rom[10930]='h0000227b;
    rd_cycle[10931] = 1'b1;  wr_cycle[10931] = 1'b0;  addr_rom[10931]='h00001f38;  wr_data_rom[10931]='h00000000;
    rd_cycle[10932] = 1'b0;  wr_cycle[10932] = 1'b1;  addr_rom[10932]='h00000544;  wr_data_rom[10932]='h000037ff;
    rd_cycle[10933] = 1'b0;  wr_cycle[10933] = 1'b1;  addr_rom[10933]='h000007bc;  wr_data_rom[10933]='h0000114e;
    rd_cycle[10934] = 1'b0;  wr_cycle[10934] = 1'b1;  addr_rom[10934]='h00003cc0;  wr_data_rom[10934]='h00002107;
    rd_cycle[10935] = 1'b0;  wr_cycle[10935] = 1'b1;  addr_rom[10935]='h000029f8;  wr_data_rom[10935]='h00002f47;
    rd_cycle[10936] = 1'b1;  wr_cycle[10936] = 1'b0;  addr_rom[10936]='h00003fc8;  wr_data_rom[10936]='h00000000;
    rd_cycle[10937] = 1'b0;  wr_cycle[10937] = 1'b1;  addr_rom[10937]='h00001ac8;  wr_data_rom[10937]='h00000189;
    rd_cycle[10938] = 1'b1;  wr_cycle[10938] = 1'b0;  addr_rom[10938]='h00001e50;  wr_data_rom[10938]='h00000000;
    rd_cycle[10939] = 1'b0;  wr_cycle[10939] = 1'b1;  addr_rom[10939]='h00000d20;  wr_data_rom[10939]='h00003cdb;
    rd_cycle[10940] = 1'b1;  wr_cycle[10940] = 1'b0;  addr_rom[10940]='h00000464;  wr_data_rom[10940]='h00000000;
    rd_cycle[10941] = 1'b1;  wr_cycle[10941] = 1'b0;  addr_rom[10941]='h00000bc8;  wr_data_rom[10941]='h00000000;
    rd_cycle[10942] = 1'b0;  wr_cycle[10942] = 1'b1;  addr_rom[10942]='h000033e4;  wr_data_rom[10942]='h00000af5;
    rd_cycle[10943] = 1'b1;  wr_cycle[10943] = 1'b0;  addr_rom[10943]='h00003eb4;  wr_data_rom[10943]='h00000000;
    rd_cycle[10944] = 1'b1;  wr_cycle[10944] = 1'b0;  addr_rom[10944]='h00001b50;  wr_data_rom[10944]='h00000000;
    rd_cycle[10945] = 1'b1;  wr_cycle[10945] = 1'b0;  addr_rom[10945]='h00000c78;  wr_data_rom[10945]='h00000000;
    rd_cycle[10946] = 1'b1;  wr_cycle[10946] = 1'b0;  addr_rom[10946]='h000029a0;  wr_data_rom[10946]='h00000000;
    rd_cycle[10947] = 1'b0;  wr_cycle[10947] = 1'b1;  addr_rom[10947]='h000018f4;  wr_data_rom[10947]='h00003967;
    rd_cycle[10948] = 1'b1;  wr_cycle[10948] = 1'b0;  addr_rom[10948]='h000017e0;  wr_data_rom[10948]='h00000000;
    rd_cycle[10949] = 1'b1;  wr_cycle[10949] = 1'b0;  addr_rom[10949]='h00003860;  wr_data_rom[10949]='h00000000;
    rd_cycle[10950] = 1'b1;  wr_cycle[10950] = 1'b0;  addr_rom[10950]='h00000c10;  wr_data_rom[10950]='h00000000;
    rd_cycle[10951] = 1'b0;  wr_cycle[10951] = 1'b1;  addr_rom[10951]='h00002118;  wr_data_rom[10951]='h00001c91;
    rd_cycle[10952] = 1'b0;  wr_cycle[10952] = 1'b1;  addr_rom[10952]='h000024a8;  wr_data_rom[10952]='h000032f4;
    rd_cycle[10953] = 1'b1;  wr_cycle[10953] = 1'b0;  addr_rom[10953]='h00001214;  wr_data_rom[10953]='h00000000;
    rd_cycle[10954] = 1'b1;  wr_cycle[10954] = 1'b0;  addr_rom[10954]='h0000225c;  wr_data_rom[10954]='h00000000;
    rd_cycle[10955] = 1'b1;  wr_cycle[10955] = 1'b0;  addr_rom[10955]='h000027a4;  wr_data_rom[10955]='h00000000;
    rd_cycle[10956] = 1'b1;  wr_cycle[10956] = 1'b0;  addr_rom[10956]='h00003464;  wr_data_rom[10956]='h00000000;
    rd_cycle[10957] = 1'b1;  wr_cycle[10957] = 1'b0;  addr_rom[10957]='h0000291c;  wr_data_rom[10957]='h00000000;
    rd_cycle[10958] = 1'b0;  wr_cycle[10958] = 1'b1;  addr_rom[10958]='h00002e68;  wr_data_rom[10958]='h00001604;
    rd_cycle[10959] = 1'b1;  wr_cycle[10959] = 1'b0;  addr_rom[10959]='h000039ac;  wr_data_rom[10959]='h00000000;
    rd_cycle[10960] = 1'b0;  wr_cycle[10960] = 1'b1;  addr_rom[10960]='h00002fe0;  wr_data_rom[10960]='h00001844;
    rd_cycle[10961] = 1'b1;  wr_cycle[10961] = 1'b0;  addr_rom[10961]='h00002904;  wr_data_rom[10961]='h00000000;
    rd_cycle[10962] = 1'b0;  wr_cycle[10962] = 1'b1;  addr_rom[10962]='h00001638;  wr_data_rom[10962]='h0000294d;
    rd_cycle[10963] = 1'b1;  wr_cycle[10963] = 1'b0;  addr_rom[10963]='h0000357c;  wr_data_rom[10963]='h00000000;
    rd_cycle[10964] = 1'b1;  wr_cycle[10964] = 1'b0;  addr_rom[10964]='h00002e0c;  wr_data_rom[10964]='h00000000;
    rd_cycle[10965] = 1'b1;  wr_cycle[10965] = 1'b0;  addr_rom[10965]='h00003ab0;  wr_data_rom[10965]='h00000000;
    rd_cycle[10966] = 1'b0;  wr_cycle[10966] = 1'b1;  addr_rom[10966]='h000035b4;  wr_data_rom[10966]='h00002083;
    rd_cycle[10967] = 1'b0;  wr_cycle[10967] = 1'b1;  addr_rom[10967]='h0000217c;  wr_data_rom[10967]='h00001d00;
    rd_cycle[10968] = 1'b0;  wr_cycle[10968] = 1'b1;  addr_rom[10968]='h00000930;  wr_data_rom[10968]='h000006fe;
    rd_cycle[10969] = 1'b1;  wr_cycle[10969] = 1'b0;  addr_rom[10969]='h00003d40;  wr_data_rom[10969]='h00000000;
    rd_cycle[10970] = 1'b0;  wr_cycle[10970] = 1'b1;  addr_rom[10970]='h00003e74;  wr_data_rom[10970]='h00003c88;
    rd_cycle[10971] = 1'b0;  wr_cycle[10971] = 1'b1;  addr_rom[10971]='h00002af0;  wr_data_rom[10971]='h00002bb8;
    rd_cycle[10972] = 1'b0;  wr_cycle[10972] = 1'b1;  addr_rom[10972]='h0000284c;  wr_data_rom[10972]='h000022eb;
    rd_cycle[10973] = 1'b1;  wr_cycle[10973] = 1'b0;  addr_rom[10973]='h000002bc;  wr_data_rom[10973]='h00000000;
    rd_cycle[10974] = 1'b0;  wr_cycle[10974] = 1'b1;  addr_rom[10974]='h0000292c;  wr_data_rom[10974]='h000026f5;
    rd_cycle[10975] = 1'b1;  wr_cycle[10975] = 1'b0;  addr_rom[10975]='h000037e0;  wr_data_rom[10975]='h00000000;
    rd_cycle[10976] = 1'b1;  wr_cycle[10976] = 1'b0;  addr_rom[10976]='h00003bb4;  wr_data_rom[10976]='h00000000;
    rd_cycle[10977] = 1'b0;  wr_cycle[10977] = 1'b1;  addr_rom[10977]='h000010ac;  wr_data_rom[10977]='h00003af5;
    rd_cycle[10978] = 1'b1;  wr_cycle[10978] = 1'b0;  addr_rom[10978]='h000001e8;  wr_data_rom[10978]='h00000000;
    rd_cycle[10979] = 1'b0;  wr_cycle[10979] = 1'b1;  addr_rom[10979]='h00002a10;  wr_data_rom[10979]='h00001812;
    rd_cycle[10980] = 1'b1;  wr_cycle[10980] = 1'b0;  addr_rom[10980]='h00003b48;  wr_data_rom[10980]='h00000000;
    rd_cycle[10981] = 1'b0;  wr_cycle[10981] = 1'b1;  addr_rom[10981]='h00002340;  wr_data_rom[10981]='h00001dd6;
    rd_cycle[10982] = 1'b0;  wr_cycle[10982] = 1'b1;  addr_rom[10982]='h00002580;  wr_data_rom[10982]='h00000318;
    rd_cycle[10983] = 1'b1;  wr_cycle[10983] = 1'b0;  addr_rom[10983]='h00002850;  wr_data_rom[10983]='h00000000;
    rd_cycle[10984] = 1'b0;  wr_cycle[10984] = 1'b1;  addr_rom[10984]='h000014a4;  wr_data_rom[10984]='h00002c44;
    rd_cycle[10985] = 1'b1;  wr_cycle[10985] = 1'b0;  addr_rom[10985]='h00001f98;  wr_data_rom[10985]='h00000000;
    rd_cycle[10986] = 1'b1;  wr_cycle[10986] = 1'b0;  addr_rom[10986]='h00000b40;  wr_data_rom[10986]='h00000000;
    rd_cycle[10987] = 1'b1;  wr_cycle[10987] = 1'b0;  addr_rom[10987]='h00002c10;  wr_data_rom[10987]='h00000000;
    rd_cycle[10988] = 1'b1;  wr_cycle[10988] = 1'b0;  addr_rom[10988]='h00000040;  wr_data_rom[10988]='h00000000;
    rd_cycle[10989] = 1'b0;  wr_cycle[10989] = 1'b1;  addr_rom[10989]='h00003f40;  wr_data_rom[10989]='h00003a25;
    rd_cycle[10990] = 1'b1;  wr_cycle[10990] = 1'b0;  addr_rom[10990]='h00002cac;  wr_data_rom[10990]='h00000000;
    rd_cycle[10991] = 1'b0;  wr_cycle[10991] = 1'b1;  addr_rom[10991]='h000037e0;  wr_data_rom[10991]='h00002de4;
    rd_cycle[10992] = 1'b1;  wr_cycle[10992] = 1'b0;  addr_rom[10992]='h00002d48;  wr_data_rom[10992]='h00000000;
    rd_cycle[10993] = 1'b0;  wr_cycle[10993] = 1'b1;  addr_rom[10993]='h00002024;  wr_data_rom[10993]='h00003e84;
    rd_cycle[10994] = 1'b1;  wr_cycle[10994] = 1'b0;  addr_rom[10994]='h00000584;  wr_data_rom[10994]='h00000000;
    rd_cycle[10995] = 1'b0;  wr_cycle[10995] = 1'b1;  addr_rom[10995]='h00003eac;  wr_data_rom[10995]='h00001f75;
    rd_cycle[10996] = 1'b0;  wr_cycle[10996] = 1'b1;  addr_rom[10996]='h00003480;  wr_data_rom[10996]='h000006cd;
    rd_cycle[10997] = 1'b1;  wr_cycle[10997] = 1'b0;  addr_rom[10997]='h00000f78;  wr_data_rom[10997]='h00000000;
    rd_cycle[10998] = 1'b1;  wr_cycle[10998] = 1'b0;  addr_rom[10998]='h00003218;  wr_data_rom[10998]='h00000000;
    rd_cycle[10999] = 1'b0;  wr_cycle[10999] = 1'b1;  addr_rom[10999]='h00003e58;  wr_data_rom[10999]='h000037b1;
    rd_cycle[11000] = 1'b1;  wr_cycle[11000] = 1'b0;  addr_rom[11000]='h000013dc;  wr_data_rom[11000]='h00000000;
    rd_cycle[11001] = 1'b0;  wr_cycle[11001] = 1'b1;  addr_rom[11001]='h00000f04;  wr_data_rom[11001]='h00002dfe;
    rd_cycle[11002] = 1'b1;  wr_cycle[11002] = 1'b0;  addr_rom[11002]='h000030f8;  wr_data_rom[11002]='h00000000;
    rd_cycle[11003] = 1'b1;  wr_cycle[11003] = 1'b0;  addr_rom[11003]='h00002e84;  wr_data_rom[11003]='h00000000;
    rd_cycle[11004] = 1'b0;  wr_cycle[11004] = 1'b1;  addr_rom[11004]='h00001af0;  wr_data_rom[11004]='h00002e7d;
    rd_cycle[11005] = 1'b1;  wr_cycle[11005] = 1'b0;  addr_rom[11005]='h00002b9c;  wr_data_rom[11005]='h00000000;
    rd_cycle[11006] = 1'b1;  wr_cycle[11006] = 1'b0;  addr_rom[11006]='h0000019c;  wr_data_rom[11006]='h00000000;
    rd_cycle[11007] = 1'b0;  wr_cycle[11007] = 1'b1;  addr_rom[11007]='h00002c6c;  wr_data_rom[11007]='h00002ee6;
    rd_cycle[11008] = 1'b1;  wr_cycle[11008] = 1'b0;  addr_rom[11008]='h000034b0;  wr_data_rom[11008]='h00000000;
    rd_cycle[11009] = 1'b1;  wr_cycle[11009] = 1'b0;  addr_rom[11009]='h00001b1c;  wr_data_rom[11009]='h00000000;
    rd_cycle[11010] = 1'b1;  wr_cycle[11010] = 1'b0;  addr_rom[11010]='h00001e5c;  wr_data_rom[11010]='h00000000;
    rd_cycle[11011] = 1'b0;  wr_cycle[11011] = 1'b1;  addr_rom[11011]='h00000420;  wr_data_rom[11011]='h00003f5d;
    rd_cycle[11012] = 1'b0;  wr_cycle[11012] = 1'b1;  addr_rom[11012]='h00002f10;  wr_data_rom[11012]='h00003d1a;
    rd_cycle[11013] = 1'b1;  wr_cycle[11013] = 1'b0;  addr_rom[11013]='h000010a8;  wr_data_rom[11013]='h00000000;
    rd_cycle[11014] = 1'b1;  wr_cycle[11014] = 1'b0;  addr_rom[11014]='h00000b18;  wr_data_rom[11014]='h00000000;
    rd_cycle[11015] = 1'b1;  wr_cycle[11015] = 1'b0;  addr_rom[11015]='h000028d0;  wr_data_rom[11015]='h00000000;
    rd_cycle[11016] = 1'b1;  wr_cycle[11016] = 1'b0;  addr_rom[11016]='h0000353c;  wr_data_rom[11016]='h00000000;
    rd_cycle[11017] = 1'b1;  wr_cycle[11017] = 1'b0;  addr_rom[11017]='h00002bac;  wr_data_rom[11017]='h00000000;
    rd_cycle[11018] = 1'b0;  wr_cycle[11018] = 1'b1;  addr_rom[11018]='h00001f50;  wr_data_rom[11018]='h00003d91;
    rd_cycle[11019] = 1'b1;  wr_cycle[11019] = 1'b0;  addr_rom[11019]='h0000236c;  wr_data_rom[11019]='h00000000;
    rd_cycle[11020] = 1'b0;  wr_cycle[11020] = 1'b1;  addr_rom[11020]='h00002284;  wr_data_rom[11020]='h00003ec5;
    rd_cycle[11021] = 1'b0;  wr_cycle[11021] = 1'b1;  addr_rom[11021]='h00003d94;  wr_data_rom[11021]='h00002928;
    rd_cycle[11022] = 1'b0;  wr_cycle[11022] = 1'b1;  addr_rom[11022]='h000039bc;  wr_data_rom[11022]='h00000e67;
    rd_cycle[11023] = 1'b1;  wr_cycle[11023] = 1'b0;  addr_rom[11023]='h00003e08;  wr_data_rom[11023]='h00000000;
    rd_cycle[11024] = 1'b0;  wr_cycle[11024] = 1'b1;  addr_rom[11024]='h00000de4;  wr_data_rom[11024]='h00003757;
    rd_cycle[11025] = 1'b1;  wr_cycle[11025] = 1'b0;  addr_rom[11025]='h00000fb4;  wr_data_rom[11025]='h00000000;
    rd_cycle[11026] = 1'b1;  wr_cycle[11026] = 1'b0;  addr_rom[11026]='h0000315c;  wr_data_rom[11026]='h00000000;
    rd_cycle[11027] = 1'b0;  wr_cycle[11027] = 1'b1;  addr_rom[11027]='h00000284;  wr_data_rom[11027]='h000015b8;
    rd_cycle[11028] = 1'b1;  wr_cycle[11028] = 1'b0;  addr_rom[11028]='h000028fc;  wr_data_rom[11028]='h00000000;
    rd_cycle[11029] = 1'b0;  wr_cycle[11029] = 1'b1;  addr_rom[11029]='h00003bc0;  wr_data_rom[11029]='h00000286;
    rd_cycle[11030] = 1'b0;  wr_cycle[11030] = 1'b1;  addr_rom[11030]='h00000a40;  wr_data_rom[11030]='h0000310c;
    rd_cycle[11031] = 1'b1;  wr_cycle[11031] = 1'b0;  addr_rom[11031]='h00001b5c;  wr_data_rom[11031]='h00000000;
    rd_cycle[11032] = 1'b1;  wr_cycle[11032] = 1'b0;  addr_rom[11032]='h00003130;  wr_data_rom[11032]='h00000000;
    rd_cycle[11033] = 1'b1;  wr_cycle[11033] = 1'b0;  addr_rom[11033]='h00002ba0;  wr_data_rom[11033]='h00000000;
    rd_cycle[11034] = 1'b1;  wr_cycle[11034] = 1'b0;  addr_rom[11034]='h000002b8;  wr_data_rom[11034]='h00000000;
    rd_cycle[11035] = 1'b1;  wr_cycle[11035] = 1'b0;  addr_rom[11035]='h00002e8c;  wr_data_rom[11035]='h00000000;
    rd_cycle[11036] = 1'b0;  wr_cycle[11036] = 1'b1;  addr_rom[11036]='h0000214c;  wr_data_rom[11036]='h00001adc;
    rd_cycle[11037] = 1'b0;  wr_cycle[11037] = 1'b1;  addr_rom[11037]='h00001494;  wr_data_rom[11037]='h000011c5;
    rd_cycle[11038] = 1'b1;  wr_cycle[11038] = 1'b0;  addr_rom[11038]='h00000ff0;  wr_data_rom[11038]='h00000000;
    rd_cycle[11039] = 1'b0;  wr_cycle[11039] = 1'b1;  addr_rom[11039]='h0000054c;  wr_data_rom[11039]='h00002c0b;
    rd_cycle[11040] = 1'b0;  wr_cycle[11040] = 1'b1;  addr_rom[11040]='h00001afc;  wr_data_rom[11040]='h00000e41;
    rd_cycle[11041] = 1'b1;  wr_cycle[11041] = 1'b0;  addr_rom[11041]='h000016c0;  wr_data_rom[11041]='h00000000;
    rd_cycle[11042] = 1'b1;  wr_cycle[11042] = 1'b0;  addr_rom[11042]='h00000fdc;  wr_data_rom[11042]='h00000000;
    rd_cycle[11043] = 1'b0;  wr_cycle[11043] = 1'b1;  addr_rom[11043]='h000000a8;  wr_data_rom[11043]='h00002c87;
    rd_cycle[11044] = 1'b1;  wr_cycle[11044] = 1'b0;  addr_rom[11044]='h00003e50;  wr_data_rom[11044]='h00000000;
    rd_cycle[11045] = 1'b0;  wr_cycle[11045] = 1'b1;  addr_rom[11045]='h00000444;  wr_data_rom[11045]='h000023b8;
    rd_cycle[11046] = 1'b0;  wr_cycle[11046] = 1'b1;  addr_rom[11046]='h00003084;  wr_data_rom[11046]='h00000fa8;
    rd_cycle[11047] = 1'b0;  wr_cycle[11047] = 1'b1;  addr_rom[11047]='h00000300;  wr_data_rom[11047]='h00001bf5;
    rd_cycle[11048] = 1'b0;  wr_cycle[11048] = 1'b1;  addr_rom[11048]='h00000f88;  wr_data_rom[11048]='h000002f1;
    rd_cycle[11049] = 1'b0;  wr_cycle[11049] = 1'b1;  addr_rom[11049]='h000029a8;  wr_data_rom[11049]='h00003b94;
    rd_cycle[11050] = 1'b1;  wr_cycle[11050] = 1'b0;  addr_rom[11050]='h00003734;  wr_data_rom[11050]='h00000000;
    rd_cycle[11051] = 1'b0;  wr_cycle[11051] = 1'b1;  addr_rom[11051]='h00001be8;  wr_data_rom[11051]='h000001e4;
    rd_cycle[11052] = 1'b1;  wr_cycle[11052] = 1'b0;  addr_rom[11052]='h000035ec;  wr_data_rom[11052]='h00000000;
    rd_cycle[11053] = 1'b0;  wr_cycle[11053] = 1'b1;  addr_rom[11053]='h000006f0;  wr_data_rom[11053]='h000009a0;
    rd_cycle[11054] = 1'b1;  wr_cycle[11054] = 1'b0;  addr_rom[11054]='h00002698;  wr_data_rom[11054]='h00000000;
    rd_cycle[11055] = 1'b1;  wr_cycle[11055] = 1'b0;  addr_rom[11055]='h00002bb8;  wr_data_rom[11055]='h00000000;
    rd_cycle[11056] = 1'b0;  wr_cycle[11056] = 1'b1;  addr_rom[11056]='h00002170;  wr_data_rom[11056]='h000022b7;
    rd_cycle[11057] = 1'b0;  wr_cycle[11057] = 1'b1;  addr_rom[11057]='h00002244;  wr_data_rom[11057]='h000025a5;
    rd_cycle[11058] = 1'b1;  wr_cycle[11058] = 1'b0;  addr_rom[11058]='h0000058c;  wr_data_rom[11058]='h00000000;
    rd_cycle[11059] = 1'b0;  wr_cycle[11059] = 1'b1;  addr_rom[11059]='h00000fd8;  wr_data_rom[11059]='h00003526;
    rd_cycle[11060] = 1'b1;  wr_cycle[11060] = 1'b0;  addr_rom[11060]='h00000b80;  wr_data_rom[11060]='h00000000;
    rd_cycle[11061] = 1'b0;  wr_cycle[11061] = 1'b1;  addr_rom[11061]='h000013dc;  wr_data_rom[11061]='h000034ed;
    rd_cycle[11062] = 1'b0;  wr_cycle[11062] = 1'b1;  addr_rom[11062]='h000027b4;  wr_data_rom[11062]='h0000154a;
    rd_cycle[11063] = 1'b0;  wr_cycle[11063] = 1'b1;  addr_rom[11063]='h000015c4;  wr_data_rom[11063]='h000035ce;
    rd_cycle[11064] = 1'b1;  wr_cycle[11064] = 1'b0;  addr_rom[11064]='h00000200;  wr_data_rom[11064]='h00000000;
    rd_cycle[11065] = 1'b0;  wr_cycle[11065] = 1'b1;  addr_rom[11065]='h00000a50;  wr_data_rom[11065]='h000003b1;
    rd_cycle[11066] = 1'b0;  wr_cycle[11066] = 1'b1;  addr_rom[11066]='h00001648;  wr_data_rom[11066]='h00001480;
    rd_cycle[11067] = 1'b0;  wr_cycle[11067] = 1'b1;  addr_rom[11067]='h00001cb4;  wr_data_rom[11067]='h00002cbd;
    rd_cycle[11068] = 1'b1;  wr_cycle[11068] = 1'b0;  addr_rom[11068]='h00003c00;  wr_data_rom[11068]='h00000000;
    rd_cycle[11069] = 1'b1;  wr_cycle[11069] = 1'b0;  addr_rom[11069]='h0000267c;  wr_data_rom[11069]='h00000000;
    rd_cycle[11070] = 1'b1;  wr_cycle[11070] = 1'b0;  addr_rom[11070]='h000032d8;  wr_data_rom[11070]='h00000000;
    rd_cycle[11071] = 1'b1;  wr_cycle[11071] = 1'b0;  addr_rom[11071]='h00001b54;  wr_data_rom[11071]='h00000000;
    rd_cycle[11072] = 1'b1;  wr_cycle[11072] = 1'b0;  addr_rom[11072]='h00002310;  wr_data_rom[11072]='h00000000;
    rd_cycle[11073] = 1'b1;  wr_cycle[11073] = 1'b0;  addr_rom[11073]='h00003a44;  wr_data_rom[11073]='h00000000;
    rd_cycle[11074] = 1'b1;  wr_cycle[11074] = 1'b0;  addr_rom[11074]='h000013e8;  wr_data_rom[11074]='h00000000;
    rd_cycle[11075] = 1'b0;  wr_cycle[11075] = 1'b1;  addr_rom[11075]='h000038d0;  wr_data_rom[11075]='h00002373;
    rd_cycle[11076] = 1'b1;  wr_cycle[11076] = 1'b0;  addr_rom[11076]='h000021ac;  wr_data_rom[11076]='h00000000;
    rd_cycle[11077] = 1'b0;  wr_cycle[11077] = 1'b1;  addr_rom[11077]='h00000410;  wr_data_rom[11077]='h00000b0c;
    rd_cycle[11078] = 1'b0;  wr_cycle[11078] = 1'b1;  addr_rom[11078]='h000019e4;  wr_data_rom[11078]='h00002226;
    rd_cycle[11079] = 1'b1;  wr_cycle[11079] = 1'b0;  addr_rom[11079]='h00003b6c;  wr_data_rom[11079]='h00000000;
    rd_cycle[11080] = 1'b1;  wr_cycle[11080] = 1'b0;  addr_rom[11080]='h00003380;  wr_data_rom[11080]='h00000000;
    rd_cycle[11081] = 1'b1;  wr_cycle[11081] = 1'b0;  addr_rom[11081]='h000025c4;  wr_data_rom[11081]='h00000000;
    rd_cycle[11082] = 1'b0;  wr_cycle[11082] = 1'b1;  addr_rom[11082]='h00002dcc;  wr_data_rom[11082]='h00003c0c;
    rd_cycle[11083] = 1'b0;  wr_cycle[11083] = 1'b1;  addr_rom[11083]='h00001c44;  wr_data_rom[11083]='h00000ee1;
    rd_cycle[11084] = 1'b1;  wr_cycle[11084] = 1'b0;  addr_rom[11084]='h0000101c;  wr_data_rom[11084]='h00000000;
    rd_cycle[11085] = 1'b0;  wr_cycle[11085] = 1'b1;  addr_rom[11085]='h00002528;  wr_data_rom[11085]='h00001e56;
    rd_cycle[11086] = 1'b1;  wr_cycle[11086] = 1'b0;  addr_rom[11086]='h0000181c;  wr_data_rom[11086]='h00000000;
    rd_cycle[11087] = 1'b1;  wr_cycle[11087] = 1'b0;  addr_rom[11087]='h00000c80;  wr_data_rom[11087]='h00000000;
    rd_cycle[11088] = 1'b0;  wr_cycle[11088] = 1'b1;  addr_rom[11088]='h00000238;  wr_data_rom[11088]='h000000b0;
    rd_cycle[11089] = 1'b1;  wr_cycle[11089] = 1'b0;  addr_rom[11089]='h000032f0;  wr_data_rom[11089]='h00000000;
    rd_cycle[11090] = 1'b0;  wr_cycle[11090] = 1'b1;  addr_rom[11090]='h00003358;  wr_data_rom[11090]='h000011e9;
    rd_cycle[11091] = 1'b1;  wr_cycle[11091] = 1'b0;  addr_rom[11091]='h000007c8;  wr_data_rom[11091]='h00000000;
    rd_cycle[11092] = 1'b1;  wr_cycle[11092] = 1'b0;  addr_rom[11092]='h00002990;  wr_data_rom[11092]='h00000000;
    rd_cycle[11093] = 1'b1;  wr_cycle[11093] = 1'b0;  addr_rom[11093]='h0000143c;  wr_data_rom[11093]='h00000000;
    rd_cycle[11094] = 1'b0;  wr_cycle[11094] = 1'b1;  addr_rom[11094]='h00001120;  wr_data_rom[11094]='h00003091;
    rd_cycle[11095] = 1'b0;  wr_cycle[11095] = 1'b1;  addr_rom[11095]='h00002544;  wr_data_rom[11095]='h00003d73;
    rd_cycle[11096] = 1'b1;  wr_cycle[11096] = 1'b0;  addr_rom[11096]='h00000e18;  wr_data_rom[11096]='h00000000;
    rd_cycle[11097] = 1'b0;  wr_cycle[11097] = 1'b1;  addr_rom[11097]='h00001cc8;  wr_data_rom[11097]='h00003a1f;
    rd_cycle[11098] = 1'b1;  wr_cycle[11098] = 1'b0;  addr_rom[11098]='h00001b4c;  wr_data_rom[11098]='h00000000;
    rd_cycle[11099] = 1'b0;  wr_cycle[11099] = 1'b1;  addr_rom[11099]='h00002a4c;  wr_data_rom[11099]='h00002c90;
    rd_cycle[11100] = 1'b1;  wr_cycle[11100] = 1'b0;  addr_rom[11100]='h00002638;  wr_data_rom[11100]='h00000000;
    rd_cycle[11101] = 1'b1;  wr_cycle[11101] = 1'b0;  addr_rom[11101]='h00002274;  wr_data_rom[11101]='h00000000;
    rd_cycle[11102] = 1'b1;  wr_cycle[11102] = 1'b0;  addr_rom[11102]='h0000288c;  wr_data_rom[11102]='h00000000;
    rd_cycle[11103] = 1'b0;  wr_cycle[11103] = 1'b1;  addr_rom[11103]='h0000169c;  wr_data_rom[11103]='h00001b12;
    rd_cycle[11104] = 1'b0;  wr_cycle[11104] = 1'b1;  addr_rom[11104]='h00002ab8;  wr_data_rom[11104]='h00003305;
    rd_cycle[11105] = 1'b0;  wr_cycle[11105] = 1'b1;  addr_rom[11105]='h00000990;  wr_data_rom[11105]='h00003cbc;
    rd_cycle[11106] = 1'b1;  wr_cycle[11106] = 1'b0;  addr_rom[11106]='h000009e4;  wr_data_rom[11106]='h00000000;
    rd_cycle[11107] = 1'b0;  wr_cycle[11107] = 1'b1;  addr_rom[11107]='h0000053c;  wr_data_rom[11107]='h000007f4;
    rd_cycle[11108] = 1'b1;  wr_cycle[11108] = 1'b0;  addr_rom[11108]='h00002388;  wr_data_rom[11108]='h00000000;
    rd_cycle[11109] = 1'b1;  wr_cycle[11109] = 1'b0;  addr_rom[11109]='h00001fd4;  wr_data_rom[11109]='h00000000;
    rd_cycle[11110] = 1'b0;  wr_cycle[11110] = 1'b1;  addr_rom[11110]='h00003a0c;  wr_data_rom[11110]='h0000144f;
    rd_cycle[11111] = 1'b1;  wr_cycle[11111] = 1'b0;  addr_rom[11111]='h000016e8;  wr_data_rom[11111]='h00000000;
    rd_cycle[11112] = 1'b0;  wr_cycle[11112] = 1'b1;  addr_rom[11112]='h00001b58;  wr_data_rom[11112]='h00003d9b;
    rd_cycle[11113] = 1'b1;  wr_cycle[11113] = 1'b0;  addr_rom[11113]='h000010fc;  wr_data_rom[11113]='h00000000;
    rd_cycle[11114] = 1'b1;  wr_cycle[11114] = 1'b0;  addr_rom[11114]='h0000327c;  wr_data_rom[11114]='h00000000;
    rd_cycle[11115] = 1'b0;  wr_cycle[11115] = 1'b1;  addr_rom[11115]='h00000e1c;  wr_data_rom[11115]='h000028bd;
    rd_cycle[11116] = 1'b1;  wr_cycle[11116] = 1'b0;  addr_rom[11116]='h000000c0;  wr_data_rom[11116]='h00000000;
    rd_cycle[11117] = 1'b1;  wr_cycle[11117] = 1'b0;  addr_rom[11117]='h00001138;  wr_data_rom[11117]='h00000000;
    rd_cycle[11118] = 1'b1;  wr_cycle[11118] = 1'b0;  addr_rom[11118]='h00000768;  wr_data_rom[11118]='h00000000;
    rd_cycle[11119] = 1'b0;  wr_cycle[11119] = 1'b1;  addr_rom[11119]='h000012fc;  wr_data_rom[11119]='h0000313d;
    rd_cycle[11120] = 1'b0;  wr_cycle[11120] = 1'b1;  addr_rom[11120]='h00001ff8;  wr_data_rom[11120]='h000008d1;
    rd_cycle[11121] = 1'b0;  wr_cycle[11121] = 1'b1;  addr_rom[11121]='h00000be4;  wr_data_rom[11121]='h000038b0;
    rd_cycle[11122] = 1'b0;  wr_cycle[11122] = 1'b1;  addr_rom[11122]='h000022ec;  wr_data_rom[11122]='h00000d22;
    rd_cycle[11123] = 1'b1;  wr_cycle[11123] = 1'b0;  addr_rom[11123]='h00003f28;  wr_data_rom[11123]='h00000000;
    rd_cycle[11124] = 1'b1;  wr_cycle[11124] = 1'b0;  addr_rom[11124]='h00001cac;  wr_data_rom[11124]='h00000000;
    rd_cycle[11125] = 1'b0;  wr_cycle[11125] = 1'b1;  addr_rom[11125]='h00000f84;  wr_data_rom[11125]='h00000c42;
    rd_cycle[11126] = 1'b1;  wr_cycle[11126] = 1'b0;  addr_rom[11126]='h00003104;  wr_data_rom[11126]='h00000000;
    rd_cycle[11127] = 1'b0;  wr_cycle[11127] = 1'b1;  addr_rom[11127]='h000000f4;  wr_data_rom[11127]='h0000026e;
    rd_cycle[11128] = 1'b0;  wr_cycle[11128] = 1'b1;  addr_rom[11128]='h00000edc;  wr_data_rom[11128]='h00001371;
    rd_cycle[11129] = 1'b0;  wr_cycle[11129] = 1'b1;  addr_rom[11129]='h00002538;  wr_data_rom[11129]='h0000073c;
    rd_cycle[11130] = 1'b1;  wr_cycle[11130] = 1'b0;  addr_rom[11130]='h0000303c;  wr_data_rom[11130]='h00000000;
    rd_cycle[11131] = 1'b1;  wr_cycle[11131] = 1'b0;  addr_rom[11131]='h000028b4;  wr_data_rom[11131]='h00000000;
    rd_cycle[11132] = 1'b0;  wr_cycle[11132] = 1'b1;  addr_rom[11132]='h000039ec;  wr_data_rom[11132]='h00003974;
    rd_cycle[11133] = 1'b0;  wr_cycle[11133] = 1'b1;  addr_rom[11133]='h000004b0;  wr_data_rom[11133]='h00002d1e;
    rd_cycle[11134] = 1'b1;  wr_cycle[11134] = 1'b0;  addr_rom[11134]='h00003a3c;  wr_data_rom[11134]='h00000000;
    rd_cycle[11135] = 1'b1;  wr_cycle[11135] = 1'b0;  addr_rom[11135]='h00001d54;  wr_data_rom[11135]='h00000000;
    rd_cycle[11136] = 1'b1;  wr_cycle[11136] = 1'b0;  addr_rom[11136]='h00003fd8;  wr_data_rom[11136]='h00000000;
    rd_cycle[11137] = 1'b1;  wr_cycle[11137] = 1'b0;  addr_rom[11137]='h00002318;  wr_data_rom[11137]='h00000000;
    rd_cycle[11138] = 1'b0;  wr_cycle[11138] = 1'b1;  addr_rom[11138]='h000022b0;  wr_data_rom[11138]='h00001dcf;
    rd_cycle[11139] = 1'b0;  wr_cycle[11139] = 1'b1;  addr_rom[11139]='h00002b94;  wr_data_rom[11139]='h0000290e;
    rd_cycle[11140] = 1'b0;  wr_cycle[11140] = 1'b1;  addr_rom[11140]='h000014ec;  wr_data_rom[11140]='h0000175a;
    rd_cycle[11141] = 1'b0;  wr_cycle[11141] = 1'b1;  addr_rom[11141]='h00000034;  wr_data_rom[11141]='h00002bac;
    rd_cycle[11142] = 1'b0;  wr_cycle[11142] = 1'b1;  addr_rom[11142]='h00000af8;  wr_data_rom[11142]='h000005b0;
    rd_cycle[11143] = 1'b1;  wr_cycle[11143] = 1'b0;  addr_rom[11143]='h00000bb4;  wr_data_rom[11143]='h00000000;
    rd_cycle[11144] = 1'b1;  wr_cycle[11144] = 1'b0;  addr_rom[11144]='h00002ff0;  wr_data_rom[11144]='h00000000;
    rd_cycle[11145] = 1'b1;  wr_cycle[11145] = 1'b0;  addr_rom[11145]='h00002eb8;  wr_data_rom[11145]='h00000000;
    rd_cycle[11146] = 1'b1;  wr_cycle[11146] = 1'b0;  addr_rom[11146]='h000015f8;  wr_data_rom[11146]='h00000000;
    rd_cycle[11147] = 1'b0;  wr_cycle[11147] = 1'b1;  addr_rom[11147]='h00000b14;  wr_data_rom[11147]='h000003f3;
    rd_cycle[11148] = 1'b1;  wr_cycle[11148] = 1'b0;  addr_rom[11148]='h00001c7c;  wr_data_rom[11148]='h00000000;
    rd_cycle[11149] = 1'b0;  wr_cycle[11149] = 1'b1;  addr_rom[11149]='h00002c6c;  wr_data_rom[11149]='h00003448;
    rd_cycle[11150] = 1'b0;  wr_cycle[11150] = 1'b1;  addr_rom[11150]='h00003190;  wr_data_rom[11150]='h000001b2;
    rd_cycle[11151] = 1'b0;  wr_cycle[11151] = 1'b1;  addr_rom[11151]='h00001ae0;  wr_data_rom[11151]='h00000025;
    rd_cycle[11152] = 1'b0;  wr_cycle[11152] = 1'b1;  addr_rom[11152]='h000028c0;  wr_data_rom[11152]='h00003401;
    rd_cycle[11153] = 1'b1;  wr_cycle[11153] = 1'b0;  addr_rom[11153]='h00000fe4;  wr_data_rom[11153]='h00000000;
    rd_cycle[11154] = 1'b1;  wr_cycle[11154] = 1'b0;  addr_rom[11154]='h00002274;  wr_data_rom[11154]='h00000000;
    rd_cycle[11155] = 1'b0;  wr_cycle[11155] = 1'b1;  addr_rom[11155]='h00002858;  wr_data_rom[11155]='h000018e0;
    rd_cycle[11156] = 1'b0;  wr_cycle[11156] = 1'b1;  addr_rom[11156]='h00001520;  wr_data_rom[11156]='h00002a54;
    rd_cycle[11157] = 1'b1;  wr_cycle[11157] = 1'b0;  addr_rom[11157]='h00000900;  wr_data_rom[11157]='h00000000;
    rd_cycle[11158] = 1'b1;  wr_cycle[11158] = 1'b0;  addr_rom[11158]='h00001bf8;  wr_data_rom[11158]='h00000000;
    rd_cycle[11159] = 1'b1;  wr_cycle[11159] = 1'b0;  addr_rom[11159]='h000037d8;  wr_data_rom[11159]='h00000000;
    rd_cycle[11160] = 1'b1;  wr_cycle[11160] = 1'b0;  addr_rom[11160]='h00002344;  wr_data_rom[11160]='h00000000;
    rd_cycle[11161] = 1'b0;  wr_cycle[11161] = 1'b1;  addr_rom[11161]='h00002954;  wr_data_rom[11161]='h000022c3;
    rd_cycle[11162] = 1'b1;  wr_cycle[11162] = 1'b0;  addr_rom[11162]='h000032a8;  wr_data_rom[11162]='h00000000;
    rd_cycle[11163] = 1'b1;  wr_cycle[11163] = 1'b0;  addr_rom[11163]='h000034e8;  wr_data_rom[11163]='h00000000;
    rd_cycle[11164] = 1'b0;  wr_cycle[11164] = 1'b1;  addr_rom[11164]='h00000288;  wr_data_rom[11164]='h00001d81;
    rd_cycle[11165] = 1'b1;  wr_cycle[11165] = 1'b0;  addr_rom[11165]='h00003eb0;  wr_data_rom[11165]='h00000000;
    rd_cycle[11166] = 1'b1;  wr_cycle[11166] = 1'b0;  addr_rom[11166]='h00000120;  wr_data_rom[11166]='h00000000;
    rd_cycle[11167] = 1'b1;  wr_cycle[11167] = 1'b0;  addr_rom[11167]='h00001a4c;  wr_data_rom[11167]='h00000000;
    rd_cycle[11168] = 1'b1;  wr_cycle[11168] = 1'b0;  addr_rom[11168]='h0000093c;  wr_data_rom[11168]='h00000000;
    rd_cycle[11169] = 1'b0;  wr_cycle[11169] = 1'b1;  addr_rom[11169]='h000001fc;  wr_data_rom[11169]='h000005f9;
    rd_cycle[11170] = 1'b1;  wr_cycle[11170] = 1'b0;  addr_rom[11170]='h00003510;  wr_data_rom[11170]='h00000000;
    rd_cycle[11171] = 1'b1;  wr_cycle[11171] = 1'b0;  addr_rom[11171]='h000018f0;  wr_data_rom[11171]='h00000000;
    rd_cycle[11172] = 1'b0;  wr_cycle[11172] = 1'b1;  addr_rom[11172]='h00002cbc;  wr_data_rom[11172]='h000004e1;
    rd_cycle[11173] = 1'b1;  wr_cycle[11173] = 1'b0;  addr_rom[11173]='h00003d14;  wr_data_rom[11173]='h00000000;
    rd_cycle[11174] = 1'b1;  wr_cycle[11174] = 1'b0;  addr_rom[11174]='h00001348;  wr_data_rom[11174]='h00000000;
    rd_cycle[11175] = 1'b1;  wr_cycle[11175] = 1'b0;  addr_rom[11175]='h000023b0;  wr_data_rom[11175]='h00000000;
    rd_cycle[11176] = 1'b1;  wr_cycle[11176] = 1'b0;  addr_rom[11176]='h00000e78;  wr_data_rom[11176]='h00000000;
    rd_cycle[11177] = 1'b0;  wr_cycle[11177] = 1'b1;  addr_rom[11177]='h00001f70;  wr_data_rom[11177]='h00001d2d;
    rd_cycle[11178] = 1'b1;  wr_cycle[11178] = 1'b0;  addr_rom[11178]='h00003d48;  wr_data_rom[11178]='h00000000;
    rd_cycle[11179] = 1'b1;  wr_cycle[11179] = 1'b0;  addr_rom[11179]='h000024c8;  wr_data_rom[11179]='h00000000;
    rd_cycle[11180] = 1'b1;  wr_cycle[11180] = 1'b0;  addr_rom[11180]='h000038a4;  wr_data_rom[11180]='h00000000;
    rd_cycle[11181] = 1'b1;  wr_cycle[11181] = 1'b0;  addr_rom[11181]='h000005c8;  wr_data_rom[11181]='h00000000;
    rd_cycle[11182] = 1'b0;  wr_cycle[11182] = 1'b1;  addr_rom[11182]='h00003d38;  wr_data_rom[11182]='h00003f10;
    rd_cycle[11183] = 1'b1;  wr_cycle[11183] = 1'b0;  addr_rom[11183]='h00000684;  wr_data_rom[11183]='h00000000;
    rd_cycle[11184] = 1'b1;  wr_cycle[11184] = 1'b0;  addr_rom[11184]='h00002130;  wr_data_rom[11184]='h00000000;
    rd_cycle[11185] = 1'b1;  wr_cycle[11185] = 1'b0;  addr_rom[11185]='h00000524;  wr_data_rom[11185]='h00000000;
    rd_cycle[11186] = 1'b1;  wr_cycle[11186] = 1'b0;  addr_rom[11186]='h00002214;  wr_data_rom[11186]='h00000000;
    rd_cycle[11187] = 1'b0;  wr_cycle[11187] = 1'b1;  addr_rom[11187]='h0000132c;  wr_data_rom[11187]='h00003ccd;
    rd_cycle[11188] = 1'b0;  wr_cycle[11188] = 1'b1;  addr_rom[11188]='h00003430;  wr_data_rom[11188]='h00003ef9;
    rd_cycle[11189] = 1'b1;  wr_cycle[11189] = 1'b0;  addr_rom[11189]='h00000d68;  wr_data_rom[11189]='h00000000;
    rd_cycle[11190] = 1'b1;  wr_cycle[11190] = 1'b0;  addr_rom[11190]='h00001bec;  wr_data_rom[11190]='h00000000;
    rd_cycle[11191] = 1'b1;  wr_cycle[11191] = 1'b0;  addr_rom[11191]='h00003664;  wr_data_rom[11191]='h00000000;
    rd_cycle[11192] = 1'b1;  wr_cycle[11192] = 1'b0;  addr_rom[11192]='h00003b40;  wr_data_rom[11192]='h00000000;
    rd_cycle[11193] = 1'b0;  wr_cycle[11193] = 1'b1;  addr_rom[11193]='h00000dfc;  wr_data_rom[11193]='h00002bfb;
    rd_cycle[11194] = 1'b1;  wr_cycle[11194] = 1'b0;  addr_rom[11194]='h0000253c;  wr_data_rom[11194]='h00000000;
    rd_cycle[11195] = 1'b0;  wr_cycle[11195] = 1'b1;  addr_rom[11195]='h00002588;  wr_data_rom[11195]='h000026b3;
    rd_cycle[11196] = 1'b1;  wr_cycle[11196] = 1'b0;  addr_rom[11196]='h00001b18;  wr_data_rom[11196]='h00000000;
    rd_cycle[11197] = 1'b0;  wr_cycle[11197] = 1'b1;  addr_rom[11197]='h0000325c;  wr_data_rom[11197]='h00003941;
    rd_cycle[11198] = 1'b1;  wr_cycle[11198] = 1'b0;  addr_rom[11198]='h000020fc;  wr_data_rom[11198]='h00000000;
    rd_cycle[11199] = 1'b0;  wr_cycle[11199] = 1'b1;  addr_rom[11199]='h00002100;  wr_data_rom[11199]='h00001d8b;
    rd_cycle[11200] = 1'b1;  wr_cycle[11200] = 1'b0;  addr_rom[11200]='h00000930;  wr_data_rom[11200]='h00000000;
    rd_cycle[11201] = 1'b1;  wr_cycle[11201] = 1'b0;  addr_rom[11201]='h0000289c;  wr_data_rom[11201]='h00000000;
    rd_cycle[11202] = 1'b1;  wr_cycle[11202] = 1'b0;  addr_rom[11202]='h000026dc;  wr_data_rom[11202]='h00000000;
    rd_cycle[11203] = 1'b1;  wr_cycle[11203] = 1'b0;  addr_rom[11203]='h00001a20;  wr_data_rom[11203]='h00000000;
    rd_cycle[11204] = 1'b0;  wr_cycle[11204] = 1'b1;  addr_rom[11204]='h00001d04;  wr_data_rom[11204]='h000017f7;
    rd_cycle[11205] = 1'b1;  wr_cycle[11205] = 1'b0;  addr_rom[11205]='h00001e9c;  wr_data_rom[11205]='h00000000;
    rd_cycle[11206] = 1'b0;  wr_cycle[11206] = 1'b1;  addr_rom[11206]='h00003138;  wr_data_rom[11206]='h00000443;
    rd_cycle[11207] = 1'b1;  wr_cycle[11207] = 1'b0;  addr_rom[11207]='h00000408;  wr_data_rom[11207]='h00000000;
    rd_cycle[11208] = 1'b0;  wr_cycle[11208] = 1'b1;  addr_rom[11208]='h00002db0;  wr_data_rom[11208]='h00002618;
    rd_cycle[11209] = 1'b1;  wr_cycle[11209] = 1'b0;  addr_rom[11209]='h0000070c;  wr_data_rom[11209]='h00000000;
    rd_cycle[11210] = 1'b1;  wr_cycle[11210] = 1'b0;  addr_rom[11210]='h00001560;  wr_data_rom[11210]='h00000000;
    rd_cycle[11211] = 1'b0;  wr_cycle[11211] = 1'b1;  addr_rom[11211]='h000030a0;  wr_data_rom[11211]='h00002f52;
    rd_cycle[11212] = 1'b1;  wr_cycle[11212] = 1'b0;  addr_rom[11212]='h000009e4;  wr_data_rom[11212]='h00000000;
    rd_cycle[11213] = 1'b0;  wr_cycle[11213] = 1'b1;  addr_rom[11213]='h000011d8;  wr_data_rom[11213]='h00000cd8;
    rd_cycle[11214] = 1'b0;  wr_cycle[11214] = 1'b1;  addr_rom[11214]='h000032f0;  wr_data_rom[11214]='h000017d7;
    rd_cycle[11215] = 1'b0;  wr_cycle[11215] = 1'b1;  addr_rom[11215]='h00002f3c;  wr_data_rom[11215]='h00002a08;
    rd_cycle[11216] = 1'b1;  wr_cycle[11216] = 1'b0;  addr_rom[11216]='h00003a90;  wr_data_rom[11216]='h00000000;
    rd_cycle[11217] = 1'b0;  wr_cycle[11217] = 1'b1;  addr_rom[11217]='h00003f64;  wr_data_rom[11217]='h00000a82;
    rd_cycle[11218] = 1'b1;  wr_cycle[11218] = 1'b0;  addr_rom[11218]='h0000192c;  wr_data_rom[11218]='h00000000;
    rd_cycle[11219] = 1'b0;  wr_cycle[11219] = 1'b1;  addr_rom[11219]='h00002054;  wr_data_rom[11219]='h0000271f;
    rd_cycle[11220] = 1'b1;  wr_cycle[11220] = 1'b0;  addr_rom[11220]='h00003e5c;  wr_data_rom[11220]='h00000000;
    rd_cycle[11221] = 1'b1;  wr_cycle[11221] = 1'b0;  addr_rom[11221]='h00001e70;  wr_data_rom[11221]='h00000000;
    rd_cycle[11222] = 1'b1;  wr_cycle[11222] = 1'b0;  addr_rom[11222]='h0000322c;  wr_data_rom[11222]='h00000000;
    rd_cycle[11223] = 1'b1;  wr_cycle[11223] = 1'b0;  addr_rom[11223]='h00000da4;  wr_data_rom[11223]='h00000000;
    rd_cycle[11224] = 1'b1;  wr_cycle[11224] = 1'b0;  addr_rom[11224]='h000036dc;  wr_data_rom[11224]='h00000000;
    rd_cycle[11225] = 1'b1;  wr_cycle[11225] = 1'b0;  addr_rom[11225]='h00000500;  wr_data_rom[11225]='h00000000;
    rd_cycle[11226] = 1'b1;  wr_cycle[11226] = 1'b0;  addr_rom[11226]='h00003118;  wr_data_rom[11226]='h00000000;
    rd_cycle[11227] = 1'b1;  wr_cycle[11227] = 1'b0;  addr_rom[11227]='h000004c0;  wr_data_rom[11227]='h00000000;
    rd_cycle[11228] = 1'b1;  wr_cycle[11228] = 1'b0;  addr_rom[11228]='h00002d2c;  wr_data_rom[11228]='h00000000;
    rd_cycle[11229] = 1'b1;  wr_cycle[11229] = 1'b0;  addr_rom[11229]='h00001dbc;  wr_data_rom[11229]='h00000000;
    rd_cycle[11230] = 1'b1;  wr_cycle[11230] = 1'b0;  addr_rom[11230]='h00001ecc;  wr_data_rom[11230]='h00000000;
    rd_cycle[11231] = 1'b1;  wr_cycle[11231] = 1'b0;  addr_rom[11231]='h00002ad0;  wr_data_rom[11231]='h00000000;
    rd_cycle[11232] = 1'b1;  wr_cycle[11232] = 1'b0;  addr_rom[11232]='h00000914;  wr_data_rom[11232]='h00000000;
    rd_cycle[11233] = 1'b1;  wr_cycle[11233] = 1'b0;  addr_rom[11233]='h000026d8;  wr_data_rom[11233]='h00000000;
    rd_cycle[11234] = 1'b1;  wr_cycle[11234] = 1'b0;  addr_rom[11234]='h0000323c;  wr_data_rom[11234]='h00000000;
    rd_cycle[11235] = 1'b1;  wr_cycle[11235] = 1'b0;  addr_rom[11235]='h0000351c;  wr_data_rom[11235]='h00000000;
    rd_cycle[11236] = 1'b0;  wr_cycle[11236] = 1'b1;  addr_rom[11236]='h00000a80;  wr_data_rom[11236]='h00003d3a;
    rd_cycle[11237] = 1'b1;  wr_cycle[11237] = 1'b0;  addr_rom[11237]='h000029a8;  wr_data_rom[11237]='h00000000;
    rd_cycle[11238] = 1'b0;  wr_cycle[11238] = 1'b1;  addr_rom[11238]='h00001390;  wr_data_rom[11238]='h00003000;
    rd_cycle[11239] = 1'b0;  wr_cycle[11239] = 1'b1;  addr_rom[11239]='h00001568;  wr_data_rom[11239]='h00003067;
    rd_cycle[11240] = 1'b1;  wr_cycle[11240] = 1'b0;  addr_rom[11240]='h00000c60;  wr_data_rom[11240]='h00000000;
    rd_cycle[11241] = 1'b0;  wr_cycle[11241] = 1'b1;  addr_rom[11241]='h00003fc0;  wr_data_rom[11241]='h000036c3;
    rd_cycle[11242] = 1'b1;  wr_cycle[11242] = 1'b0;  addr_rom[11242]='h00000f84;  wr_data_rom[11242]='h00000000;
    rd_cycle[11243] = 1'b0;  wr_cycle[11243] = 1'b1;  addr_rom[11243]='h00003410;  wr_data_rom[11243]='h00002df8;
    rd_cycle[11244] = 1'b1;  wr_cycle[11244] = 1'b0;  addr_rom[11244]='h00003390;  wr_data_rom[11244]='h00000000;
    rd_cycle[11245] = 1'b1;  wr_cycle[11245] = 1'b0;  addr_rom[11245]='h00001330;  wr_data_rom[11245]='h00000000;
    rd_cycle[11246] = 1'b1;  wr_cycle[11246] = 1'b0;  addr_rom[11246]='h00001ba4;  wr_data_rom[11246]='h00000000;
    rd_cycle[11247] = 1'b1;  wr_cycle[11247] = 1'b0;  addr_rom[11247]='h00000db8;  wr_data_rom[11247]='h00000000;
    rd_cycle[11248] = 1'b1;  wr_cycle[11248] = 1'b0;  addr_rom[11248]='h000013c8;  wr_data_rom[11248]='h00000000;
    rd_cycle[11249] = 1'b1;  wr_cycle[11249] = 1'b0;  addr_rom[11249]='h00003d88;  wr_data_rom[11249]='h00000000;
    rd_cycle[11250] = 1'b0;  wr_cycle[11250] = 1'b1;  addr_rom[11250]='h00000230;  wr_data_rom[11250]='h00001844;
    rd_cycle[11251] = 1'b0;  wr_cycle[11251] = 1'b1;  addr_rom[11251]='h00003438;  wr_data_rom[11251]='h0000290e;
    rd_cycle[11252] = 1'b0;  wr_cycle[11252] = 1'b1;  addr_rom[11252]='h000007ec;  wr_data_rom[11252]='h00003612;
    rd_cycle[11253] = 1'b0;  wr_cycle[11253] = 1'b1;  addr_rom[11253]='h000023c0;  wr_data_rom[11253]='h00003145;
    rd_cycle[11254] = 1'b0;  wr_cycle[11254] = 1'b1;  addr_rom[11254]='h00003f94;  wr_data_rom[11254]='h000008b1;
    rd_cycle[11255] = 1'b0;  wr_cycle[11255] = 1'b1;  addr_rom[11255]='h0000269c;  wr_data_rom[11255]='h00001916;
    rd_cycle[11256] = 1'b0;  wr_cycle[11256] = 1'b1;  addr_rom[11256]='h00000520;  wr_data_rom[11256]='h00002ed7;
    rd_cycle[11257] = 1'b1;  wr_cycle[11257] = 1'b0;  addr_rom[11257]='h00001298;  wr_data_rom[11257]='h00000000;
    rd_cycle[11258] = 1'b0;  wr_cycle[11258] = 1'b1;  addr_rom[11258]='h00002f70;  wr_data_rom[11258]='h00001d7c;
    rd_cycle[11259] = 1'b0;  wr_cycle[11259] = 1'b1;  addr_rom[11259]='h00000d7c;  wr_data_rom[11259]='h00002a6b;
    rd_cycle[11260] = 1'b1;  wr_cycle[11260] = 1'b0;  addr_rom[11260]='h00000144;  wr_data_rom[11260]='h00000000;
    rd_cycle[11261] = 1'b1;  wr_cycle[11261] = 1'b0;  addr_rom[11261]='h00002b20;  wr_data_rom[11261]='h00000000;
    rd_cycle[11262] = 1'b0;  wr_cycle[11262] = 1'b1;  addr_rom[11262]='h000000b0;  wr_data_rom[11262]='h00003c78;
    rd_cycle[11263] = 1'b1;  wr_cycle[11263] = 1'b0;  addr_rom[11263]='h000031b8;  wr_data_rom[11263]='h00000000;
    rd_cycle[11264] = 1'b1;  wr_cycle[11264] = 1'b0;  addr_rom[11264]='h0000273c;  wr_data_rom[11264]='h00000000;
    rd_cycle[11265] = 1'b1;  wr_cycle[11265] = 1'b0;  addr_rom[11265]='h000017d8;  wr_data_rom[11265]='h00000000;
    rd_cycle[11266] = 1'b1;  wr_cycle[11266] = 1'b0;  addr_rom[11266]='h0000249c;  wr_data_rom[11266]='h00000000;
    rd_cycle[11267] = 1'b0;  wr_cycle[11267] = 1'b1;  addr_rom[11267]='h00000ec4;  wr_data_rom[11267]='h00000c08;
    rd_cycle[11268] = 1'b1;  wr_cycle[11268] = 1'b0;  addr_rom[11268]='h00003190;  wr_data_rom[11268]='h00000000;
    rd_cycle[11269] = 1'b0;  wr_cycle[11269] = 1'b1;  addr_rom[11269]='h00002348;  wr_data_rom[11269]='h00003689;
    rd_cycle[11270] = 1'b1;  wr_cycle[11270] = 1'b0;  addr_rom[11270]='h00001450;  wr_data_rom[11270]='h00000000;
    rd_cycle[11271] = 1'b0;  wr_cycle[11271] = 1'b1;  addr_rom[11271]='h0000247c;  wr_data_rom[11271]='h00002f45;
    rd_cycle[11272] = 1'b0;  wr_cycle[11272] = 1'b1;  addr_rom[11272]='h00002ffc;  wr_data_rom[11272]='h000029f6;
    rd_cycle[11273] = 1'b1;  wr_cycle[11273] = 1'b0;  addr_rom[11273]='h000026a4;  wr_data_rom[11273]='h00000000;
    rd_cycle[11274] = 1'b0;  wr_cycle[11274] = 1'b1;  addr_rom[11274]='h00000090;  wr_data_rom[11274]='h00001895;
    rd_cycle[11275] = 1'b1;  wr_cycle[11275] = 1'b0;  addr_rom[11275]='h0000169c;  wr_data_rom[11275]='h00000000;
    rd_cycle[11276] = 1'b0;  wr_cycle[11276] = 1'b1;  addr_rom[11276]='h00001ff8;  wr_data_rom[11276]='h000019e4;
    rd_cycle[11277] = 1'b1;  wr_cycle[11277] = 1'b0;  addr_rom[11277]='h00001310;  wr_data_rom[11277]='h00000000;
    rd_cycle[11278] = 1'b1;  wr_cycle[11278] = 1'b0;  addr_rom[11278]='h00000110;  wr_data_rom[11278]='h00000000;
    rd_cycle[11279] = 1'b1;  wr_cycle[11279] = 1'b0;  addr_rom[11279]='h00000760;  wr_data_rom[11279]='h00000000;
    rd_cycle[11280] = 1'b0;  wr_cycle[11280] = 1'b1;  addr_rom[11280]='h00001028;  wr_data_rom[11280]='h00001c89;
    rd_cycle[11281] = 1'b1;  wr_cycle[11281] = 1'b0;  addr_rom[11281]='h00001480;  wr_data_rom[11281]='h00000000;
    rd_cycle[11282] = 1'b1;  wr_cycle[11282] = 1'b0;  addr_rom[11282]='h000025ac;  wr_data_rom[11282]='h00000000;
    rd_cycle[11283] = 1'b0;  wr_cycle[11283] = 1'b1;  addr_rom[11283]='h0000087c;  wr_data_rom[11283]='h000030e0;
    rd_cycle[11284] = 1'b1;  wr_cycle[11284] = 1'b0;  addr_rom[11284]='h00001e28;  wr_data_rom[11284]='h00000000;
    rd_cycle[11285] = 1'b1;  wr_cycle[11285] = 1'b0;  addr_rom[11285]='h00001e3c;  wr_data_rom[11285]='h00000000;
    rd_cycle[11286] = 1'b0;  wr_cycle[11286] = 1'b1;  addr_rom[11286]='h00000bac;  wr_data_rom[11286]='h00002ca4;
    rd_cycle[11287] = 1'b0;  wr_cycle[11287] = 1'b1;  addr_rom[11287]='h0000248c;  wr_data_rom[11287]='h00001bc7;
    rd_cycle[11288] = 1'b0;  wr_cycle[11288] = 1'b1;  addr_rom[11288]='h000020ac;  wr_data_rom[11288]='h0000261b;
    rd_cycle[11289] = 1'b1;  wr_cycle[11289] = 1'b0;  addr_rom[11289]='h00002d00;  wr_data_rom[11289]='h00000000;
    rd_cycle[11290] = 1'b1;  wr_cycle[11290] = 1'b0;  addr_rom[11290]='h00003234;  wr_data_rom[11290]='h00000000;
    rd_cycle[11291] = 1'b1;  wr_cycle[11291] = 1'b0;  addr_rom[11291]='h00000794;  wr_data_rom[11291]='h00000000;
    rd_cycle[11292] = 1'b0;  wr_cycle[11292] = 1'b1;  addr_rom[11292]='h000017e0;  wr_data_rom[11292]='h0000399c;
    rd_cycle[11293] = 1'b0;  wr_cycle[11293] = 1'b1;  addr_rom[11293]='h000022e8;  wr_data_rom[11293]='h00000c8f;
    rd_cycle[11294] = 1'b0;  wr_cycle[11294] = 1'b1;  addr_rom[11294]='h00000430;  wr_data_rom[11294]='h00003f4c;
    rd_cycle[11295] = 1'b1;  wr_cycle[11295] = 1'b0;  addr_rom[11295]='h00002578;  wr_data_rom[11295]='h00000000;
    rd_cycle[11296] = 1'b1;  wr_cycle[11296] = 1'b0;  addr_rom[11296]='h00001c58;  wr_data_rom[11296]='h00000000;
    rd_cycle[11297] = 1'b0;  wr_cycle[11297] = 1'b1;  addr_rom[11297]='h00002ec4;  wr_data_rom[11297]='h00001b76;
    rd_cycle[11298] = 1'b1;  wr_cycle[11298] = 1'b0;  addr_rom[11298]='h00000180;  wr_data_rom[11298]='h00000000;
    rd_cycle[11299] = 1'b1;  wr_cycle[11299] = 1'b0;  addr_rom[11299]='h00003c84;  wr_data_rom[11299]='h00000000;
    rd_cycle[11300] = 1'b1;  wr_cycle[11300] = 1'b0;  addr_rom[11300]='h000003cc;  wr_data_rom[11300]='h00000000;
    rd_cycle[11301] = 1'b1;  wr_cycle[11301] = 1'b0;  addr_rom[11301]='h00002a54;  wr_data_rom[11301]='h00000000;
    rd_cycle[11302] = 1'b1;  wr_cycle[11302] = 1'b0;  addr_rom[11302]='h000000e0;  wr_data_rom[11302]='h00000000;
    rd_cycle[11303] = 1'b0;  wr_cycle[11303] = 1'b1;  addr_rom[11303]='h00001290;  wr_data_rom[11303]='h00002683;
    rd_cycle[11304] = 1'b1;  wr_cycle[11304] = 1'b0;  addr_rom[11304]='h00002f98;  wr_data_rom[11304]='h00000000;
    rd_cycle[11305] = 1'b0;  wr_cycle[11305] = 1'b1;  addr_rom[11305]='h00003fe4;  wr_data_rom[11305]='h000035a5;
    rd_cycle[11306] = 1'b0;  wr_cycle[11306] = 1'b1;  addr_rom[11306]='h00000e70;  wr_data_rom[11306]='h000028f3;
    rd_cycle[11307] = 1'b1;  wr_cycle[11307] = 1'b0;  addr_rom[11307]='h00002124;  wr_data_rom[11307]='h00000000;
    rd_cycle[11308] = 1'b1;  wr_cycle[11308] = 1'b0;  addr_rom[11308]='h000018a4;  wr_data_rom[11308]='h00000000;
    rd_cycle[11309] = 1'b0;  wr_cycle[11309] = 1'b1;  addr_rom[11309]='h00003708;  wr_data_rom[11309]='h00000dcb;
    rd_cycle[11310] = 1'b1;  wr_cycle[11310] = 1'b0;  addr_rom[11310]='h0000114c;  wr_data_rom[11310]='h00000000;
    rd_cycle[11311] = 1'b0;  wr_cycle[11311] = 1'b1;  addr_rom[11311]='h00000400;  wr_data_rom[11311]='h00000540;
    rd_cycle[11312] = 1'b1;  wr_cycle[11312] = 1'b0;  addr_rom[11312]='h0000154c;  wr_data_rom[11312]='h00000000;
    rd_cycle[11313] = 1'b0;  wr_cycle[11313] = 1'b1;  addr_rom[11313]='h00001c48;  wr_data_rom[11313]='h0000206a;
    rd_cycle[11314] = 1'b1;  wr_cycle[11314] = 1'b0;  addr_rom[11314]='h00003d30;  wr_data_rom[11314]='h00000000;
    rd_cycle[11315] = 1'b1;  wr_cycle[11315] = 1'b0;  addr_rom[11315]='h000036d8;  wr_data_rom[11315]='h00000000;
    rd_cycle[11316] = 1'b0;  wr_cycle[11316] = 1'b1;  addr_rom[11316]='h00001744;  wr_data_rom[11316]='h000005e4;
    rd_cycle[11317] = 1'b0;  wr_cycle[11317] = 1'b1;  addr_rom[11317]='h000003e4;  wr_data_rom[11317]='h0000259f;
    rd_cycle[11318] = 1'b0;  wr_cycle[11318] = 1'b1;  addr_rom[11318]='h00000174;  wr_data_rom[11318]='h000023c8;
    rd_cycle[11319] = 1'b0;  wr_cycle[11319] = 1'b1;  addr_rom[11319]='h00003d08;  wr_data_rom[11319]='h0000336d;
    rd_cycle[11320] = 1'b0;  wr_cycle[11320] = 1'b1;  addr_rom[11320]='h00000be0;  wr_data_rom[11320]='h00000374;
    rd_cycle[11321] = 1'b0;  wr_cycle[11321] = 1'b1;  addr_rom[11321]='h00003120;  wr_data_rom[11321]='h00001b28;
    rd_cycle[11322] = 1'b1;  wr_cycle[11322] = 1'b0;  addr_rom[11322]='h00003dfc;  wr_data_rom[11322]='h00000000;
    rd_cycle[11323] = 1'b0;  wr_cycle[11323] = 1'b1;  addr_rom[11323]='h00003eac;  wr_data_rom[11323]='h00002a78;
    rd_cycle[11324] = 1'b1;  wr_cycle[11324] = 1'b0;  addr_rom[11324]='h000008e4;  wr_data_rom[11324]='h00000000;
    rd_cycle[11325] = 1'b1;  wr_cycle[11325] = 1'b0;  addr_rom[11325]='h000017e8;  wr_data_rom[11325]='h00000000;
    rd_cycle[11326] = 1'b1;  wr_cycle[11326] = 1'b0;  addr_rom[11326]='h00003a08;  wr_data_rom[11326]='h00000000;
    rd_cycle[11327] = 1'b1;  wr_cycle[11327] = 1'b0;  addr_rom[11327]='h00002ef0;  wr_data_rom[11327]='h00000000;
    rd_cycle[11328] = 1'b1;  wr_cycle[11328] = 1'b0;  addr_rom[11328]='h000015dc;  wr_data_rom[11328]='h00000000;
    rd_cycle[11329] = 1'b0;  wr_cycle[11329] = 1'b1;  addr_rom[11329]='h00001498;  wr_data_rom[11329]='h00000a37;
    rd_cycle[11330] = 1'b0;  wr_cycle[11330] = 1'b1;  addr_rom[11330]='h000018a8;  wr_data_rom[11330]='h00000c0a;
    rd_cycle[11331] = 1'b1;  wr_cycle[11331] = 1'b0;  addr_rom[11331]='h000024b8;  wr_data_rom[11331]='h00000000;
    rd_cycle[11332] = 1'b1;  wr_cycle[11332] = 1'b0;  addr_rom[11332]='h00002710;  wr_data_rom[11332]='h00000000;
    rd_cycle[11333] = 1'b1;  wr_cycle[11333] = 1'b0;  addr_rom[11333]='h00003fd8;  wr_data_rom[11333]='h00000000;
    rd_cycle[11334] = 1'b0;  wr_cycle[11334] = 1'b1;  addr_rom[11334]='h000034f0;  wr_data_rom[11334]='h00003320;
    rd_cycle[11335] = 1'b1;  wr_cycle[11335] = 1'b0;  addr_rom[11335]='h00003b78;  wr_data_rom[11335]='h00000000;
    rd_cycle[11336] = 1'b1;  wr_cycle[11336] = 1'b0;  addr_rom[11336]='h00002f80;  wr_data_rom[11336]='h00000000;
    rd_cycle[11337] = 1'b0;  wr_cycle[11337] = 1'b1;  addr_rom[11337]='h000035bc;  wr_data_rom[11337]='h00001789;
    rd_cycle[11338] = 1'b0;  wr_cycle[11338] = 1'b1;  addr_rom[11338]='h0000379c;  wr_data_rom[11338]='h00002702;
    rd_cycle[11339] = 1'b1;  wr_cycle[11339] = 1'b0;  addr_rom[11339]='h00001890;  wr_data_rom[11339]='h00000000;
    rd_cycle[11340] = 1'b1;  wr_cycle[11340] = 1'b0;  addr_rom[11340]='h000018ac;  wr_data_rom[11340]='h00000000;
    rd_cycle[11341] = 1'b1;  wr_cycle[11341] = 1'b0;  addr_rom[11341]='h00000418;  wr_data_rom[11341]='h00000000;
    rd_cycle[11342] = 1'b0;  wr_cycle[11342] = 1'b1;  addr_rom[11342]='h00000138;  wr_data_rom[11342]='h00003652;
    rd_cycle[11343] = 1'b1;  wr_cycle[11343] = 1'b0;  addr_rom[11343]='h00000bd0;  wr_data_rom[11343]='h00000000;
    rd_cycle[11344] = 1'b0;  wr_cycle[11344] = 1'b1;  addr_rom[11344]='h00000db0;  wr_data_rom[11344]='h00003b37;
    rd_cycle[11345] = 1'b1;  wr_cycle[11345] = 1'b0;  addr_rom[11345]='h000015e0;  wr_data_rom[11345]='h00000000;
    rd_cycle[11346] = 1'b0;  wr_cycle[11346] = 1'b1;  addr_rom[11346]='h00001fec;  wr_data_rom[11346]='h0000307e;
    rd_cycle[11347] = 1'b1;  wr_cycle[11347] = 1'b0;  addr_rom[11347]='h00001000;  wr_data_rom[11347]='h00000000;
    rd_cycle[11348] = 1'b0;  wr_cycle[11348] = 1'b1;  addr_rom[11348]='h00003e18;  wr_data_rom[11348]='h00000e77;
    rd_cycle[11349] = 1'b0;  wr_cycle[11349] = 1'b1;  addr_rom[11349]='h00001f94;  wr_data_rom[11349]='h00002b77;
    rd_cycle[11350] = 1'b1;  wr_cycle[11350] = 1'b0;  addr_rom[11350]='h000029cc;  wr_data_rom[11350]='h00000000;
    rd_cycle[11351] = 1'b1;  wr_cycle[11351] = 1'b0;  addr_rom[11351]='h00001a08;  wr_data_rom[11351]='h00000000;
    rd_cycle[11352] = 1'b1;  wr_cycle[11352] = 1'b0;  addr_rom[11352]='h00003400;  wr_data_rom[11352]='h00000000;
    rd_cycle[11353] = 1'b1;  wr_cycle[11353] = 1'b0;  addr_rom[11353]='h000018fc;  wr_data_rom[11353]='h00000000;
    rd_cycle[11354] = 1'b0;  wr_cycle[11354] = 1'b1;  addr_rom[11354]='h0000178c;  wr_data_rom[11354]='h00002637;
    rd_cycle[11355] = 1'b1;  wr_cycle[11355] = 1'b0;  addr_rom[11355]='h00003144;  wr_data_rom[11355]='h00000000;
    rd_cycle[11356] = 1'b0;  wr_cycle[11356] = 1'b1;  addr_rom[11356]='h000025d8;  wr_data_rom[11356]='h00003b50;
    rd_cycle[11357] = 1'b1;  wr_cycle[11357] = 1'b0;  addr_rom[11357]='h00003b54;  wr_data_rom[11357]='h00000000;
    rd_cycle[11358] = 1'b1;  wr_cycle[11358] = 1'b0;  addr_rom[11358]='h00000a34;  wr_data_rom[11358]='h00000000;
    rd_cycle[11359] = 1'b1;  wr_cycle[11359] = 1'b0;  addr_rom[11359]='h000004c4;  wr_data_rom[11359]='h00000000;
    rd_cycle[11360] = 1'b0;  wr_cycle[11360] = 1'b1;  addr_rom[11360]='h00000cc8;  wr_data_rom[11360]='h00002370;
    rd_cycle[11361] = 1'b1;  wr_cycle[11361] = 1'b0;  addr_rom[11361]='h00001ed4;  wr_data_rom[11361]='h00000000;
    rd_cycle[11362] = 1'b1;  wr_cycle[11362] = 1'b0;  addr_rom[11362]='h00002794;  wr_data_rom[11362]='h00000000;
    rd_cycle[11363] = 1'b0;  wr_cycle[11363] = 1'b1;  addr_rom[11363]='h000001d8;  wr_data_rom[11363]='h00003583;
    rd_cycle[11364] = 1'b1;  wr_cycle[11364] = 1'b0;  addr_rom[11364]='h00002958;  wr_data_rom[11364]='h00000000;
    rd_cycle[11365] = 1'b1;  wr_cycle[11365] = 1'b0;  addr_rom[11365]='h0000343c;  wr_data_rom[11365]='h00000000;
    rd_cycle[11366] = 1'b0;  wr_cycle[11366] = 1'b1;  addr_rom[11366]='h00000818;  wr_data_rom[11366]='h00003608;
    rd_cycle[11367] = 1'b1;  wr_cycle[11367] = 1'b0;  addr_rom[11367]='h00000b68;  wr_data_rom[11367]='h00000000;
    rd_cycle[11368] = 1'b0;  wr_cycle[11368] = 1'b1;  addr_rom[11368]='h00003b14;  wr_data_rom[11368]='h0000127c;
    rd_cycle[11369] = 1'b0;  wr_cycle[11369] = 1'b1;  addr_rom[11369]='h00003974;  wr_data_rom[11369]='h00003fdd;
    rd_cycle[11370] = 1'b0;  wr_cycle[11370] = 1'b1;  addr_rom[11370]='h00003118;  wr_data_rom[11370]='h000015a7;
    rd_cycle[11371] = 1'b1;  wr_cycle[11371] = 1'b0;  addr_rom[11371]='h00002be0;  wr_data_rom[11371]='h00000000;
    rd_cycle[11372] = 1'b1;  wr_cycle[11372] = 1'b0;  addr_rom[11372]='h00002e1c;  wr_data_rom[11372]='h00000000;
    rd_cycle[11373] = 1'b1;  wr_cycle[11373] = 1'b0;  addr_rom[11373]='h00002584;  wr_data_rom[11373]='h00000000;
    rd_cycle[11374] = 1'b1;  wr_cycle[11374] = 1'b0;  addr_rom[11374]='h00002798;  wr_data_rom[11374]='h00000000;
    rd_cycle[11375] = 1'b0;  wr_cycle[11375] = 1'b1;  addr_rom[11375]='h00003908;  wr_data_rom[11375]='h00000106;
    rd_cycle[11376] = 1'b1;  wr_cycle[11376] = 1'b0;  addr_rom[11376]='h00003198;  wr_data_rom[11376]='h00000000;
    rd_cycle[11377] = 1'b1;  wr_cycle[11377] = 1'b0;  addr_rom[11377]='h000021fc;  wr_data_rom[11377]='h00000000;
    rd_cycle[11378] = 1'b0;  wr_cycle[11378] = 1'b1;  addr_rom[11378]='h00003868;  wr_data_rom[11378]='h00002040;
    rd_cycle[11379] = 1'b0;  wr_cycle[11379] = 1'b1;  addr_rom[11379]='h000037dc;  wr_data_rom[11379]='h00001878;
    rd_cycle[11380] = 1'b1;  wr_cycle[11380] = 1'b0;  addr_rom[11380]='h000029dc;  wr_data_rom[11380]='h00000000;
    rd_cycle[11381] = 1'b1;  wr_cycle[11381] = 1'b0;  addr_rom[11381]='h00001728;  wr_data_rom[11381]='h00000000;
    rd_cycle[11382] = 1'b1;  wr_cycle[11382] = 1'b0;  addr_rom[11382]='h00002880;  wr_data_rom[11382]='h00000000;
    rd_cycle[11383] = 1'b0;  wr_cycle[11383] = 1'b1;  addr_rom[11383]='h000034a0;  wr_data_rom[11383]='h0000111e;
    rd_cycle[11384] = 1'b1;  wr_cycle[11384] = 1'b0;  addr_rom[11384]='h00002bb8;  wr_data_rom[11384]='h00000000;
    rd_cycle[11385] = 1'b0;  wr_cycle[11385] = 1'b1;  addr_rom[11385]='h000010f0;  wr_data_rom[11385]='h00002518;
    rd_cycle[11386] = 1'b1;  wr_cycle[11386] = 1'b0;  addr_rom[11386]='h00002760;  wr_data_rom[11386]='h00000000;
    rd_cycle[11387] = 1'b1;  wr_cycle[11387] = 1'b0;  addr_rom[11387]='h0000098c;  wr_data_rom[11387]='h00000000;
    rd_cycle[11388] = 1'b0;  wr_cycle[11388] = 1'b1;  addr_rom[11388]='h000014bc;  wr_data_rom[11388]='h00003637;
    rd_cycle[11389] = 1'b1;  wr_cycle[11389] = 1'b0;  addr_rom[11389]='h00003ae8;  wr_data_rom[11389]='h00000000;
    rd_cycle[11390] = 1'b0;  wr_cycle[11390] = 1'b1;  addr_rom[11390]='h00001bb4;  wr_data_rom[11390]='h000002a1;
    rd_cycle[11391] = 1'b0;  wr_cycle[11391] = 1'b1;  addr_rom[11391]='h000009e4;  wr_data_rom[11391]='h0000252a;
    rd_cycle[11392] = 1'b0;  wr_cycle[11392] = 1'b1;  addr_rom[11392]='h00001b84;  wr_data_rom[11392]='h00000817;
    rd_cycle[11393] = 1'b0;  wr_cycle[11393] = 1'b1;  addr_rom[11393]='h00001258;  wr_data_rom[11393]='h000013bc;
    rd_cycle[11394] = 1'b1;  wr_cycle[11394] = 1'b0;  addr_rom[11394]='h00001d38;  wr_data_rom[11394]='h00000000;
    rd_cycle[11395] = 1'b0;  wr_cycle[11395] = 1'b1;  addr_rom[11395]='h00000bd8;  wr_data_rom[11395]='h000038de;
    rd_cycle[11396] = 1'b0;  wr_cycle[11396] = 1'b1;  addr_rom[11396]='h00003b38;  wr_data_rom[11396]='h00000cd0;
    rd_cycle[11397] = 1'b0;  wr_cycle[11397] = 1'b1;  addr_rom[11397]='h000017bc;  wr_data_rom[11397]='h00001864;
    rd_cycle[11398] = 1'b1;  wr_cycle[11398] = 1'b0;  addr_rom[11398]='h00003160;  wr_data_rom[11398]='h00000000;
    rd_cycle[11399] = 1'b1;  wr_cycle[11399] = 1'b0;  addr_rom[11399]='h00001768;  wr_data_rom[11399]='h00000000;
    rd_cycle[11400] = 1'b1;  wr_cycle[11400] = 1'b0;  addr_rom[11400]='h000032e8;  wr_data_rom[11400]='h00000000;
    rd_cycle[11401] = 1'b0;  wr_cycle[11401] = 1'b1;  addr_rom[11401]='h0000076c;  wr_data_rom[11401]='h000022ca;
    rd_cycle[11402] = 1'b1;  wr_cycle[11402] = 1'b0;  addr_rom[11402]='h00000288;  wr_data_rom[11402]='h00000000;
    rd_cycle[11403] = 1'b0;  wr_cycle[11403] = 1'b1;  addr_rom[11403]='h000033d0;  wr_data_rom[11403]='h00002acc;
    rd_cycle[11404] = 1'b1;  wr_cycle[11404] = 1'b0;  addr_rom[11404]='h0000382c;  wr_data_rom[11404]='h00000000;
    rd_cycle[11405] = 1'b1;  wr_cycle[11405] = 1'b0;  addr_rom[11405]='h00002ffc;  wr_data_rom[11405]='h00000000;
    rd_cycle[11406] = 1'b1;  wr_cycle[11406] = 1'b0;  addr_rom[11406]='h000008ec;  wr_data_rom[11406]='h00000000;
    rd_cycle[11407] = 1'b1;  wr_cycle[11407] = 1'b0;  addr_rom[11407]='h00001a7c;  wr_data_rom[11407]='h00000000;
    rd_cycle[11408] = 1'b0;  wr_cycle[11408] = 1'b1;  addr_rom[11408]='h00000ad0;  wr_data_rom[11408]='h000035d4;
    rd_cycle[11409] = 1'b1;  wr_cycle[11409] = 1'b0;  addr_rom[11409]='h0000116c;  wr_data_rom[11409]='h00000000;
    rd_cycle[11410] = 1'b1;  wr_cycle[11410] = 1'b0;  addr_rom[11410]='h00001304;  wr_data_rom[11410]='h00000000;
    rd_cycle[11411] = 1'b0;  wr_cycle[11411] = 1'b1;  addr_rom[11411]='h00003368;  wr_data_rom[11411]='h000016f5;
    rd_cycle[11412] = 1'b1;  wr_cycle[11412] = 1'b0;  addr_rom[11412]='h000012e8;  wr_data_rom[11412]='h00000000;
    rd_cycle[11413] = 1'b0;  wr_cycle[11413] = 1'b1;  addr_rom[11413]='h00000e68;  wr_data_rom[11413]='h00003a7b;
    rd_cycle[11414] = 1'b1;  wr_cycle[11414] = 1'b0;  addr_rom[11414]='h000026d0;  wr_data_rom[11414]='h00000000;
    rd_cycle[11415] = 1'b1;  wr_cycle[11415] = 1'b0;  addr_rom[11415]='h00001ee8;  wr_data_rom[11415]='h00000000;
    rd_cycle[11416] = 1'b1;  wr_cycle[11416] = 1'b0;  addr_rom[11416]='h00000828;  wr_data_rom[11416]='h00000000;
    rd_cycle[11417] = 1'b0;  wr_cycle[11417] = 1'b1;  addr_rom[11417]='h00000984;  wr_data_rom[11417]='h00002db5;
    rd_cycle[11418] = 1'b1;  wr_cycle[11418] = 1'b0;  addr_rom[11418]='h0000311c;  wr_data_rom[11418]='h00000000;
    rd_cycle[11419] = 1'b0;  wr_cycle[11419] = 1'b1;  addr_rom[11419]='h00002010;  wr_data_rom[11419]='h000030e3;
    rd_cycle[11420] = 1'b1;  wr_cycle[11420] = 1'b0;  addr_rom[11420]='h00001008;  wr_data_rom[11420]='h00000000;
    rd_cycle[11421] = 1'b0;  wr_cycle[11421] = 1'b1;  addr_rom[11421]='h00002b78;  wr_data_rom[11421]='h00000bec;
    rd_cycle[11422] = 1'b1;  wr_cycle[11422] = 1'b0;  addr_rom[11422]='h00001478;  wr_data_rom[11422]='h00000000;
    rd_cycle[11423] = 1'b0;  wr_cycle[11423] = 1'b1;  addr_rom[11423]='h000028bc;  wr_data_rom[11423]='h000009fd;
    rd_cycle[11424] = 1'b0;  wr_cycle[11424] = 1'b1;  addr_rom[11424]='h00000d80;  wr_data_rom[11424]='h000003c8;
    rd_cycle[11425] = 1'b1;  wr_cycle[11425] = 1'b0;  addr_rom[11425]='h000014e8;  wr_data_rom[11425]='h00000000;
    rd_cycle[11426] = 1'b1;  wr_cycle[11426] = 1'b0;  addr_rom[11426]='h00002c78;  wr_data_rom[11426]='h00000000;
    rd_cycle[11427] = 1'b1;  wr_cycle[11427] = 1'b0;  addr_rom[11427]='h00002a10;  wr_data_rom[11427]='h00000000;
    rd_cycle[11428] = 1'b0;  wr_cycle[11428] = 1'b1;  addr_rom[11428]='h00000348;  wr_data_rom[11428]='h0000342d;
    rd_cycle[11429] = 1'b1;  wr_cycle[11429] = 1'b0;  addr_rom[11429]='h00002874;  wr_data_rom[11429]='h00000000;
    rd_cycle[11430] = 1'b0;  wr_cycle[11430] = 1'b1;  addr_rom[11430]='h00000294;  wr_data_rom[11430]='h000007a7;
    rd_cycle[11431] = 1'b1;  wr_cycle[11431] = 1'b0;  addr_rom[11431]='h00000cfc;  wr_data_rom[11431]='h00000000;
    rd_cycle[11432] = 1'b1;  wr_cycle[11432] = 1'b0;  addr_rom[11432]='h000021a0;  wr_data_rom[11432]='h00000000;
    rd_cycle[11433] = 1'b0;  wr_cycle[11433] = 1'b1;  addr_rom[11433]='h0000340c;  wr_data_rom[11433]='h000038d5;
    rd_cycle[11434] = 1'b1;  wr_cycle[11434] = 1'b0;  addr_rom[11434]='h000037dc;  wr_data_rom[11434]='h00000000;
    rd_cycle[11435] = 1'b1;  wr_cycle[11435] = 1'b0;  addr_rom[11435]='h0000377c;  wr_data_rom[11435]='h00000000;
    rd_cycle[11436] = 1'b1;  wr_cycle[11436] = 1'b0;  addr_rom[11436]='h00000918;  wr_data_rom[11436]='h00000000;
    rd_cycle[11437] = 1'b1;  wr_cycle[11437] = 1'b0;  addr_rom[11437]='h00003fac;  wr_data_rom[11437]='h00000000;
    rd_cycle[11438] = 1'b1;  wr_cycle[11438] = 1'b0;  addr_rom[11438]='h00000f28;  wr_data_rom[11438]='h00000000;
    rd_cycle[11439] = 1'b1;  wr_cycle[11439] = 1'b0;  addr_rom[11439]='h00003044;  wr_data_rom[11439]='h00000000;
    rd_cycle[11440] = 1'b0;  wr_cycle[11440] = 1'b1;  addr_rom[11440]='h00001944;  wr_data_rom[11440]='h00000aaa;
    rd_cycle[11441] = 1'b1;  wr_cycle[11441] = 1'b0;  addr_rom[11441]='h00001608;  wr_data_rom[11441]='h00000000;
    rd_cycle[11442] = 1'b0;  wr_cycle[11442] = 1'b1;  addr_rom[11442]='h000011a4;  wr_data_rom[11442]='h00002ac6;
    rd_cycle[11443] = 1'b0;  wr_cycle[11443] = 1'b1;  addr_rom[11443]='h0000335c;  wr_data_rom[11443]='h00002e70;
    rd_cycle[11444] = 1'b0;  wr_cycle[11444] = 1'b1;  addr_rom[11444]='h00001d40;  wr_data_rom[11444]='h00003388;
    rd_cycle[11445] = 1'b0;  wr_cycle[11445] = 1'b1;  addr_rom[11445]='h00001344;  wr_data_rom[11445]='h00000d16;
    rd_cycle[11446] = 1'b1;  wr_cycle[11446] = 1'b0;  addr_rom[11446]='h000000d4;  wr_data_rom[11446]='h00000000;
    rd_cycle[11447] = 1'b1;  wr_cycle[11447] = 1'b0;  addr_rom[11447]='h00003ca0;  wr_data_rom[11447]='h00000000;
    rd_cycle[11448] = 1'b1;  wr_cycle[11448] = 1'b0;  addr_rom[11448]='h00000fac;  wr_data_rom[11448]='h00000000;
    rd_cycle[11449] = 1'b1;  wr_cycle[11449] = 1'b0;  addr_rom[11449]='h0000395c;  wr_data_rom[11449]='h00000000;
    rd_cycle[11450] = 1'b0;  wr_cycle[11450] = 1'b1;  addr_rom[11450]='h00003d1c;  wr_data_rom[11450]='h000028cd;
    rd_cycle[11451] = 1'b0;  wr_cycle[11451] = 1'b1;  addr_rom[11451]='h000032d8;  wr_data_rom[11451]='h000003a5;
    rd_cycle[11452] = 1'b0;  wr_cycle[11452] = 1'b1;  addr_rom[11452]='h00003fcc;  wr_data_rom[11452]='h00001cc8;
    rd_cycle[11453] = 1'b0;  wr_cycle[11453] = 1'b1;  addr_rom[11453]='h000029f0;  wr_data_rom[11453]='h00001077;
    rd_cycle[11454] = 1'b1;  wr_cycle[11454] = 1'b0;  addr_rom[11454]='h000004b4;  wr_data_rom[11454]='h00000000;
    rd_cycle[11455] = 1'b1;  wr_cycle[11455] = 1'b0;  addr_rom[11455]='h00002330;  wr_data_rom[11455]='h00000000;
    rd_cycle[11456] = 1'b1;  wr_cycle[11456] = 1'b0;  addr_rom[11456]='h000014a8;  wr_data_rom[11456]='h00000000;
    rd_cycle[11457] = 1'b0;  wr_cycle[11457] = 1'b1;  addr_rom[11457]='h0000165c;  wr_data_rom[11457]='h00001822;
    rd_cycle[11458] = 1'b1;  wr_cycle[11458] = 1'b0;  addr_rom[11458]='h00001914;  wr_data_rom[11458]='h00000000;
    rd_cycle[11459] = 1'b0;  wr_cycle[11459] = 1'b1;  addr_rom[11459]='h0000122c;  wr_data_rom[11459]='h00002d06;
    rd_cycle[11460] = 1'b0;  wr_cycle[11460] = 1'b1;  addr_rom[11460]='h00001bf8;  wr_data_rom[11460]='h00002ada;
    rd_cycle[11461] = 1'b0;  wr_cycle[11461] = 1'b1;  addr_rom[11461]='h00000900;  wr_data_rom[11461]='h000019ed;
    rd_cycle[11462] = 1'b1;  wr_cycle[11462] = 1'b0;  addr_rom[11462]='h00002c14;  wr_data_rom[11462]='h00000000;
    rd_cycle[11463] = 1'b1;  wr_cycle[11463] = 1'b0;  addr_rom[11463]='h000007e8;  wr_data_rom[11463]='h00000000;
    rd_cycle[11464] = 1'b1;  wr_cycle[11464] = 1'b0;  addr_rom[11464]='h0000143c;  wr_data_rom[11464]='h00000000;
    rd_cycle[11465] = 1'b0;  wr_cycle[11465] = 1'b1;  addr_rom[11465]='h00003a0c;  wr_data_rom[11465]='h000012ff;
    rd_cycle[11466] = 1'b1;  wr_cycle[11466] = 1'b0;  addr_rom[11466]='h00002d00;  wr_data_rom[11466]='h00000000;
    rd_cycle[11467] = 1'b1;  wr_cycle[11467] = 1'b0;  addr_rom[11467]='h000024e4;  wr_data_rom[11467]='h00000000;
    rd_cycle[11468] = 1'b0;  wr_cycle[11468] = 1'b1;  addr_rom[11468]='h000038a4;  wr_data_rom[11468]='h00003397;
    rd_cycle[11469] = 1'b0;  wr_cycle[11469] = 1'b1;  addr_rom[11469]='h00002d3c;  wr_data_rom[11469]='h00000f22;
    rd_cycle[11470] = 1'b0;  wr_cycle[11470] = 1'b1;  addr_rom[11470]='h00001b7c;  wr_data_rom[11470]='h0000066a;
    rd_cycle[11471] = 1'b0;  wr_cycle[11471] = 1'b1;  addr_rom[11471]='h00003d50;  wr_data_rom[11471]='h00001f74;
    rd_cycle[11472] = 1'b0;  wr_cycle[11472] = 1'b1;  addr_rom[11472]='h00000c08;  wr_data_rom[11472]='h0000173d;
    rd_cycle[11473] = 1'b1;  wr_cycle[11473] = 1'b0;  addr_rom[11473]='h000018fc;  wr_data_rom[11473]='h00000000;
    rd_cycle[11474] = 1'b0;  wr_cycle[11474] = 1'b1;  addr_rom[11474]='h00001ca4;  wr_data_rom[11474]='h00003d11;
    rd_cycle[11475] = 1'b1;  wr_cycle[11475] = 1'b0;  addr_rom[11475]='h00003784;  wr_data_rom[11475]='h00000000;
    rd_cycle[11476] = 1'b0;  wr_cycle[11476] = 1'b1;  addr_rom[11476]='h000014c0;  wr_data_rom[11476]='h00000c9f;
    rd_cycle[11477] = 1'b1;  wr_cycle[11477] = 1'b0;  addr_rom[11477]='h00001170;  wr_data_rom[11477]='h00000000;
    rd_cycle[11478] = 1'b0;  wr_cycle[11478] = 1'b1;  addr_rom[11478]='h00000670;  wr_data_rom[11478]='h000002eb;
    rd_cycle[11479] = 1'b0;  wr_cycle[11479] = 1'b1;  addr_rom[11479]='h000026fc;  wr_data_rom[11479]='h000036aa;
    rd_cycle[11480] = 1'b0;  wr_cycle[11480] = 1'b1;  addr_rom[11480]='h000023cc;  wr_data_rom[11480]='h000030da;
    rd_cycle[11481] = 1'b1;  wr_cycle[11481] = 1'b0;  addr_rom[11481]='h00000838;  wr_data_rom[11481]='h00000000;
    rd_cycle[11482] = 1'b0;  wr_cycle[11482] = 1'b1;  addr_rom[11482]='h0000342c;  wr_data_rom[11482]='h00001010;
    rd_cycle[11483] = 1'b0;  wr_cycle[11483] = 1'b1;  addr_rom[11483]='h00001024;  wr_data_rom[11483]='h00003c9c;
    rd_cycle[11484] = 1'b1;  wr_cycle[11484] = 1'b0;  addr_rom[11484]='h00002410;  wr_data_rom[11484]='h00000000;
    rd_cycle[11485] = 1'b0;  wr_cycle[11485] = 1'b1;  addr_rom[11485]='h00001fd0;  wr_data_rom[11485]='h000000f9;
    rd_cycle[11486] = 1'b0;  wr_cycle[11486] = 1'b1;  addr_rom[11486]='h0000085c;  wr_data_rom[11486]='h000035e0;
    rd_cycle[11487] = 1'b0;  wr_cycle[11487] = 1'b1;  addr_rom[11487]='h000001f4;  wr_data_rom[11487]='h0000155b;
    rd_cycle[11488] = 1'b1;  wr_cycle[11488] = 1'b0;  addr_rom[11488]='h0000000c;  wr_data_rom[11488]='h00000000;
    rd_cycle[11489] = 1'b1;  wr_cycle[11489] = 1'b0;  addr_rom[11489]='h00000bcc;  wr_data_rom[11489]='h00000000;
    rd_cycle[11490] = 1'b0;  wr_cycle[11490] = 1'b1;  addr_rom[11490]='h000000bc;  wr_data_rom[11490]='h000033ee;
    rd_cycle[11491] = 1'b1;  wr_cycle[11491] = 1'b0;  addr_rom[11491]='h000023f8;  wr_data_rom[11491]='h00000000;
    rd_cycle[11492] = 1'b1;  wr_cycle[11492] = 1'b0;  addr_rom[11492]='h00002838;  wr_data_rom[11492]='h00000000;
    rd_cycle[11493] = 1'b0;  wr_cycle[11493] = 1'b1;  addr_rom[11493]='h00002dfc;  wr_data_rom[11493]='h000029ae;
    rd_cycle[11494] = 1'b0;  wr_cycle[11494] = 1'b1;  addr_rom[11494]='h00000164;  wr_data_rom[11494]='h0000233d;
    rd_cycle[11495] = 1'b0;  wr_cycle[11495] = 1'b1;  addr_rom[11495]='h00002980;  wr_data_rom[11495]='h0000325c;
    rd_cycle[11496] = 1'b0;  wr_cycle[11496] = 1'b1;  addr_rom[11496]='h00002f40;  wr_data_rom[11496]='h000017b9;
    rd_cycle[11497] = 1'b0;  wr_cycle[11497] = 1'b1;  addr_rom[11497]='h00002dcc;  wr_data_rom[11497]='h00003451;
    rd_cycle[11498] = 1'b0;  wr_cycle[11498] = 1'b1;  addr_rom[11498]='h00001758;  wr_data_rom[11498]='h000010ff;
    rd_cycle[11499] = 1'b1;  wr_cycle[11499] = 1'b0;  addr_rom[11499]='h00003e14;  wr_data_rom[11499]='h00000000;
    rd_cycle[11500] = 1'b0;  wr_cycle[11500] = 1'b1;  addr_rom[11500]='h000027f0;  wr_data_rom[11500]='h00003cb2;
    rd_cycle[11501] = 1'b0;  wr_cycle[11501] = 1'b1;  addr_rom[11501]='h000010a8;  wr_data_rom[11501]='h000032ee;
    rd_cycle[11502] = 1'b0;  wr_cycle[11502] = 1'b1;  addr_rom[11502]='h000007c0;  wr_data_rom[11502]='h00001834;
    rd_cycle[11503] = 1'b1;  wr_cycle[11503] = 1'b0;  addr_rom[11503]='h000030c8;  wr_data_rom[11503]='h00000000;
    rd_cycle[11504] = 1'b0;  wr_cycle[11504] = 1'b1;  addr_rom[11504]='h0000192c;  wr_data_rom[11504]='h00003f46;
    rd_cycle[11505] = 1'b0;  wr_cycle[11505] = 1'b1;  addr_rom[11505]='h00000ae4;  wr_data_rom[11505]='h0000187d;
    rd_cycle[11506] = 1'b0;  wr_cycle[11506] = 1'b1;  addr_rom[11506]='h00002d4c;  wr_data_rom[11506]='h00003b89;
    rd_cycle[11507] = 1'b0;  wr_cycle[11507] = 1'b1;  addr_rom[11507]='h000030ac;  wr_data_rom[11507]='h00001f57;
    rd_cycle[11508] = 1'b1;  wr_cycle[11508] = 1'b0;  addr_rom[11508]='h000025b8;  wr_data_rom[11508]='h00000000;
    rd_cycle[11509] = 1'b1;  wr_cycle[11509] = 1'b0;  addr_rom[11509]='h00003610;  wr_data_rom[11509]='h00000000;
    rd_cycle[11510] = 1'b0;  wr_cycle[11510] = 1'b1;  addr_rom[11510]='h00001c50;  wr_data_rom[11510]='h00001dcc;
    rd_cycle[11511] = 1'b1;  wr_cycle[11511] = 1'b0;  addr_rom[11511]='h000037b8;  wr_data_rom[11511]='h00000000;
    rd_cycle[11512] = 1'b1;  wr_cycle[11512] = 1'b0;  addr_rom[11512]='h00001238;  wr_data_rom[11512]='h00000000;
    rd_cycle[11513] = 1'b0;  wr_cycle[11513] = 1'b1;  addr_rom[11513]='h00001598;  wr_data_rom[11513]='h00003e31;
    rd_cycle[11514] = 1'b0;  wr_cycle[11514] = 1'b1;  addr_rom[11514]='h00000da8;  wr_data_rom[11514]='h00003f08;
    rd_cycle[11515] = 1'b0;  wr_cycle[11515] = 1'b1;  addr_rom[11515]='h00002460;  wr_data_rom[11515]='h000005bf;
    rd_cycle[11516] = 1'b0;  wr_cycle[11516] = 1'b1;  addr_rom[11516]='h00002030;  wr_data_rom[11516]='h00000dbb;
    rd_cycle[11517] = 1'b1;  wr_cycle[11517] = 1'b0;  addr_rom[11517]='h00001e40;  wr_data_rom[11517]='h00000000;
    rd_cycle[11518] = 1'b1;  wr_cycle[11518] = 1'b0;  addr_rom[11518]='h000003d4;  wr_data_rom[11518]='h00000000;
    rd_cycle[11519] = 1'b0;  wr_cycle[11519] = 1'b1;  addr_rom[11519]='h00002564;  wr_data_rom[11519]='h00003a2e;
    rd_cycle[11520] = 1'b1;  wr_cycle[11520] = 1'b0;  addr_rom[11520]='h00002790;  wr_data_rom[11520]='h00000000;
    rd_cycle[11521] = 1'b1;  wr_cycle[11521] = 1'b0;  addr_rom[11521]='h00002c84;  wr_data_rom[11521]='h00000000;
    rd_cycle[11522] = 1'b0;  wr_cycle[11522] = 1'b1;  addr_rom[11522]='h00001d48;  wr_data_rom[11522]='h00002ba9;
    rd_cycle[11523] = 1'b1;  wr_cycle[11523] = 1'b0;  addr_rom[11523]='h00003340;  wr_data_rom[11523]='h00000000;
    rd_cycle[11524] = 1'b1;  wr_cycle[11524] = 1'b0;  addr_rom[11524]='h000005a4;  wr_data_rom[11524]='h00000000;
    rd_cycle[11525] = 1'b1;  wr_cycle[11525] = 1'b0;  addr_rom[11525]='h000018d0;  wr_data_rom[11525]='h00000000;
    rd_cycle[11526] = 1'b0;  wr_cycle[11526] = 1'b1;  addr_rom[11526]='h00002258;  wr_data_rom[11526]='h0000381c;
    rd_cycle[11527] = 1'b0;  wr_cycle[11527] = 1'b1;  addr_rom[11527]='h0000215c;  wr_data_rom[11527]='h00001d75;
    rd_cycle[11528] = 1'b1;  wr_cycle[11528] = 1'b0;  addr_rom[11528]='h00003598;  wr_data_rom[11528]='h00000000;
    rd_cycle[11529] = 1'b0;  wr_cycle[11529] = 1'b1;  addr_rom[11529]='h00001074;  wr_data_rom[11529]='h00001989;
    rd_cycle[11530] = 1'b0;  wr_cycle[11530] = 1'b1;  addr_rom[11530]='h000037c8;  wr_data_rom[11530]='h00000637;
    rd_cycle[11531] = 1'b0;  wr_cycle[11531] = 1'b1;  addr_rom[11531]='h00001f70;  wr_data_rom[11531]='h00002923;
    rd_cycle[11532] = 1'b1;  wr_cycle[11532] = 1'b0;  addr_rom[11532]='h00002414;  wr_data_rom[11532]='h00000000;
    rd_cycle[11533] = 1'b1;  wr_cycle[11533] = 1'b0;  addr_rom[11533]='h00001850;  wr_data_rom[11533]='h00000000;
    rd_cycle[11534] = 1'b0;  wr_cycle[11534] = 1'b1;  addr_rom[11534]='h00000b1c;  wr_data_rom[11534]='h00002885;
    rd_cycle[11535] = 1'b1;  wr_cycle[11535] = 1'b0;  addr_rom[11535]='h00003c6c;  wr_data_rom[11535]='h00000000;
    rd_cycle[11536] = 1'b0;  wr_cycle[11536] = 1'b1;  addr_rom[11536]='h00001d80;  wr_data_rom[11536]='h000038db;
    rd_cycle[11537] = 1'b1;  wr_cycle[11537] = 1'b0;  addr_rom[11537]='h00003800;  wr_data_rom[11537]='h00000000;
    rd_cycle[11538] = 1'b0;  wr_cycle[11538] = 1'b1;  addr_rom[11538]='h00003f40;  wr_data_rom[11538]='h000022a2;
    rd_cycle[11539] = 1'b1;  wr_cycle[11539] = 1'b0;  addr_rom[11539]='h000005e8;  wr_data_rom[11539]='h00000000;
    rd_cycle[11540] = 1'b0;  wr_cycle[11540] = 1'b1;  addr_rom[11540]='h000038e4;  wr_data_rom[11540]='h000007d6;
    rd_cycle[11541] = 1'b1;  wr_cycle[11541] = 1'b0;  addr_rom[11541]='h0000242c;  wr_data_rom[11541]='h00000000;
    rd_cycle[11542] = 1'b1;  wr_cycle[11542] = 1'b0;  addr_rom[11542]='h000025f8;  wr_data_rom[11542]='h00000000;
    rd_cycle[11543] = 1'b0;  wr_cycle[11543] = 1'b1;  addr_rom[11543]='h00001adc;  wr_data_rom[11543]='h00000edd;
    rd_cycle[11544] = 1'b1;  wr_cycle[11544] = 1'b0;  addr_rom[11544]='h00001960;  wr_data_rom[11544]='h00000000;
    rd_cycle[11545] = 1'b0;  wr_cycle[11545] = 1'b1;  addr_rom[11545]='h00000970;  wr_data_rom[11545]='h00003617;
    rd_cycle[11546] = 1'b1;  wr_cycle[11546] = 1'b0;  addr_rom[11546]='h00003a7c;  wr_data_rom[11546]='h00000000;
    rd_cycle[11547] = 1'b1;  wr_cycle[11547] = 1'b0;  addr_rom[11547]='h00001a90;  wr_data_rom[11547]='h00000000;
    rd_cycle[11548] = 1'b1;  wr_cycle[11548] = 1'b0;  addr_rom[11548]='h0000215c;  wr_data_rom[11548]='h00000000;
    rd_cycle[11549] = 1'b0;  wr_cycle[11549] = 1'b1;  addr_rom[11549]='h000038c0;  wr_data_rom[11549]='h00003c15;
    rd_cycle[11550] = 1'b0;  wr_cycle[11550] = 1'b1;  addr_rom[11550]='h00001c24;  wr_data_rom[11550]='h000039c3;
    rd_cycle[11551] = 1'b1;  wr_cycle[11551] = 1'b0;  addr_rom[11551]='h00003d1c;  wr_data_rom[11551]='h00000000;
    rd_cycle[11552] = 1'b0;  wr_cycle[11552] = 1'b1;  addr_rom[11552]='h0000026c;  wr_data_rom[11552]='h0000200e;
    rd_cycle[11553] = 1'b0;  wr_cycle[11553] = 1'b1;  addr_rom[11553]='h00003b08;  wr_data_rom[11553]='h000017a0;
    rd_cycle[11554] = 1'b0;  wr_cycle[11554] = 1'b1;  addr_rom[11554]='h00000cf0;  wr_data_rom[11554]='h000031a9;
    rd_cycle[11555] = 1'b1;  wr_cycle[11555] = 1'b0;  addr_rom[11555]='h000019b0;  wr_data_rom[11555]='h00000000;
    rd_cycle[11556] = 1'b1;  wr_cycle[11556] = 1'b0;  addr_rom[11556]='h000014d0;  wr_data_rom[11556]='h00000000;
    rd_cycle[11557] = 1'b1;  wr_cycle[11557] = 1'b0;  addr_rom[11557]='h00001568;  wr_data_rom[11557]='h00000000;
    rd_cycle[11558] = 1'b0;  wr_cycle[11558] = 1'b1;  addr_rom[11558]='h00001b74;  wr_data_rom[11558]='h000007dc;
    rd_cycle[11559] = 1'b0;  wr_cycle[11559] = 1'b1;  addr_rom[11559]='h000007d0;  wr_data_rom[11559]='h000030b4;
    rd_cycle[11560] = 1'b0;  wr_cycle[11560] = 1'b1;  addr_rom[11560]='h000016e4;  wr_data_rom[11560]='h000002ed;
    rd_cycle[11561] = 1'b1;  wr_cycle[11561] = 1'b0;  addr_rom[11561]='h0000252c;  wr_data_rom[11561]='h00000000;
    rd_cycle[11562] = 1'b0;  wr_cycle[11562] = 1'b1;  addr_rom[11562]='h00000bec;  wr_data_rom[11562]='h00003776;
    rd_cycle[11563] = 1'b0;  wr_cycle[11563] = 1'b1;  addr_rom[11563]='h00001a80;  wr_data_rom[11563]='h00002a0b;
    rd_cycle[11564] = 1'b1;  wr_cycle[11564] = 1'b0;  addr_rom[11564]='h00002bdc;  wr_data_rom[11564]='h00000000;
    rd_cycle[11565] = 1'b1;  wr_cycle[11565] = 1'b0;  addr_rom[11565]='h00003404;  wr_data_rom[11565]='h00000000;
    rd_cycle[11566] = 1'b0;  wr_cycle[11566] = 1'b1;  addr_rom[11566]='h000019d8;  wr_data_rom[11566]='h00000f99;
    rd_cycle[11567] = 1'b1;  wr_cycle[11567] = 1'b0;  addr_rom[11567]='h000004c0;  wr_data_rom[11567]='h00000000;
    rd_cycle[11568] = 1'b1;  wr_cycle[11568] = 1'b0;  addr_rom[11568]='h0000386c;  wr_data_rom[11568]='h00000000;
    rd_cycle[11569] = 1'b0;  wr_cycle[11569] = 1'b1;  addr_rom[11569]='h000025fc;  wr_data_rom[11569]='h000036c3;
    rd_cycle[11570] = 1'b0;  wr_cycle[11570] = 1'b1;  addr_rom[11570]='h00003ee4;  wr_data_rom[11570]='h00002344;
    rd_cycle[11571] = 1'b1;  wr_cycle[11571] = 1'b0;  addr_rom[11571]='h00001ea8;  wr_data_rom[11571]='h00000000;
    rd_cycle[11572] = 1'b1;  wr_cycle[11572] = 1'b0;  addr_rom[11572]='h00003084;  wr_data_rom[11572]='h00000000;
    rd_cycle[11573] = 1'b0;  wr_cycle[11573] = 1'b1;  addr_rom[11573]='h000015a4;  wr_data_rom[11573]='h000008e4;
    rd_cycle[11574] = 1'b0;  wr_cycle[11574] = 1'b1;  addr_rom[11574]='h00000898;  wr_data_rom[11574]='h00000db1;
    rd_cycle[11575] = 1'b0;  wr_cycle[11575] = 1'b1;  addr_rom[11575]='h00001e6c;  wr_data_rom[11575]='h00000d3f;
    rd_cycle[11576] = 1'b1;  wr_cycle[11576] = 1'b0;  addr_rom[11576]='h00000634;  wr_data_rom[11576]='h00000000;
    rd_cycle[11577] = 1'b0;  wr_cycle[11577] = 1'b1;  addr_rom[11577]='h00003a48;  wr_data_rom[11577]='h00001323;
    rd_cycle[11578] = 1'b1;  wr_cycle[11578] = 1'b0;  addr_rom[11578]='h000017a4;  wr_data_rom[11578]='h00000000;
    rd_cycle[11579] = 1'b1;  wr_cycle[11579] = 1'b0;  addr_rom[11579]='h00000950;  wr_data_rom[11579]='h00000000;
    rd_cycle[11580] = 1'b0;  wr_cycle[11580] = 1'b1;  addr_rom[11580]='h00001648;  wr_data_rom[11580]='h000032b6;
    rd_cycle[11581] = 1'b1;  wr_cycle[11581] = 1'b0;  addr_rom[11581]='h00003498;  wr_data_rom[11581]='h00000000;
    rd_cycle[11582] = 1'b0;  wr_cycle[11582] = 1'b1;  addr_rom[11582]='h00003ab8;  wr_data_rom[11582]='h00003054;
    rd_cycle[11583] = 1'b1;  wr_cycle[11583] = 1'b0;  addr_rom[11583]='h00002738;  wr_data_rom[11583]='h00000000;
    rd_cycle[11584] = 1'b1;  wr_cycle[11584] = 1'b0;  addr_rom[11584]='h00000868;  wr_data_rom[11584]='h00000000;
    rd_cycle[11585] = 1'b0;  wr_cycle[11585] = 1'b1;  addr_rom[11585]='h00002934;  wr_data_rom[11585]='h00003770;
    rd_cycle[11586] = 1'b1;  wr_cycle[11586] = 1'b0;  addr_rom[11586]='h00002484;  wr_data_rom[11586]='h00000000;
    rd_cycle[11587] = 1'b1;  wr_cycle[11587] = 1'b0;  addr_rom[11587]='h00000b4c;  wr_data_rom[11587]='h00000000;
    rd_cycle[11588] = 1'b1;  wr_cycle[11588] = 1'b0;  addr_rom[11588]='h00001e88;  wr_data_rom[11588]='h00000000;
    rd_cycle[11589] = 1'b1;  wr_cycle[11589] = 1'b0;  addr_rom[11589]='h00002b2c;  wr_data_rom[11589]='h00000000;
    rd_cycle[11590] = 1'b0;  wr_cycle[11590] = 1'b1;  addr_rom[11590]='h00000c0c;  wr_data_rom[11590]='h000010b6;
    rd_cycle[11591] = 1'b1;  wr_cycle[11591] = 1'b0;  addr_rom[11591]='h00001b84;  wr_data_rom[11591]='h00000000;
    rd_cycle[11592] = 1'b0;  wr_cycle[11592] = 1'b1;  addr_rom[11592]='h00000710;  wr_data_rom[11592]='h00002673;
    rd_cycle[11593] = 1'b0;  wr_cycle[11593] = 1'b1;  addr_rom[11593]='h0000181c;  wr_data_rom[11593]='h00001b30;
    rd_cycle[11594] = 1'b0;  wr_cycle[11594] = 1'b1;  addr_rom[11594]='h00002f4c;  wr_data_rom[11594]='h000006ac;
    rd_cycle[11595] = 1'b0;  wr_cycle[11595] = 1'b1;  addr_rom[11595]='h00003418;  wr_data_rom[11595]='h00003342;
    rd_cycle[11596] = 1'b0;  wr_cycle[11596] = 1'b1;  addr_rom[11596]='h00000390;  wr_data_rom[11596]='h00002c89;
    rd_cycle[11597] = 1'b0;  wr_cycle[11597] = 1'b1;  addr_rom[11597]='h00002614;  wr_data_rom[11597]='h0000248d;
    rd_cycle[11598] = 1'b0;  wr_cycle[11598] = 1'b1;  addr_rom[11598]='h000034c0;  wr_data_rom[11598]='h00002e55;
    rd_cycle[11599] = 1'b1;  wr_cycle[11599] = 1'b0;  addr_rom[11599]='h0000204c;  wr_data_rom[11599]='h00000000;
    rd_cycle[11600] = 1'b1;  wr_cycle[11600] = 1'b0;  addr_rom[11600]='h000034a0;  wr_data_rom[11600]='h00000000;
    rd_cycle[11601] = 1'b1;  wr_cycle[11601] = 1'b0;  addr_rom[11601]='h00002654;  wr_data_rom[11601]='h00000000;
    rd_cycle[11602] = 1'b1;  wr_cycle[11602] = 1'b0;  addr_rom[11602]='h00000a38;  wr_data_rom[11602]='h00000000;
    rd_cycle[11603] = 1'b1;  wr_cycle[11603] = 1'b0;  addr_rom[11603]='h00003014;  wr_data_rom[11603]='h00000000;
    rd_cycle[11604] = 1'b1;  wr_cycle[11604] = 1'b0;  addr_rom[11604]='h00001078;  wr_data_rom[11604]='h00000000;
    rd_cycle[11605] = 1'b0;  wr_cycle[11605] = 1'b1;  addr_rom[11605]='h000024c8;  wr_data_rom[11605]='h0000371b;
    rd_cycle[11606] = 1'b1;  wr_cycle[11606] = 1'b0;  addr_rom[11606]='h00002c2c;  wr_data_rom[11606]='h00000000;
    rd_cycle[11607] = 1'b1;  wr_cycle[11607] = 1'b0;  addr_rom[11607]='h00002058;  wr_data_rom[11607]='h00000000;
    rd_cycle[11608] = 1'b0;  wr_cycle[11608] = 1'b1;  addr_rom[11608]='h000028f4;  wr_data_rom[11608]='h000036c9;
    rd_cycle[11609] = 1'b0;  wr_cycle[11609] = 1'b1;  addr_rom[11609]='h0000251c;  wr_data_rom[11609]='h00001693;
    rd_cycle[11610] = 1'b0;  wr_cycle[11610] = 1'b1;  addr_rom[11610]='h00003b0c;  wr_data_rom[11610]='h00000666;
    rd_cycle[11611] = 1'b0;  wr_cycle[11611] = 1'b1;  addr_rom[11611]='h00001b30;  wr_data_rom[11611]='h00003534;
    rd_cycle[11612] = 1'b1;  wr_cycle[11612] = 1'b0;  addr_rom[11612]='h00003034;  wr_data_rom[11612]='h00000000;
    rd_cycle[11613] = 1'b0;  wr_cycle[11613] = 1'b1;  addr_rom[11613]='h00003368;  wr_data_rom[11613]='h00001b48;
    rd_cycle[11614] = 1'b1;  wr_cycle[11614] = 1'b0;  addr_rom[11614]='h000019c0;  wr_data_rom[11614]='h00000000;
    rd_cycle[11615] = 1'b0;  wr_cycle[11615] = 1'b1;  addr_rom[11615]='h0000347c;  wr_data_rom[11615]='h0000149f;
    rd_cycle[11616] = 1'b0;  wr_cycle[11616] = 1'b1;  addr_rom[11616]='h00002fcc;  wr_data_rom[11616]='h0000040c;
    rd_cycle[11617] = 1'b0;  wr_cycle[11617] = 1'b1;  addr_rom[11617]='h00003ae0;  wr_data_rom[11617]='h00000fba;
    rd_cycle[11618] = 1'b0;  wr_cycle[11618] = 1'b1;  addr_rom[11618]='h0000140c;  wr_data_rom[11618]='h00002979;
    rd_cycle[11619] = 1'b1;  wr_cycle[11619] = 1'b0;  addr_rom[11619]='h000007d4;  wr_data_rom[11619]='h00000000;
    rd_cycle[11620] = 1'b1;  wr_cycle[11620] = 1'b0;  addr_rom[11620]='h00001004;  wr_data_rom[11620]='h00000000;
    rd_cycle[11621] = 1'b0;  wr_cycle[11621] = 1'b1;  addr_rom[11621]='h00001ec8;  wr_data_rom[11621]='h00001e48;
    rd_cycle[11622] = 1'b1;  wr_cycle[11622] = 1'b0;  addr_rom[11622]='h000026b0;  wr_data_rom[11622]='h00000000;
    rd_cycle[11623] = 1'b1;  wr_cycle[11623] = 1'b0;  addr_rom[11623]='h000036a0;  wr_data_rom[11623]='h00000000;
    rd_cycle[11624] = 1'b1;  wr_cycle[11624] = 1'b0;  addr_rom[11624]='h000005cc;  wr_data_rom[11624]='h00000000;
    rd_cycle[11625] = 1'b1;  wr_cycle[11625] = 1'b0;  addr_rom[11625]='h00001f68;  wr_data_rom[11625]='h00000000;
    rd_cycle[11626] = 1'b0;  wr_cycle[11626] = 1'b1;  addr_rom[11626]='h00002ed8;  wr_data_rom[11626]='h00001043;
    rd_cycle[11627] = 1'b0;  wr_cycle[11627] = 1'b1;  addr_rom[11627]='h00001cb4;  wr_data_rom[11627]='h00002d1f;
    rd_cycle[11628] = 1'b0;  wr_cycle[11628] = 1'b1;  addr_rom[11628]='h000015c4;  wr_data_rom[11628]='h00001720;
    rd_cycle[11629] = 1'b0;  wr_cycle[11629] = 1'b1;  addr_rom[11629]='h000008f0;  wr_data_rom[11629]='h00000236;
    rd_cycle[11630] = 1'b1;  wr_cycle[11630] = 1'b0;  addr_rom[11630]='h00002460;  wr_data_rom[11630]='h00000000;
    rd_cycle[11631] = 1'b0;  wr_cycle[11631] = 1'b1;  addr_rom[11631]='h00002888;  wr_data_rom[11631]='h00000615;
    rd_cycle[11632] = 1'b1;  wr_cycle[11632] = 1'b0;  addr_rom[11632]='h000001d4;  wr_data_rom[11632]='h00000000;
    rd_cycle[11633] = 1'b1;  wr_cycle[11633] = 1'b0;  addr_rom[11633]='h00000314;  wr_data_rom[11633]='h00000000;
    rd_cycle[11634] = 1'b1;  wr_cycle[11634] = 1'b0;  addr_rom[11634]='h00001060;  wr_data_rom[11634]='h00000000;
    rd_cycle[11635] = 1'b1;  wr_cycle[11635] = 1'b0;  addr_rom[11635]='h0000131c;  wr_data_rom[11635]='h00000000;
    rd_cycle[11636] = 1'b0;  wr_cycle[11636] = 1'b1;  addr_rom[11636]='h00000d00;  wr_data_rom[11636]='h000019f1;
    rd_cycle[11637] = 1'b1;  wr_cycle[11637] = 1'b0;  addr_rom[11637]='h000026f0;  wr_data_rom[11637]='h00000000;
    rd_cycle[11638] = 1'b0;  wr_cycle[11638] = 1'b1;  addr_rom[11638]='h00003c98;  wr_data_rom[11638]='h00003491;
    rd_cycle[11639] = 1'b0;  wr_cycle[11639] = 1'b1;  addr_rom[11639]='h00003758;  wr_data_rom[11639]='h00002073;
    rd_cycle[11640] = 1'b1;  wr_cycle[11640] = 1'b0;  addr_rom[11640]='h0000004c;  wr_data_rom[11640]='h00000000;
    rd_cycle[11641] = 1'b0;  wr_cycle[11641] = 1'b1;  addr_rom[11641]='h00003300;  wr_data_rom[11641]='h00003fc9;
    rd_cycle[11642] = 1'b1;  wr_cycle[11642] = 1'b0;  addr_rom[11642]='h00002160;  wr_data_rom[11642]='h00000000;
    rd_cycle[11643] = 1'b1;  wr_cycle[11643] = 1'b0;  addr_rom[11643]='h000021e0;  wr_data_rom[11643]='h00000000;
    rd_cycle[11644] = 1'b1;  wr_cycle[11644] = 1'b0;  addr_rom[11644]='h00002160;  wr_data_rom[11644]='h00000000;
    rd_cycle[11645] = 1'b1;  wr_cycle[11645] = 1'b0;  addr_rom[11645]='h00001ee0;  wr_data_rom[11645]='h00000000;
    rd_cycle[11646] = 1'b1;  wr_cycle[11646] = 1'b0;  addr_rom[11646]='h00002c40;  wr_data_rom[11646]='h00000000;
    rd_cycle[11647] = 1'b0;  wr_cycle[11647] = 1'b1;  addr_rom[11647]='h000034c0;  wr_data_rom[11647]='h00002df7;
    rd_cycle[11648] = 1'b0;  wr_cycle[11648] = 1'b1;  addr_rom[11648]='h00003710;  wr_data_rom[11648]='h00003406;
    rd_cycle[11649] = 1'b0;  wr_cycle[11649] = 1'b1;  addr_rom[11649]='h00001b78;  wr_data_rom[11649]='h000007f9;
    rd_cycle[11650] = 1'b1;  wr_cycle[11650] = 1'b0;  addr_rom[11650]='h0000331c;  wr_data_rom[11650]='h00000000;
    rd_cycle[11651] = 1'b1;  wr_cycle[11651] = 1'b0;  addr_rom[11651]='h00002e6c;  wr_data_rom[11651]='h00000000;
    rd_cycle[11652] = 1'b0;  wr_cycle[11652] = 1'b1;  addr_rom[11652]='h00002c2c;  wr_data_rom[11652]='h00001b82;
    rd_cycle[11653] = 1'b0;  wr_cycle[11653] = 1'b1;  addr_rom[11653]='h000001b8;  wr_data_rom[11653]='h0000365b;
    rd_cycle[11654] = 1'b1;  wr_cycle[11654] = 1'b0;  addr_rom[11654]='h00002160;  wr_data_rom[11654]='h00000000;
    rd_cycle[11655] = 1'b1;  wr_cycle[11655] = 1'b0;  addr_rom[11655]='h00001064;  wr_data_rom[11655]='h00000000;
    rd_cycle[11656] = 1'b1;  wr_cycle[11656] = 1'b0;  addr_rom[11656]='h00001b24;  wr_data_rom[11656]='h00000000;
    rd_cycle[11657] = 1'b1;  wr_cycle[11657] = 1'b0;  addr_rom[11657]='h000008e0;  wr_data_rom[11657]='h00000000;
    rd_cycle[11658] = 1'b1;  wr_cycle[11658] = 1'b0;  addr_rom[11658]='h00003660;  wr_data_rom[11658]='h00000000;
    rd_cycle[11659] = 1'b1;  wr_cycle[11659] = 1'b0;  addr_rom[11659]='h00003b1c;  wr_data_rom[11659]='h00000000;
    rd_cycle[11660] = 1'b1;  wr_cycle[11660] = 1'b0;  addr_rom[11660]='h000029d8;  wr_data_rom[11660]='h00000000;
    rd_cycle[11661] = 1'b0;  wr_cycle[11661] = 1'b1;  addr_rom[11661]='h00003f04;  wr_data_rom[11661]='h00003cf7;
    rd_cycle[11662] = 1'b1;  wr_cycle[11662] = 1'b0;  addr_rom[11662]='h00003bb4;  wr_data_rom[11662]='h00000000;
    rd_cycle[11663] = 1'b0;  wr_cycle[11663] = 1'b1;  addr_rom[11663]='h00000484;  wr_data_rom[11663]='h00001f18;
    rd_cycle[11664] = 1'b1;  wr_cycle[11664] = 1'b0;  addr_rom[11664]='h00001b0c;  wr_data_rom[11664]='h00000000;
    rd_cycle[11665] = 1'b0;  wr_cycle[11665] = 1'b1;  addr_rom[11665]='h0000272c;  wr_data_rom[11665]='h00002e6c;
    rd_cycle[11666] = 1'b0;  wr_cycle[11666] = 1'b1;  addr_rom[11666]='h00002884;  wr_data_rom[11666]='h0000278d;
    rd_cycle[11667] = 1'b0;  wr_cycle[11667] = 1'b1;  addr_rom[11667]='h00001708;  wr_data_rom[11667]='h00002f06;
    rd_cycle[11668] = 1'b0;  wr_cycle[11668] = 1'b1;  addr_rom[11668]='h00002860;  wr_data_rom[11668]='h00002454;
    rd_cycle[11669] = 1'b0;  wr_cycle[11669] = 1'b1;  addr_rom[11669]='h00003458;  wr_data_rom[11669]='h000026bb;
    rd_cycle[11670] = 1'b0;  wr_cycle[11670] = 1'b1;  addr_rom[11670]='h000025ac;  wr_data_rom[11670]='h0000241f;
    rd_cycle[11671] = 1'b0;  wr_cycle[11671] = 1'b1;  addr_rom[11671]='h00000438;  wr_data_rom[11671]='h00000e9b;
    rd_cycle[11672] = 1'b1;  wr_cycle[11672] = 1'b0;  addr_rom[11672]='h00003234;  wr_data_rom[11672]='h00000000;
    rd_cycle[11673] = 1'b1;  wr_cycle[11673] = 1'b0;  addr_rom[11673]='h000002c4;  wr_data_rom[11673]='h00000000;
    rd_cycle[11674] = 1'b0;  wr_cycle[11674] = 1'b1;  addr_rom[11674]='h00000dbc;  wr_data_rom[11674]='h000000b5;
    rd_cycle[11675] = 1'b0;  wr_cycle[11675] = 1'b1;  addr_rom[11675]='h00000940;  wr_data_rom[11675]='h00003707;
    rd_cycle[11676] = 1'b1;  wr_cycle[11676] = 1'b0;  addr_rom[11676]='h00002d68;  wr_data_rom[11676]='h00000000;
    rd_cycle[11677] = 1'b0;  wr_cycle[11677] = 1'b1;  addr_rom[11677]='h00001e50;  wr_data_rom[11677]='h000015d8;
    rd_cycle[11678] = 1'b0;  wr_cycle[11678] = 1'b1;  addr_rom[11678]='h00002e84;  wr_data_rom[11678]='h00003248;
    rd_cycle[11679] = 1'b1;  wr_cycle[11679] = 1'b0;  addr_rom[11679]='h00000934;  wr_data_rom[11679]='h00000000;
    rd_cycle[11680] = 1'b0;  wr_cycle[11680] = 1'b1;  addr_rom[11680]='h0000189c;  wr_data_rom[11680]='h00002b4d;
    rd_cycle[11681] = 1'b1;  wr_cycle[11681] = 1'b0;  addr_rom[11681]='h00001958;  wr_data_rom[11681]='h00000000;
    rd_cycle[11682] = 1'b0;  wr_cycle[11682] = 1'b1;  addr_rom[11682]='h00003f48;  wr_data_rom[11682]='h00002573;
    rd_cycle[11683] = 1'b0;  wr_cycle[11683] = 1'b1;  addr_rom[11683]='h00002a4c;  wr_data_rom[11683]='h0000103c;
    rd_cycle[11684] = 1'b0;  wr_cycle[11684] = 1'b1;  addr_rom[11684]='h0000247c;  wr_data_rom[11684]='h0000365d;
    rd_cycle[11685] = 1'b1;  wr_cycle[11685] = 1'b0;  addr_rom[11685]='h00000fe8;  wr_data_rom[11685]='h00000000;
    rd_cycle[11686] = 1'b1;  wr_cycle[11686] = 1'b0;  addr_rom[11686]='h00000c6c;  wr_data_rom[11686]='h00000000;
    rd_cycle[11687] = 1'b0;  wr_cycle[11687] = 1'b1;  addr_rom[11687]='h00001528;  wr_data_rom[11687]='h00001098;
    rd_cycle[11688] = 1'b1;  wr_cycle[11688] = 1'b0;  addr_rom[11688]='h0000171c;  wr_data_rom[11688]='h00000000;
    rd_cycle[11689] = 1'b0;  wr_cycle[11689] = 1'b1;  addr_rom[11689]='h00003f78;  wr_data_rom[11689]='h00000211;
    rd_cycle[11690] = 1'b1;  wr_cycle[11690] = 1'b0;  addr_rom[11690]='h000030c0;  wr_data_rom[11690]='h00000000;
    rd_cycle[11691] = 1'b1;  wr_cycle[11691] = 1'b0;  addr_rom[11691]='h00001e6c;  wr_data_rom[11691]='h00000000;
    rd_cycle[11692] = 1'b1;  wr_cycle[11692] = 1'b0;  addr_rom[11692]='h000011d8;  wr_data_rom[11692]='h00000000;
    rd_cycle[11693] = 1'b1;  wr_cycle[11693] = 1'b0;  addr_rom[11693]='h00001c18;  wr_data_rom[11693]='h00000000;
    rd_cycle[11694] = 1'b0;  wr_cycle[11694] = 1'b1;  addr_rom[11694]='h00001954;  wr_data_rom[11694]='h00002ba5;
    rd_cycle[11695] = 1'b1;  wr_cycle[11695] = 1'b0;  addr_rom[11695]='h000025f0;  wr_data_rom[11695]='h00000000;
    rd_cycle[11696] = 1'b1;  wr_cycle[11696] = 1'b0;  addr_rom[11696]='h00002f6c;  wr_data_rom[11696]='h00000000;
    rd_cycle[11697] = 1'b1;  wr_cycle[11697] = 1'b0;  addr_rom[11697]='h00003f5c;  wr_data_rom[11697]='h00000000;
    rd_cycle[11698] = 1'b0;  wr_cycle[11698] = 1'b1;  addr_rom[11698]='h0000218c;  wr_data_rom[11698]='h000014d0;
    rd_cycle[11699] = 1'b1;  wr_cycle[11699] = 1'b0;  addr_rom[11699]='h00001408;  wr_data_rom[11699]='h00000000;
    rd_cycle[11700] = 1'b1;  wr_cycle[11700] = 1'b0;  addr_rom[11700]='h00001c40;  wr_data_rom[11700]='h00000000;
    rd_cycle[11701] = 1'b0;  wr_cycle[11701] = 1'b1;  addr_rom[11701]='h00002a24;  wr_data_rom[11701]='h00002a47;
    rd_cycle[11702] = 1'b1;  wr_cycle[11702] = 1'b0;  addr_rom[11702]='h00001428;  wr_data_rom[11702]='h00000000;
    rd_cycle[11703] = 1'b0;  wr_cycle[11703] = 1'b1;  addr_rom[11703]='h00000d68;  wr_data_rom[11703]='h00000602;
    rd_cycle[11704] = 1'b1;  wr_cycle[11704] = 1'b0;  addr_rom[11704]='h00001844;  wr_data_rom[11704]='h00000000;
    rd_cycle[11705] = 1'b0;  wr_cycle[11705] = 1'b1;  addr_rom[11705]='h000030c8;  wr_data_rom[11705]='h00003ea2;
    rd_cycle[11706] = 1'b0;  wr_cycle[11706] = 1'b1;  addr_rom[11706]='h00000c80;  wr_data_rom[11706]='h00001808;
    rd_cycle[11707] = 1'b0;  wr_cycle[11707] = 1'b1;  addr_rom[11707]='h00003460;  wr_data_rom[11707]='h0000037a;
    rd_cycle[11708] = 1'b0;  wr_cycle[11708] = 1'b1;  addr_rom[11708]='h00002654;  wr_data_rom[11708]='h0000341d;
    rd_cycle[11709] = 1'b1;  wr_cycle[11709] = 1'b0;  addr_rom[11709]='h00002c9c;  wr_data_rom[11709]='h00000000;
    rd_cycle[11710] = 1'b1;  wr_cycle[11710] = 1'b0;  addr_rom[11710]='h00002680;  wr_data_rom[11710]='h00000000;
    rd_cycle[11711] = 1'b0;  wr_cycle[11711] = 1'b1;  addr_rom[11711]='h00002fe4;  wr_data_rom[11711]='h0000377e;
    rd_cycle[11712] = 1'b0;  wr_cycle[11712] = 1'b1;  addr_rom[11712]='h00001508;  wr_data_rom[11712]='h00001b5c;
    rd_cycle[11713] = 1'b0;  wr_cycle[11713] = 1'b1;  addr_rom[11713]='h000022a4;  wr_data_rom[11713]='h00000796;
    rd_cycle[11714] = 1'b1;  wr_cycle[11714] = 1'b0;  addr_rom[11714]='h00003834;  wr_data_rom[11714]='h00000000;
    rd_cycle[11715] = 1'b1;  wr_cycle[11715] = 1'b0;  addr_rom[11715]='h000035f8;  wr_data_rom[11715]='h00000000;
    rd_cycle[11716] = 1'b0;  wr_cycle[11716] = 1'b1;  addr_rom[11716]='h00001864;  wr_data_rom[11716]='h00002c16;
    rd_cycle[11717] = 1'b0;  wr_cycle[11717] = 1'b1;  addr_rom[11717]='h000009b4;  wr_data_rom[11717]='h0000070a;
    rd_cycle[11718] = 1'b1;  wr_cycle[11718] = 1'b0;  addr_rom[11718]='h00000d54;  wr_data_rom[11718]='h00000000;
    rd_cycle[11719] = 1'b0;  wr_cycle[11719] = 1'b1;  addr_rom[11719]='h00001c90;  wr_data_rom[11719]='h0000314a;
    rd_cycle[11720] = 1'b1;  wr_cycle[11720] = 1'b0;  addr_rom[11720]='h0000276c;  wr_data_rom[11720]='h00000000;
    rd_cycle[11721] = 1'b0;  wr_cycle[11721] = 1'b1;  addr_rom[11721]='h00001b20;  wr_data_rom[11721]='h00000241;
    rd_cycle[11722] = 1'b1;  wr_cycle[11722] = 1'b0;  addr_rom[11722]='h000023a8;  wr_data_rom[11722]='h00000000;
    rd_cycle[11723] = 1'b0;  wr_cycle[11723] = 1'b1;  addr_rom[11723]='h00003b70;  wr_data_rom[11723]='h000031c7;
    rd_cycle[11724] = 1'b1;  wr_cycle[11724] = 1'b0;  addr_rom[11724]='h00000960;  wr_data_rom[11724]='h00000000;
    rd_cycle[11725] = 1'b0;  wr_cycle[11725] = 1'b1;  addr_rom[11725]='h0000296c;  wr_data_rom[11725]='h000020bc;
    rd_cycle[11726] = 1'b1;  wr_cycle[11726] = 1'b0;  addr_rom[11726]='h00001f54;  wr_data_rom[11726]='h00000000;
    rd_cycle[11727] = 1'b0;  wr_cycle[11727] = 1'b1;  addr_rom[11727]='h0000154c;  wr_data_rom[11727]='h00002716;
    rd_cycle[11728] = 1'b1;  wr_cycle[11728] = 1'b0;  addr_rom[11728]='h00003574;  wr_data_rom[11728]='h00000000;
    rd_cycle[11729] = 1'b0;  wr_cycle[11729] = 1'b1;  addr_rom[11729]='h00003dc0;  wr_data_rom[11729]='h000036b3;
    rd_cycle[11730] = 1'b1;  wr_cycle[11730] = 1'b0;  addr_rom[11730]='h00003f04;  wr_data_rom[11730]='h00000000;
    rd_cycle[11731] = 1'b0;  wr_cycle[11731] = 1'b1;  addr_rom[11731]='h00000d00;  wr_data_rom[11731]='h0000232a;
    rd_cycle[11732] = 1'b0;  wr_cycle[11732] = 1'b1;  addr_rom[11732]='h00001d00;  wr_data_rom[11732]='h000007bb;
    rd_cycle[11733] = 1'b1;  wr_cycle[11733] = 1'b0;  addr_rom[11733]='h00003cf4;  wr_data_rom[11733]='h00000000;
    rd_cycle[11734] = 1'b0;  wr_cycle[11734] = 1'b1;  addr_rom[11734]='h00002110;  wr_data_rom[11734]='h00003dbc;
    rd_cycle[11735] = 1'b1;  wr_cycle[11735] = 1'b0;  addr_rom[11735]='h0000171c;  wr_data_rom[11735]='h00000000;
    rd_cycle[11736] = 1'b1;  wr_cycle[11736] = 1'b0;  addr_rom[11736]='h00003720;  wr_data_rom[11736]='h00000000;
    rd_cycle[11737] = 1'b1;  wr_cycle[11737] = 1'b0;  addr_rom[11737]='h00002b24;  wr_data_rom[11737]='h00000000;
    rd_cycle[11738] = 1'b1;  wr_cycle[11738] = 1'b0;  addr_rom[11738]='h00002318;  wr_data_rom[11738]='h00000000;
    rd_cycle[11739] = 1'b1;  wr_cycle[11739] = 1'b0;  addr_rom[11739]='h000004bc;  wr_data_rom[11739]='h00000000;
    rd_cycle[11740] = 1'b0;  wr_cycle[11740] = 1'b1;  addr_rom[11740]='h000034d4;  wr_data_rom[11740]='h00002e25;
    rd_cycle[11741] = 1'b1;  wr_cycle[11741] = 1'b0;  addr_rom[11741]='h00001a54;  wr_data_rom[11741]='h00000000;
    rd_cycle[11742] = 1'b0;  wr_cycle[11742] = 1'b1;  addr_rom[11742]='h00003ca0;  wr_data_rom[11742]='h00003db5;
    rd_cycle[11743] = 1'b0;  wr_cycle[11743] = 1'b1;  addr_rom[11743]='h000038d8;  wr_data_rom[11743]='h00000e3e;
    rd_cycle[11744] = 1'b0;  wr_cycle[11744] = 1'b1;  addr_rom[11744]='h00001254;  wr_data_rom[11744]='h000019a4;
    rd_cycle[11745] = 1'b0;  wr_cycle[11745] = 1'b1;  addr_rom[11745]='h00003e9c;  wr_data_rom[11745]='h00000aec;
    rd_cycle[11746] = 1'b1;  wr_cycle[11746] = 1'b0;  addr_rom[11746]='h000003a0;  wr_data_rom[11746]='h00000000;
    rd_cycle[11747] = 1'b1;  wr_cycle[11747] = 1'b0;  addr_rom[11747]='h00001770;  wr_data_rom[11747]='h00000000;
    rd_cycle[11748] = 1'b0;  wr_cycle[11748] = 1'b1;  addr_rom[11748]='h00001370;  wr_data_rom[11748]='h000015b5;
    rd_cycle[11749] = 1'b0;  wr_cycle[11749] = 1'b1;  addr_rom[11749]='h00003664;  wr_data_rom[11749]='h0000369f;
    rd_cycle[11750] = 1'b1;  wr_cycle[11750] = 1'b0;  addr_rom[11750]='h000024dc;  wr_data_rom[11750]='h00000000;
    rd_cycle[11751] = 1'b0;  wr_cycle[11751] = 1'b1;  addr_rom[11751]='h00002614;  wr_data_rom[11751]='h00000efa;
    rd_cycle[11752] = 1'b1;  wr_cycle[11752] = 1'b0;  addr_rom[11752]='h0000157c;  wr_data_rom[11752]='h00000000;
    rd_cycle[11753] = 1'b0;  wr_cycle[11753] = 1'b1;  addr_rom[11753]='h00000308;  wr_data_rom[11753]='h00002431;
    rd_cycle[11754] = 1'b1;  wr_cycle[11754] = 1'b0;  addr_rom[11754]='h00003b6c;  wr_data_rom[11754]='h00000000;
    rd_cycle[11755] = 1'b0;  wr_cycle[11755] = 1'b1;  addr_rom[11755]='h00001d44;  wr_data_rom[11755]='h000009c4;
    rd_cycle[11756] = 1'b1;  wr_cycle[11756] = 1'b0;  addr_rom[11756]='h00003dd4;  wr_data_rom[11756]='h00000000;
    rd_cycle[11757] = 1'b0;  wr_cycle[11757] = 1'b1;  addr_rom[11757]='h00002610;  wr_data_rom[11757]='h00000d1d;
    rd_cycle[11758] = 1'b1;  wr_cycle[11758] = 1'b0;  addr_rom[11758]='h00002888;  wr_data_rom[11758]='h00000000;
    rd_cycle[11759] = 1'b1;  wr_cycle[11759] = 1'b0;  addr_rom[11759]='h00001394;  wr_data_rom[11759]='h00000000;
    rd_cycle[11760] = 1'b1;  wr_cycle[11760] = 1'b0;  addr_rom[11760]='h0000365c;  wr_data_rom[11760]='h00000000;
    rd_cycle[11761] = 1'b1;  wr_cycle[11761] = 1'b0;  addr_rom[11761]='h00000688;  wr_data_rom[11761]='h00000000;
    rd_cycle[11762] = 1'b0;  wr_cycle[11762] = 1'b1;  addr_rom[11762]='h00002978;  wr_data_rom[11762]='h00002620;
    rd_cycle[11763] = 1'b0;  wr_cycle[11763] = 1'b1;  addr_rom[11763]='h00003e6c;  wr_data_rom[11763]='h00001bab;
    rd_cycle[11764] = 1'b0;  wr_cycle[11764] = 1'b1;  addr_rom[11764]='h00000c00;  wr_data_rom[11764]='h00003db4;
    rd_cycle[11765] = 1'b0;  wr_cycle[11765] = 1'b1;  addr_rom[11765]='h00003718;  wr_data_rom[11765]='h00000928;
    rd_cycle[11766] = 1'b0;  wr_cycle[11766] = 1'b1;  addr_rom[11766]='h000015ec;  wr_data_rom[11766]='h00003122;
    rd_cycle[11767] = 1'b1;  wr_cycle[11767] = 1'b0;  addr_rom[11767]='h0000370c;  wr_data_rom[11767]='h00000000;
    rd_cycle[11768] = 1'b1;  wr_cycle[11768] = 1'b0;  addr_rom[11768]='h00000c5c;  wr_data_rom[11768]='h00000000;
    rd_cycle[11769] = 1'b0;  wr_cycle[11769] = 1'b1;  addr_rom[11769]='h00001b04;  wr_data_rom[11769]='h0000070e;
    rd_cycle[11770] = 1'b1;  wr_cycle[11770] = 1'b0;  addr_rom[11770]='h000009f4;  wr_data_rom[11770]='h00000000;
    rd_cycle[11771] = 1'b1;  wr_cycle[11771] = 1'b0;  addr_rom[11771]='h00003dd4;  wr_data_rom[11771]='h00000000;
    rd_cycle[11772] = 1'b1;  wr_cycle[11772] = 1'b0;  addr_rom[11772]='h00002bec;  wr_data_rom[11772]='h00000000;
    rd_cycle[11773] = 1'b1;  wr_cycle[11773] = 1'b0;  addr_rom[11773]='h000011b4;  wr_data_rom[11773]='h00000000;
    rd_cycle[11774] = 1'b0;  wr_cycle[11774] = 1'b1;  addr_rom[11774]='h00001f78;  wr_data_rom[11774]='h000030a0;
    rd_cycle[11775] = 1'b0;  wr_cycle[11775] = 1'b1;  addr_rom[11775]='h000014f4;  wr_data_rom[11775]='h000013df;
    rd_cycle[11776] = 1'b1;  wr_cycle[11776] = 1'b0;  addr_rom[11776]='h000038fc;  wr_data_rom[11776]='h00000000;
    rd_cycle[11777] = 1'b1;  wr_cycle[11777] = 1'b0;  addr_rom[11777]='h00001a68;  wr_data_rom[11777]='h00000000;
    rd_cycle[11778] = 1'b1;  wr_cycle[11778] = 1'b0;  addr_rom[11778]='h00001d00;  wr_data_rom[11778]='h00000000;
    rd_cycle[11779] = 1'b1;  wr_cycle[11779] = 1'b0;  addr_rom[11779]='h00001160;  wr_data_rom[11779]='h00000000;
    rd_cycle[11780] = 1'b0;  wr_cycle[11780] = 1'b1;  addr_rom[11780]='h00000634;  wr_data_rom[11780]='h00000211;
    rd_cycle[11781] = 1'b1;  wr_cycle[11781] = 1'b0;  addr_rom[11781]='h00002244;  wr_data_rom[11781]='h00000000;
    rd_cycle[11782] = 1'b0;  wr_cycle[11782] = 1'b1;  addr_rom[11782]='h00001b08;  wr_data_rom[11782]='h000029eb;
    rd_cycle[11783] = 1'b1;  wr_cycle[11783] = 1'b0;  addr_rom[11783]='h00003fac;  wr_data_rom[11783]='h00000000;
    rd_cycle[11784] = 1'b1;  wr_cycle[11784] = 1'b0;  addr_rom[11784]='h00000a8c;  wr_data_rom[11784]='h00000000;
    rd_cycle[11785] = 1'b0;  wr_cycle[11785] = 1'b1;  addr_rom[11785]='h00001200;  wr_data_rom[11785]='h00002fd5;
    rd_cycle[11786] = 1'b1;  wr_cycle[11786] = 1'b0;  addr_rom[11786]='h00003120;  wr_data_rom[11786]='h00000000;
    rd_cycle[11787] = 1'b1;  wr_cycle[11787] = 1'b0;  addr_rom[11787]='h00002288;  wr_data_rom[11787]='h00000000;
    rd_cycle[11788] = 1'b0;  wr_cycle[11788] = 1'b1;  addr_rom[11788]='h0000164c;  wr_data_rom[11788]='h00003ee5;
    rd_cycle[11789] = 1'b1;  wr_cycle[11789] = 1'b0;  addr_rom[11789]='h00000338;  wr_data_rom[11789]='h00000000;
    rd_cycle[11790] = 1'b0;  wr_cycle[11790] = 1'b1;  addr_rom[11790]='h000022ec;  wr_data_rom[11790]='h00000991;
    rd_cycle[11791] = 1'b1;  wr_cycle[11791] = 1'b0;  addr_rom[11791]='h0000151c;  wr_data_rom[11791]='h00000000;
    rd_cycle[11792] = 1'b0;  wr_cycle[11792] = 1'b1;  addr_rom[11792]='h00003d3c;  wr_data_rom[11792]='h000023bf;
    rd_cycle[11793] = 1'b1;  wr_cycle[11793] = 1'b0;  addr_rom[11793]='h0000241c;  wr_data_rom[11793]='h00000000;
    rd_cycle[11794] = 1'b1;  wr_cycle[11794] = 1'b0;  addr_rom[11794]='h00003fe8;  wr_data_rom[11794]='h00000000;
    rd_cycle[11795] = 1'b0;  wr_cycle[11795] = 1'b1;  addr_rom[11795]='h000026f8;  wr_data_rom[11795]='h00000a23;
    rd_cycle[11796] = 1'b1;  wr_cycle[11796] = 1'b0;  addr_rom[11796]='h000006d0;  wr_data_rom[11796]='h00000000;
    rd_cycle[11797] = 1'b0;  wr_cycle[11797] = 1'b1;  addr_rom[11797]='h0000353c;  wr_data_rom[11797]='h0000303f;
    rd_cycle[11798] = 1'b1;  wr_cycle[11798] = 1'b0;  addr_rom[11798]='h00000200;  wr_data_rom[11798]='h00000000;
    rd_cycle[11799] = 1'b1;  wr_cycle[11799] = 1'b0;  addr_rom[11799]='h000005e4;  wr_data_rom[11799]='h00000000;
    rd_cycle[11800] = 1'b1;  wr_cycle[11800] = 1'b0;  addr_rom[11800]='h00003504;  wr_data_rom[11800]='h00000000;
    rd_cycle[11801] = 1'b0;  wr_cycle[11801] = 1'b1;  addr_rom[11801]='h00000bc4;  wr_data_rom[11801]='h00001ea7;
    rd_cycle[11802] = 1'b1;  wr_cycle[11802] = 1'b0;  addr_rom[11802]='h000024f0;  wr_data_rom[11802]='h00000000;
    rd_cycle[11803] = 1'b1;  wr_cycle[11803] = 1'b0;  addr_rom[11803]='h00002264;  wr_data_rom[11803]='h00000000;
    rd_cycle[11804] = 1'b1;  wr_cycle[11804] = 1'b0;  addr_rom[11804]='h00000430;  wr_data_rom[11804]='h00000000;
    rd_cycle[11805] = 1'b0;  wr_cycle[11805] = 1'b1;  addr_rom[11805]='h00003be4;  wr_data_rom[11805]='h00000d3c;
    rd_cycle[11806] = 1'b1;  wr_cycle[11806] = 1'b0;  addr_rom[11806]='h00003be0;  wr_data_rom[11806]='h00000000;
    rd_cycle[11807] = 1'b0;  wr_cycle[11807] = 1'b1;  addr_rom[11807]='h00003b08;  wr_data_rom[11807]='h00002675;
    rd_cycle[11808] = 1'b0;  wr_cycle[11808] = 1'b1;  addr_rom[11808]='h000010e4;  wr_data_rom[11808]='h00001a5d;
    rd_cycle[11809] = 1'b1;  wr_cycle[11809] = 1'b0;  addr_rom[11809]='h00002cdc;  wr_data_rom[11809]='h00000000;
    rd_cycle[11810] = 1'b0;  wr_cycle[11810] = 1'b1;  addr_rom[11810]='h00002258;  wr_data_rom[11810]='h00003acb;
    rd_cycle[11811] = 1'b1;  wr_cycle[11811] = 1'b0;  addr_rom[11811]='h0000126c;  wr_data_rom[11811]='h00000000;
    rd_cycle[11812] = 1'b0;  wr_cycle[11812] = 1'b1;  addr_rom[11812]='h00002ed0;  wr_data_rom[11812]='h000017fc;
    rd_cycle[11813] = 1'b1;  wr_cycle[11813] = 1'b0;  addr_rom[11813]='h00001bac;  wr_data_rom[11813]='h00000000;
    rd_cycle[11814] = 1'b1;  wr_cycle[11814] = 1'b0;  addr_rom[11814]='h0000023c;  wr_data_rom[11814]='h00000000;
    rd_cycle[11815] = 1'b0;  wr_cycle[11815] = 1'b1;  addr_rom[11815]='h00001000;  wr_data_rom[11815]='h00000760;
    rd_cycle[11816] = 1'b0;  wr_cycle[11816] = 1'b1;  addr_rom[11816]='h00000994;  wr_data_rom[11816]='h00003161;
    rd_cycle[11817] = 1'b0;  wr_cycle[11817] = 1'b1;  addr_rom[11817]='h00000a5c;  wr_data_rom[11817]='h00001414;
    rd_cycle[11818] = 1'b1;  wr_cycle[11818] = 1'b0;  addr_rom[11818]='h000029c8;  wr_data_rom[11818]='h00000000;
    rd_cycle[11819] = 1'b1;  wr_cycle[11819] = 1'b0;  addr_rom[11819]='h00002af4;  wr_data_rom[11819]='h00000000;
    rd_cycle[11820] = 1'b1;  wr_cycle[11820] = 1'b0;  addr_rom[11820]='h00001c7c;  wr_data_rom[11820]='h00000000;
    rd_cycle[11821] = 1'b1;  wr_cycle[11821] = 1'b0;  addr_rom[11821]='h0000265c;  wr_data_rom[11821]='h00000000;
    rd_cycle[11822] = 1'b1;  wr_cycle[11822] = 1'b0;  addr_rom[11822]='h00003b48;  wr_data_rom[11822]='h00000000;
    rd_cycle[11823] = 1'b0;  wr_cycle[11823] = 1'b1;  addr_rom[11823]='h00001ca4;  wr_data_rom[11823]='h000030b6;
    rd_cycle[11824] = 1'b1;  wr_cycle[11824] = 1'b0;  addr_rom[11824]='h00001a14;  wr_data_rom[11824]='h00000000;
    rd_cycle[11825] = 1'b1;  wr_cycle[11825] = 1'b0;  addr_rom[11825]='h00002b50;  wr_data_rom[11825]='h00000000;
    rd_cycle[11826] = 1'b1;  wr_cycle[11826] = 1'b0;  addr_rom[11826]='h00002bc0;  wr_data_rom[11826]='h00000000;
    rd_cycle[11827] = 1'b0;  wr_cycle[11827] = 1'b1;  addr_rom[11827]='h00003bac;  wr_data_rom[11827]='h00002a2d;
    rd_cycle[11828] = 1'b0;  wr_cycle[11828] = 1'b1;  addr_rom[11828]='h000005e8;  wr_data_rom[11828]='h00000e76;
    rd_cycle[11829] = 1'b0;  wr_cycle[11829] = 1'b1;  addr_rom[11829]='h00003160;  wr_data_rom[11829]='h00003395;
    rd_cycle[11830] = 1'b0;  wr_cycle[11830] = 1'b1;  addr_rom[11830]='h00000088;  wr_data_rom[11830]='h000031ff;
    rd_cycle[11831] = 1'b1;  wr_cycle[11831] = 1'b0;  addr_rom[11831]='h0000058c;  wr_data_rom[11831]='h00000000;
    rd_cycle[11832] = 1'b0;  wr_cycle[11832] = 1'b1;  addr_rom[11832]='h00001dec;  wr_data_rom[11832]='h000026c3;
    rd_cycle[11833] = 1'b0;  wr_cycle[11833] = 1'b1;  addr_rom[11833]='h00003da0;  wr_data_rom[11833]='h00000bbc;
    rd_cycle[11834] = 1'b1;  wr_cycle[11834] = 1'b0;  addr_rom[11834]='h000002ac;  wr_data_rom[11834]='h00000000;
    rd_cycle[11835] = 1'b1;  wr_cycle[11835] = 1'b0;  addr_rom[11835]='h00001070;  wr_data_rom[11835]='h00000000;
    rd_cycle[11836] = 1'b1;  wr_cycle[11836] = 1'b0;  addr_rom[11836]='h00003918;  wr_data_rom[11836]='h00000000;
    rd_cycle[11837] = 1'b1;  wr_cycle[11837] = 1'b0;  addr_rom[11837]='h000012fc;  wr_data_rom[11837]='h00000000;
    rd_cycle[11838] = 1'b1;  wr_cycle[11838] = 1'b0;  addr_rom[11838]='h00001c4c;  wr_data_rom[11838]='h00000000;
    rd_cycle[11839] = 1'b1;  wr_cycle[11839] = 1'b0;  addr_rom[11839]='h00003c20;  wr_data_rom[11839]='h00000000;
    rd_cycle[11840] = 1'b1;  wr_cycle[11840] = 1'b0;  addr_rom[11840]='h00001764;  wr_data_rom[11840]='h00000000;
    rd_cycle[11841] = 1'b1;  wr_cycle[11841] = 1'b0;  addr_rom[11841]='h00003dd4;  wr_data_rom[11841]='h00000000;
    rd_cycle[11842] = 1'b1;  wr_cycle[11842] = 1'b0;  addr_rom[11842]='h00001320;  wr_data_rom[11842]='h00000000;
    rd_cycle[11843] = 1'b0;  wr_cycle[11843] = 1'b1;  addr_rom[11843]='h000004f0;  wr_data_rom[11843]='h00003d73;
    rd_cycle[11844] = 1'b1;  wr_cycle[11844] = 1'b0;  addr_rom[11844]='h00003f20;  wr_data_rom[11844]='h00000000;
    rd_cycle[11845] = 1'b0;  wr_cycle[11845] = 1'b1;  addr_rom[11845]='h000022c8;  wr_data_rom[11845]='h00002e80;
    rd_cycle[11846] = 1'b1;  wr_cycle[11846] = 1'b0;  addr_rom[11846]='h00000934;  wr_data_rom[11846]='h00000000;
    rd_cycle[11847] = 1'b0;  wr_cycle[11847] = 1'b1;  addr_rom[11847]='h00003d3c;  wr_data_rom[11847]='h000031c2;
    rd_cycle[11848] = 1'b0;  wr_cycle[11848] = 1'b1;  addr_rom[11848]='h00001fc8;  wr_data_rom[11848]='h000030d9;
    rd_cycle[11849] = 1'b0;  wr_cycle[11849] = 1'b1;  addr_rom[11849]='h00000498;  wr_data_rom[11849]='h000003d5;
    rd_cycle[11850] = 1'b1;  wr_cycle[11850] = 1'b0;  addr_rom[11850]='h00002cd8;  wr_data_rom[11850]='h00000000;
    rd_cycle[11851] = 1'b0;  wr_cycle[11851] = 1'b1;  addr_rom[11851]='h00002008;  wr_data_rom[11851]='h00001950;
    rd_cycle[11852] = 1'b1;  wr_cycle[11852] = 1'b0;  addr_rom[11852]='h000031ec;  wr_data_rom[11852]='h00000000;
    rd_cycle[11853] = 1'b1;  wr_cycle[11853] = 1'b0;  addr_rom[11853]='h00001cb0;  wr_data_rom[11853]='h00000000;
    rd_cycle[11854] = 1'b0;  wr_cycle[11854] = 1'b1;  addr_rom[11854]='h000031e0;  wr_data_rom[11854]='h000009a6;
    rd_cycle[11855] = 1'b1;  wr_cycle[11855] = 1'b0;  addr_rom[11855]='h00002e80;  wr_data_rom[11855]='h00000000;
    rd_cycle[11856] = 1'b0;  wr_cycle[11856] = 1'b1;  addr_rom[11856]='h000022ec;  wr_data_rom[11856]='h0000360f;
    rd_cycle[11857] = 1'b0;  wr_cycle[11857] = 1'b1;  addr_rom[11857]='h00000b4c;  wr_data_rom[11857]='h00000a33;
    rd_cycle[11858] = 1'b0;  wr_cycle[11858] = 1'b1;  addr_rom[11858]='h000026b4;  wr_data_rom[11858]='h00000629;
    rd_cycle[11859] = 1'b1;  wr_cycle[11859] = 1'b0;  addr_rom[11859]='h00003034;  wr_data_rom[11859]='h00000000;
    rd_cycle[11860] = 1'b1;  wr_cycle[11860] = 1'b0;  addr_rom[11860]='h000019b4;  wr_data_rom[11860]='h00000000;
    rd_cycle[11861] = 1'b0;  wr_cycle[11861] = 1'b1;  addr_rom[11861]='h000033f0;  wr_data_rom[11861]='h0000336f;
    rd_cycle[11862] = 1'b0;  wr_cycle[11862] = 1'b1;  addr_rom[11862]='h0000132c;  wr_data_rom[11862]='h000010d5;
    rd_cycle[11863] = 1'b0;  wr_cycle[11863] = 1'b1;  addr_rom[11863]='h00002ba0;  wr_data_rom[11863]='h000034a3;
    rd_cycle[11864] = 1'b0;  wr_cycle[11864] = 1'b1;  addr_rom[11864]='h0000263c;  wr_data_rom[11864]='h000036b4;
    rd_cycle[11865] = 1'b0;  wr_cycle[11865] = 1'b1;  addr_rom[11865]='h00002ff4;  wr_data_rom[11865]='h00003b72;
    rd_cycle[11866] = 1'b0;  wr_cycle[11866] = 1'b1;  addr_rom[11866]='h00000610;  wr_data_rom[11866]='h0000087e;
    rd_cycle[11867] = 1'b1;  wr_cycle[11867] = 1'b0;  addr_rom[11867]='h00001190;  wr_data_rom[11867]='h00000000;
    rd_cycle[11868] = 1'b0;  wr_cycle[11868] = 1'b1;  addr_rom[11868]='h0000004c;  wr_data_rom[11868]='h00002b1a;
    rd_cycle[11869] = 1'b0;  wr_cycle[11869] = 1'b1;  addr_rom[11869]='h000017c4;  wr_data_rom[11869]='h00000b68;
    rd_cycle[11870] = 1'b0;  wr_cycle[11870] = 1'b1;  addr_rom[11870]='h00003928;  wr_data_rom[11870]='h000003fa;
    rd_cycle[11871] = 1'b0;  wr_cycle[11871] = 1'b1;  addr_rom[11871]='h00001be8;  wr_data_rom[11871]='h00001c2b;
    rd_cycle[11872] = 1'b0;  wr_cycle[11872] = 1'b1;  addr_rom[11872]='h00000338;  wr_data_rom[11872]='h00000702;
    rd_cycle[11873] = 1'b0;  wr_cycle[11873] = 1'b1;  addr_rom[11873]='h00000834;  wr_data_rom[11873]='h00000fb5;
    rd_cycle[11874] = 1'b1;  wr_cycle[11874] = 1'b0;  addr_rom[11874]='h00000894;  wr_data_rom[11874]='h00000000;
    rd_cycle[11875] = 1'b0;  wr_cycle[11875] = 1'b1;  addr_rom[11875]='h00000f9c;  wr_data_rom[11875]='h00002b2c;
    rd_cycle[11876] = 1'b0;  wr_cycle[11876] = 1'b1;  addr_rom[11876]='h0000219c;  wr_data_rom[11876]='h00003ec6;
    rd_cycle[11877] = 1'b1;  wr_cycle[11877] = 1'b0;  addr_rom[11877]='h00003780;  wr_data_rom[11877]='h00000000;
    rd_cycle[11878] = 1'b0;  wr_cycle[11878] = 1'b1;  addr_rom[11878]='h00003c90;  wr_data_rom[11878]='h0000369f;
    rd_cycle[11879] = 1'b0;  wr_cycle[11879] = 1'b1;  addr_rom[11879]='h00000404;  wr_data_rom[11879]='h00000c8a;
    rd_cycle[11880] = 1'b1;  wr_cycle[11880] = 1'b0;  addr_rom[11880]='h00000178;  wr_data_rom[11880]='h00000000;
    rd_cycle[11881] = 1'b0;  wr_cycle[11881] = 1'b1;  addr_rom[11881]='h00000bd4;  wr_data_rom[11881]='h00003fdf;
    rd_cycle[11882] = 1'b0;  wr_cycle[11882] = 1'b1;  addr_rom[11882]='h000005f8;  wr_data_rom[11882]='h00001275;
    rd_cycle[11883] = 1'b1;  wr_cycle[11883] = 1'b0;  addr_rom[11883]='h00002158;  wr_data_rom[11883]='h00000000;
    rd_cycle[11884] = 1'b0;  wr_cycle[11884] = 1'b1;  addr_rom[11884]='h000004d4;  wr_data_rom[11884]='h000032eb;
    rd_cycle[11885] = 1'b1;  wr_cycle[11885] = 1'b0;  addr_rom[11885]='h00001dfc;  wr_data_rom[11885]='h00000000;
    rd_cycle[11886] = 1'b0;  wr_cycle[11886] = 1'b1;  addr_rom[11886]='h00002438;  wr_data_rom[11886]='h00001cee;
    rd_cycle[11887] = 1'b0;  wr_cycle[11887] = 1'b1;  addr_rom[11887]='h000026b8;  wr_data_rom[11887]='h0000239f;
    rd_cycle[11888] = 1'b1;  wr_cycle[11888] = 1'b0;  addr_rom[11888]='h00001240;  wr_data_rom[11888]='h00000000;
    rd_cycle[11889] = 1'b0;  wr_cycle[11889] = 1'b1;  addr_rom[11889]='h00001e4c;  wr_data_rom[11889]='h000017fe;
    rd_cycle[11890] = 1'b0;  wr_cycle[11890] = 1'b1;  addr_rom[11890]='h00000114;  wr_data_rom[11890]='h00000162;
    rd_cycle[11891] = 1'b0;  wr_cycle[11891] = 1'b1;  addr_rom[11891]='h00003114;  wr_data_rom[11891]='h00001e4f;
    rd_cycle[11892] = 1'b0;  wr_cycle[11892] = 1'b1;  addr_rom[11892]='h00001ca4;  wr_data_rom[11892]='h00003882;
    rd_cycle[11893] = 1'b1;  wr_cycle[11893] = 1'b0;  addr_rom[11893]='h0000271c;  wr_data_rom[11893]='h00000000;
    rd_cycle[11894] = 1'b0;  wr_cycle[11894] = 1'b1;  addr_rom[11894]='h00003244;  wr_data_rom[11894]='h000012f0;
    rd_cycle[11895] = 1'b0;  wr_cycle[11895] = 1'b1;  addr_rom[11895]='h00002f58;  wr_data_rom[11895]='h000022e3;
    rd_cycle[11896] = 1'b0;  wr_cycle[11896] = 1'b1;  addr_rom[11896]='h00002718;  wr_data_rom[11896]='h0000318a;
    rd_cycle[11897] = 1'b0;  wr_cycle[11897] = 1'b1;  addr_rom[11897]='h00000f88;  wr_data_rom[11897]='h00000a2e;
    rd_cycle[11898] = 1'b0;  wr_cycle[11898] = 1'b1;  addr_rom[11898]='h00000494;  wr_data_rom[11898]='h00003dd0;
    rd_cycle[11899] = 1'b0;  wr_cycle[11899] = 1'b1;  addr_rom[11899]='h00002698;  wr_data_rom[11899]='h00001b8f;
    rd_cycle[11900] = 1'b1;  wr_cycle[11900] = 1'b0;  addr_rom[11900]='h00001c6c;  wr_data_rom[11900]='h00000000;
    rd_cycle[11901] = 1'b1;  wr_cycle[11901] = 1'b0;  addr_rom[11901]='h00000278;  wr_data_rom[11901]='h00000000;
    rd_cycle[11902] = 1'b1;  wr_cycle[11902] = 1'b0;  addr_rom[11902]='h00001a78;  wr_data_rom[11902]='h00000000;
    rd_cycle[11903] = 1'b1;  wr_cycle[11903] = 1'b0;  addr_rom[11903]='h000027d8;  wr_data_rom[11903]='h00000000;
    rd_cycle[11904] = 1'b1;  wr_cycle[11904] = 1'b0;  addr_rom[11904]='h00000a2c;  wr_data_rom[11904]='h00000000;
    rd_cycle[11905] = 1'b1;  wr_cycle[11905] = 1'b0;  addr_rom[11905]='h000009fc;  wr_data_rom[11905]='h00000000;
    rd_cycle[11906] = 1'b1;  wr_cycle[11906] = 1'b0;  addr_rom[11906]='h00002888;  wr_data_rom[11906]='h00000000;
    rd_cycle[11907] = 1'b0;  wr_cycle[11907] = 1'b1;  addr_rom[11907]='h000035e8;  wr_data_rom[11907]='h0000195b;
    rd_cycle[11908] = 1'b1;  wr_cycle[11908] = 1'b0;  addr_rom[11908]='h00001698;  wr_data_rom[11908]='h00000000;
    rd_cycle[11909] = 1'b0;  wr_cycle[11909] = 1'b1;  addr_rom[11909]='h0000178c;  wr_data_rom[11909]='h00000878;
    rd_cycle[11910] = 1'b1;  wr_cycle[11910] = 1'b0;  addr_rom[11910]='h0000280c;  wr_data_rom[11910]='h00000000;
    rd_cycle[11911] = 1'b0;  wr_cycle[11911] = 1'b1;  addr_rom[11911]='h00003014;  wr_data_rom[11911]='h00001f7e;
    rd_cycle[11912] = 1'b0;  wr_cycle[11912] = 1'b1;  addr_rom[11912]='h00002ccc;  wr_data_rom[11912]='h00002b9c;
    rd_cycle[11913] = 1'b1;  wr_cycle[11913] = 1'b0;  addr_rom[11913]='h000014dc;  wr_data_rom[11913]='h00000000;
    rd_cycle[11914] = 1'b0;  wr_cycle[11914] = 1'b1;  addr_rom[11914]='h0000026c;  wr_data_rom[11914]='h00002e78;
    rd_cycle[11915] = 1'b0;  wr_cycle[11915] = 1'b1;  addr_rom[11915]='h00002e6c;  wr_data_rom[11915]='h00000420;
    rd_cycle[11916] = 1'b0;  wr_cycle[11916] = 1'b1;  addr_rom[11916]='h00000ca0;  wr_data_rom[11916]='h00000fdd;
    rd_cycle[11917] = 1'b0;  wr_cycle[11917] = 1'b1;  addr_rom[11917]='h00000234;  wr_data_rom[11917]='h0000273b;
    rd_cycle[11918] = 1'b0;  wr_cycle[11918] = 1'b1;  addr_rom[11918]='h0000111c;  wr_data_rom[11918]='h000002e8;
    rd_cycle[11919] = 1'b0;  wr_cycle[11919] = 1'b1;  addr_rom[11919]='h00002ca8;  wr_data_rom[11919]='h00000aa1;
    rd_cycle[11920] = 1'b0;  wr_cycle[11920] = 1'b1;  addr_rom[11920]='h00000be0;  wr_data_rom[11920]='h00003b3c;
    rd_cycle[11921] = 1'b1;  wr_cycle[11921] = 1'b0;  addr_rom[11921]='h0000295c;  wr_data_rom[11921]='h00000000;
    rd_cycle[11922] = 1'b1;  wr_cycle[11922] = 1'b0;  addr_rom[11922]='h00003164;  wr_data_rom[11922]='h00000000;
    rd_cycle[11923] = 1'b1;  wr_cycle[11923] = 1'b0;  addr_rom[11923]='h000035f0;  wr_data_rom[11923]='h00000000;
    rd_cycle[11924] = 1'b0;  wr_cycle[11924] = 1'b1;  addr_rom[11924]='h000031a8;  wr_data_rom[11924]='h00002171;
    rd_cycle[11925] = 1'b1;  wr_cycle[11925] = 1'b0;  addr_rom[11925]='h00001348;  wr_data_rom[11925]='h00000000;
    rd_cycle[11926] = 1'b0;  wr_cycle[11926] = 1'b1;  addr_rom[11926]='h0000341c;  wr_data_rom[11926]='h00002556;
    rd_cycle[11927] = 1'b1;  wr_cycle[11927] = 1'b0;  addr_rom[11927]='h00000dd4;  wr_data_rom[11927]='h00000000;
    rd_cycle[11928] = 1'b1;  wr_cycle[11928] = 1'b0;  addr_rom[11928]='h000038cc;  wr_data_rom[11928]='h00000000;
    rd_cycle[11929] = 1'b1;  wr_cycle[11929] = 1'b0;  addr_rom[11929]='h00003f74;  wr_data_rom[11929]='h00000000;
    rd_cycle[11930] = 1'b1;  wr_cycle[11930] = 1'b0;  addr_rom[11930]='h00003fec;  wr_data_rom[11930]='h00000000;
    rd_cycle[11931] = 1'b0;  wr_cycle[11931] = 1'b1;  addr_rom[11931]='h00001768;  wr_data_rom[11931]='h00002025;
    rd_cycle[11932] = 1'b1;  wr_cycle[11932] = 1'b0;  addr_rom[11932]='h00003398;  wr_data_rom[11932]='h00000000;
    rd_cycle[11933] = 1'b1;  wr_cycle[11933] = 1'b0;  addr_rom[11933]='h00002840;  wr_data_rom[11933]='h00000000;
    rd_cycle[11934] = 1'b1;  wr_cycle[11934] = 1'b0;  addr_rom[11934]='h00002f54;  wr_data_rom[11934]='h00000000;
    rd_cycle[11935] = 1'b0;  wr_cycle[11935] = 1'b1;  addr_rom[11935]='h00000c38;  wr_data_rom[11935]='h000014d9;
    rd_cycle[11936] = 1'b1;  wr_cycle[11936] = 1'b0;  addr_rom[11936]='h00003e9c;  wr_data_rom[11936]='h00000000;
    rd_cycle[11937] = 1'b0;  wr_cycle[11937] = 1'b1;  addr_rom[11937]='h00000cb0;  wr_data_rom[11937]='h00002230;
    rd_cycle[11938] = 1'b0;  wr_cycle[11938] = 1'b1;  addr_rom[11938]='h00003cc0;  wr_data_rom[11938]='h000006b9;
    rd_cycle[11939] = 1'b1;  wr_cycle[11939] = 1'b0;  addr_rom[11939]='h00000ab8;  wr_data_rom[11939]='h00000000;
    rd_cycle[11940] = 1'b0;  wr_cycle[11940] = 1'b1;  addr_rom[11940]='h000029b0;  wr_data_rom[11940]='h00002c60;
    rd_cycle[11941] = 1'b0;  wr_cycle[11941] = 1'b1;  addr_rom[11941]='h00003854;  wr_data_rom[11941]='h00002404;
    rd_cycle[11942] = 1'b1;  wr_cycle[11942] = 1'b0;  addr_rom[11942]='h000034b8;  wr_data_rom[11942]='h00000000;
    rd_cycle[11943] = 1'b0;  wr_cycle[11943] = 1'b1;  addr_rom[11943]='h000021ec;  wr_data_rom[11943]='h00003730;
    rd_cycle[11944] = 1'b1;  wr_cycle[11944] = 1'b0;  addr_rom[11944]='h0000108c;  wr_data_rom[11944]='h00000000;
    rd_cycle[11945] = 1'b1;  wr_cycle[11945] = 1'b0;  addr_rom[11945]='h00002174;  wr_data_rom[11945]='h00000000;
    rd_cycle[11946] = 1'b0;  wr_cycle[11946] = 1'b1;  addr_rom[11946]='h000037dc;  wr_data_rom[11946]='h00003186;
    rd_cycle[11947] = 1'b0;  wr_cycle[11947] = 1'b1;  addr_rom[11947]='h00001a64;  wr_data_rom[11947]='h00003aaa;
    rd_cycle[11948] = 1'b0;  wr_cycle[11948] = 1'b1;  addr_rom[11948]='h00003e78;  wr_data_rom[11948]='h0000376b;
    rd_cycle[11949] = 1'b1;  wr_cycle[11949] = 1'b0;  addr_rom[11949]='h00000b00;  wr_data_rom[11949]='h00000000;
    rd_cycle[11950] = 1'b1;  wr_cycle[11950] = 1'b0;  addr_rom[11950]='h00003fb0;  wr_data_rom[11950]='h00000000;
    rd_cycle[11951] = 1'b0;  wr_cycle[11951] = 1'b1;  addr_rom[11951]='h000008bc;  wr_data_rom[11951]='h0000076f;
    rd_cycle[11952] = 1'b0;  wr_cycle[11952] = 1'b1;  addr_rom[11952]='h00001f2c;  wr_data_rom[11952]='h000006fb;
    rd_cycle[11953] = 1'b0;  wr_cycle[11953] = 1'b1;  addr_rom[11953]='h00003ad8;  wr_data_rom[11953]='h00002c4f;
    rd_cycle[11954] = 1'b1;  wr_cycle[11954] = 1'b0;  addr_rom[11954]='h000023f4;  wr_data_rom[11954]='h00000000;
    rd_cycle[11955] = 1'b1;  wr_cycle[11955] = 1'b0;  addr_rom[11955]='h000026d4;  wr_data_rom[11955]='h00000000;
    rd_cycle[11956] = 1'b1;  wr_cycle[11956] = 1'b0;  addr_rom[11956]='h00002914;  wr_data_rom[11956]='h00000000;
    rd_cycle[11957] = 1'b0;  wr_cycle[11957] = 1'b1;  addr_rom[11957]='h00000e04;  wr_data_rom[11957]='h00000bad;
    rd_cycle[11958] = 1'b1;  wr_cycle[11958] = 1'b0;  addr_rom[11958]='h00002b7c;  wr_data_rom[11958]='h00000000;
    rd_cycle[11959] = 1'b0;  wr_cycle[11959] = 1'b1;  addr_rom[11959]='h00002088;  wr_data_rom[11959]='h00000649;
    rd_cycle[11960] = 1'b1;  wr_cycle[11960] = 1'b0;  addr_rom[11960]='h00000f84;  wr_data_rom[11960]='h00000000;
    rd_cycle[11961] = 1'b1;  wr_cycle[11961] = 1'b0;  addr_rom[11961]='h00002a64;  wr_data_rom[11961]='h00000000;
    rd_cycle[11962] = 1'b1;  wr_cycle[11962] = 1'b0;  addr_rom[11962]='h00002098;  wr_data_rom[11962]='h00000000;
    rd_cycle[11963] = 1'b0;  wr_cycle[11963] = 1'b1;  addr_rom[11963]='h0000175c;  wr_data_rom[11963]='h00003153;
    rd_cycle[11964] = 1'b0;  wr_cycle[11964] = 1'b1;  addr_rom[11964]='h000034a4;  wr_data_rom[11964]='h0000009c;
    rd_cycle[11965] = 1'b0;  wr_cycle[11965] = 1'b1;  addr_rom[11965]='h0000252c;  wr_data_rom[11965]='h00002e7f;
    rd_cycle[11966] = 1'b0;  wr_cycle[11966] = 1'b1;  addr_rom[11966]='h00001cfc;  wr_data_rom[11966]='h00001e82;
    rd_cycle[11967] = 1'b1;  wr_cycle[11967] = 1'b0;  addr_rom[11967]='h00002794;  wr_data_rom[11967]='h00000000;
    rd_cycle[11968] = 1'b0;  wr_cycle[11968] = 1'b1;  addr_rom[11968]='h00003fe0;  wr_data_rom[11968]='h0000070b;
    rd_cycle[11969] = 1'b0;  wr_cycle[11969] = 1'b1;  addr_rom[11969]='h00003604;  wr_data_rom[11969]='h00002b72;
    rd_cycle[11970] = 1'b0;  wr_cycle[11970] = 1'b1;  addr_rom[11970]='h00002280;  wr_data_rom[11970]='h0000249f;
    rd_cycle[11971] = 1'b1;  wr_cycle[11971] = 1'b0;  addr_rom[11971]='h000013b8;  wr_data_rom[11971]='h00000000;
    rd_cycle[11972] = 1'b0;  wr_cycle[11972] = 1'b1;  addr_rom[11972]='h00000a30;  wr_data_rom[11972]='h000029c7;
    rd_cycle[11973] = 1'b1;  wr_cycle[11973] = 1'b0;  addr_rom[11973]='h00001db4;  wr_data_rom[11973]='h00000000;
    rd_cycle[11974] = 1'b1;  wr_cycle[11974] = 1'b0;  addr_rom[11974]='h00000a3c;  wr_data_rom[11974]='h00000000;
    rd_cycle[11975] = 1'b0;  wr_cycle[11975] = 1'b1;  addr_rom[11975]='h00001ca8;  wr_data_rom[11975]='h000036af;
    rd_cycle[11976] = 1'b1;  wr_cycle[11976] = 1'b0;  addr_rom[11976]='h000004b4;  wr_data_rom[11976]='h00000000;
    rd_cycle[11977] = 1'b0;  wr_cycle[11977] = 1'b1;  addr_rom[11977]='h000036e8;  wr_data_rom[11977]='h000001f3;
    rd_cycle[11978] = 1'b1;  wr_cycle[11978] = 1'b0;  addr_rom[11978]='h000015e8;  wr_data_rom[11978]='h00000000;
    rd_cycle[11979] = 1'b1;  wr_cycle[11979] = 1'b0;  addr_rom[11979]='h00001654;  wr_data_rom[11979]='h00000000;
    rd_cycle[11980] = 1'b0;  wr_cycle[11980] = 1'b1;  addr_rom[11980]='h00003f84;  wr_data_rom[11980]='h00001192;
    rd_cycle[11981] = 1'b0;  wr_cycle[11981] = 1'b1;  addr_rom[11981]='h00000e1c;  wr_data_rom[11981]='h00001d71;
    rd_cycle[11982] = 1'b1;  wr_cycle[11982] = 1'b0;  addr_rom[11982]='h00000b30;  wr_data_rom[11982]='h00000000;
    rd_cycle[11983] = 1'b1;  wr_cycle[11983] = 1'b0;  addr_rom[11983]='h00001048;  wr_data_rom[11983]='h00000000;
    rd_cycle[11984] = 1'b1;  wr_cycle[11984] = 1'b0;  addr_rom[11984]='h00003908;  wr_data_rom[11984]='h00000000;
    rd_cycle[11985] = 1'b0;  wr_cycle[11985] = 1'b1;  addr_rom[11985]='h0000182c;  wr_data_rom[11985]='h000021a7;
    rd_cycle[11986] = 1'b0;  wr_cycle[11986] = 1'b1;  addr_rom[11986]='h00003090;  wr_data_rom[11986]='h0000071f;
    rd_cycle[11987] = 1'b1;  wr_cycle[11987] = 1'b0;  addr_rom[11987]='h0000256c;  wr_data_rom[11987]='h00000000;
    rd_cycle[11988] = 1'b0;  wr_cycle[11988] = 1'b1;  addr_rom[11988]='h000031bc;  wr_data_rom[11988]='h00003b1d;
    rd_cycle[11989] = 1'b0;  wr_cycle[11989] = 1'b1;  addr_rom[11989]='h00000964;  wr_data_rom[11989]='h000025ed;
    rd_cycle[11990] = 1'b1;  wr_cycle[11990] = 1'b0;  addr_rom[11990]='h000036a0;  wr_data_rom[11990]='h00000000;
    rd_cycle[11991] = 1'b1;  wr_cycle[11991] = 1'b0;  addr_rom[11991]='h00000cfc;  wr_data_rom[11991]='h00000000;
    rd_cycle[11992] = 1'b1;  wr_cycle[11992] = 1'b0;  addr_rom[11992]='h00001dc0;  wr_data_rom[11992]='h00000000;
    rd_cycle[11993] = 1'b0;  wr_cycle[11993] = 1'b1;  addr_rom[11993]='h00003b1c;  wr_data_rom[11993]='h00000af1;
    rd_cycle[11994] = 1'b0;  wr_cycle[11994] = 1'b1;  addr_rom[11994]='h00001ee4;  wr_data_rom[11994]='h000034c0;
    rd_cycle[11995] = 1'b1;  wr_cycle[11995] = 1'b0;  addr_rom[11995]='h00002100;  wr_data_rom[11995]='h00000000;
    rd_cycle[11996] = 1'b0;  wr_cycle[11996] = 1'b1;  addr_rom[11996]='h00002060;  wr_data_rom[11996]='h0000319c;
    rd_cycle[11997] = 1'b1;  wr_cycle[11997] = 1'b0;  addr_rom[11997]='h000026a0;  wr_data_rom[11997]='h00000000;
    rd_cycle[11998] = 1'b0;  wr_cycle[11998] = 1'b1;  addr_rom[11998]='h0000336c;  wr_data_rom[11998]='h00003990;
    rd_cycle[11999] = 1'b1;  wr_cycle[11999] = 1'b0;  addr_rom[11999]='h00000814;  wr_data_rom[11999]='h00000000;
    rd_cycle[12000] = 1'b0;  wr_cycle[12000] = 1'b1;  addr_rom[12000]='h0000160c;  wr_data_rom[12000]='h00001015;
    rd_cycle[12001] = 1'b1;  wr_cycle[12001] = 1'b0;  addr_rom[12001]='h000011c0;  wr_data_rom[12001]='h00000000;
    rd_cycle[12002] = 1'b0;  wr_cycle[12002] = 1'b1;  addr_rom[12002]='h00003610;  wr_data_rom[12002]='h00002625;
    rd_cycle[12003] = 1'b0;  wr_cycle[12003] = 1'b1;  addr_rom[12003]='h00003a14;  wr_data_rom[12003]='h00001f6a;
    rd_cycle[12004] = 1'b1;  wr_cycle[12004] = 1'b0;  addr_rom[12004]='h00000fe8;  wr_data_rom[12004]='h00000000;
    rd_cycle[12005] = 1'b0;  wr_cycle[12005] = 1'b1;  addr_rom[12005]='h00003f94;  wr_data_rom[12005]='h00000685;
    rd_cycle[12006] = 1'b1;  wr_cycle[12006] = 1'b0;  addr_rom[12006]='h00000338;  wr_data_rom[12006]='h00000000;
    rd_cycle[12007] = 1'b0;  wr_cycle[12007] = 1'b1;  addr_rom[12007]='h00001354;  wr_data_rom[12007]='h00000b0f;
    rd_cycle[12008] = 1'b1;  wr_cycle[12008] = 1'b0;  addr_rom[12008]='h00000a2c;  wr_data_rom[12008]='h00000000;
    rd_cycle[12009] = 1'b1;  wr_cycle[12009] = 1'b0;  addr_rom[12009]='h000019b8;  wr_data_rom[12009]='h00000000;
    rd_cycle[12010] = 1'b1;  wr_cycle[12010] = 1'b0;  addr_rom[12010]='h00000f80;  wr_data_rom[12010]='h00000000;
    rd_cycle[12011] = 1'b1;  wr_cycle[12011] = 1'b0;  addr_rom[12011]='h000023bc;  wr_data_rom[12011]='h00000000;
    rd_cycle[12012] = 1'b0;  wr_cycle[12012] = 1'b1;  addr_rom[12012]='h00002174;  wr_data_rom[12012]='h00002892;
    rd_cycle[12013] = 1'b1;  wr_cycle[12013] = 1'b0;  addr_rom[12013]='h00000340;  wr_data_rom[12013]='h00000000;
    rd_cycle[12014] = 1'b0;  wr_cycle[12014] = 1'b1;  addr_rom[12014]='h000031a0;  wr_data_rom[12014]='h00003271;
    rd_cycle[12015] = 1'b1;  wr_cycle[12015] = 1'b0;  addr_rom[12015]='h00002f2c;  wr_data_rom[12015]='h00000000;
    rd_cycle[12016] = 1'b0;  wr_cycle[12016] = 1'b1;  addr_rom[12016]='h000029a4;  wr_data_rom[12016]='h00001c89;
    rd_cycle[12017] = 1'b1;  wr_cycle[12017] = 1'b0;  addr_rom[12017]='h00002e60;  wr_data_rom[12017]='h00000000;
    rd_cycle[12018] = 1'b1;  wr_cycle[12018] = 1'b0;  addr_rom[12018]='h000030f4;  wr_data_rom[12018]='h00000000;
    rd_cycle[12019] = 1'b0;  wr_cycle[12019] = 1'b1;  addr_rom[12019]='h00002430;  wr_data_rom[12019]='h00003f3a;
    rd_cycle[12020] = 1'b1;  wr_cycle[12020] = 1'b0;  addr_rom[12020]='h00003aec;  wr_data_rom[12020]='h00000000;
    rd_cycle[12021] = 1'b0;  wr_cycle[12021] = 1'b1;  addr_rom[12021]='h00000614;  wr_data_rom[12021]='h00002d4d;
    rd_cycle[12022] = 1'b0;  wr_cycle[12022] = 1'b1;  addr_rom[12022]='h00000b28;  wr_data_rom[12022]='h00000bfa;
    rd_cycle[12023] = 1'b1;  wr_cycle[12023] = 1'b0;  addr_rom[12023]='h00003748;  wr_data_rom[12023]='h00000000;
    rd_cycle[12024] = 1'b1;  wr_cycle[12024] = 1'b0;  addr_rom[12024]='h00003128;  wr_data_rom[12024]='h00000000;
    rd_cycle[12025] = 1'b0;  wr_cycle[12025] = 1'b1;  addr_rom[12025]='h00003ecc;  wr_data_rom[12025]='h00003f0c;
    rd_cycle[12026] = 1'b1;  wr_cycle[12026] = 1'b0;  addr_rom[12026]='h0000194c;  wr_data_rom[12026]='h00000000;
    rd_cycle[12027] = 1'b1;  wr_cycle[12027] = 1'b0;  addr_rom[12027]='h0000197c;  wr_data_rom[12027]='h00000000;
    rd_cycle[12028] = 1'b1;  wr_cycle[12028] = 1'b0;  addr_rom[12028]='h000012e0;  wr_data_rom[12028]='h00000000;
    rd_cycle[12029] = 1'b0;  wr_cycle[12029] = 1'b1;  addr_rom[12029]='h000037fc;  wr_data_rom[12029]='h00001f5d;
    rd_cycle[12030] = 1'b1;  wr_cycle[12030] = 1'b0;  addr_rom[12030]='h00000c5c;  wr_data_rom[12030]='h00000000;
    rd_cycle[12031] = 1'b0;  wr_cycle[12031] = 1'b1;  addr_rom[12031]='h00001b84;  wr_data_rom[12031]='h000019c9;
    rd_cycle[12032] = 1'b1;  wr_cycle[12032] = 1'b0;  addr_rom[12032]='h000035d8;  wr_data_rom[12032]='h00000000;
    rd_cycle[12033] = 1'b0;  wr_cycle[12033] = 1'b1;  addr_rom[12033]='h0000087c;  wr_data_rom[12033]='h00002b28;
    rd_cycle[12034] = 1'b0;  wr_cycle[12034] = 1'b1;  addr_rom[12034]='h00002454;  wr_data_rom[12034]='h0000229c;
    rd_cycle[12035] = 1'b0;  wr_cycle[12035] = 1'b1;  addr_rom[12035]='h000010b8;  wr_data_rom[12035]='h00000003;
    rd_cycle[12036] = 1'b1;  wr_cycle[12036] = 1'b0;  addr_rom[12036]='h000008f4;  wr_data_rom[12036]='h00000000;
    rd_cycle[12037] = 1'b0;  wr_cycle[12037] = 1'b1;  addr_rom[12037]='h000024e0;  wr_data_rom[12037]='h000039fd;
    rd_cycle[12038] = 1'b1;  wr_cycle[12038] = 1'b0;  addr_rom[12038]='h00001894;  wr_data_rom[12038]='h00000000;
    rd_cycle[12039] = 1'b1;  wr_cycle[12039] = 1'b0;  addr_rom[12039]='h00003c18;  wr_data_rom[12039]='h00000000;
    rd_cycle[12040] = 1'b0;  wr_cycle[12040] = 1'b1;  addr_rom[12040]='h00002440;  wr_data_rom[12040]='h000035b5;
    rd_cycle[12041] = 1'b1;  wr_cycle[12041] = 1'b0;  addr_rom[12041]='h00003110;  wr_data_rom[12041]='h00000000;
    rd_cycle[12042] = 1'b0;  wr_cycle[12042] = 1'b1;  addr_rom[12042]='h00002358;  wr_data_rom[12042]='h00003caf;
    rd_cycle[12043] = 1'b0;  wr_cycle[12043] = 1'b1;  addr_rom[12043]='h00003e3c;  wr_data_rom[12043]='h00001dfc;
    rd_cycle[12044] = 1'b0;  wr_cycle[12044] = 1'b1;  addr_rom[12044]='h000026bc;  wr_data_rom[12044]='h000008f9;
    rd_cycle[12045] = 1'b1;  wr_cycle[12045] = 1'b0;  addr_rom[12045]='h0000152c;  wr_data_rom[12045]='h00000000;
    rd_cycle[12046] = 1'b1;  wr_cycle[12046] = 1'b0;  addr_rom[12046]='h00002d3c;  wr_data_rom[12046]='h00000000;
    rd_cycle[12047] = 1'b0;  wr_cycle[12047] = 1'b1;  addr_rom[12047]='h00000cbc;  wr_data_rom[12047]='h00001524;
    rd_cycle[12048] = 1'b1;  wr_cycle[12048] = 1'b0;  addr_rom[12048]='h00003934;  wr_data_rom[12048]='h00000000;
    rd_cycle[12049] = 1'b0;  wr_cycle[12049] = 1'b1;  addr_rom[12049]='h00002884;  wr_data_rom[12049]='h00003a8c;
    rd_cycle[12050] = 1'b1;  wr_cycle[12050] = 1'b0;  addr_rom[12050]='h00002978;  wr_data_rom[12050]='h00000000;
    rd_cycle[12051] = 1'b0;  wr_cycle[12051] = 1'b1;  addr_rom[12051]='h00002770;  wr_data_rom[12051]='h00003928;
    rd_cycle[12052] = 1'b0;  wr_cycle[12052] = 1'b1;  addr_rom[12052]='h00000030;  wr_data_rom[12052]='h00003ddb;
    rd_cycle[12053] = 1'b1;  wr_cycle[12053] = 1'b0;  addr_rom[12053]='h00003238;  wr_data_rom[12053]='h00000000;
    rd_cycle[12054] = 1'b0;  wr_cycle[12054] = 1'b1;  addr_rom[12054]='h000032b4;  wr_data_rom[12054]='h00000ed6;
    rd_cycle[12055] = 1'b0;  wr_cycle[12055] = 1'b1;  addr_rom[12055]='h00003944;  wr_data_rom[12055]='h00001c38;
    rd_cycle[12056] = 1'b1;  wr_cycle[12056] = 1'b0;  addr_rom[12056]='h000006a4;  wr_data_rom[12056]='h00000000;
    rd_cycle[12057] = 1'b1;  wr_cycle[12057] = 1'b0;  addr_rom[12057]='h00000ff4;  wr_data_rom[12057]='h00000000;
    rd_cycle[12058] = 1'b1;  wr_cycle[12058] = 1'b0;  addr_rom[12058]='h00001910;  wr_data_rom[12058]='h00000000;
    rd_cycle[12059] = 1'b0;  wr_cycle[12059] = 1'b1;  addr_rom[12059]='h00003b3c;  wr_data_rom[12059]='h0000182f;
    rd_cycle[12060] = 1'b0;  wr_cycle[12060] = 1'b1;  addr_rom[12060]='h000031bc;  wr_data_rom[12060]='h000021e3;
    rd_cycle[12061] = 1'b1;  wr_cycle[12061] = 1'b0;  addr_rom[12061]='h000022ec;  wr_data_rom[12061]='h00000000;
    rd_cycle[12062] = 1'b0;  wr_cycle[12062] = 1'b1;  addr_rom[12062]='h00001154;  wr_data_rom[12062]='h00003845;
    rd_cycle[12063] = 1'b0;  wr_cycle[12063] = 1'b1;  addr_rom[12063]='h000023d8;  wr_data_rom[12063]='h00002dab;
    rd_cycle[12064] = 1'b0;  wr_cycle[12064] = 1'b1;  addr_rom[12064]='h00000ca0;  wr_data_rom[12064]='h000037ff;
    rd_cycle[12065] = 1'b0;  wr_cycle[12065] = 1'b1;  addr_rom[12065]='h00000248;  wr_data_rom[12065]='h00003691;
    rd_cycle[12066] = 1'b1;  wr_cycle[12066] = 1'b0;  addr_rom[12066]='h00002a5c;  wr_data_rom[12066]='h00000000;
    rd_cycle[12067] = 1'b0;  wr_cycle[12067] = 1'b1;  addr_rom[12067]='h00001748;  wr_data_rom[12067]='h00003fb3;
    rd_cycle[12068] = 1'b1;  wr_cycle[12068] = 1'b0;  addr_rom[12068]='h00000cd4;  wr_data_rom[12068]='h00000000;
    rd_cycle[12069] = 1'b1;  wr_cycle[12069] = 1'b0;  addr_rom[12069]='h00001fbc;  wr_data_rom[12069]='h00000000;
    rd_cycle[12070] = 1'b1;  wr_cycle[12070] = 1'b0;  addr_rom[12070]='h00002100;  wr_data_rom[12070]='h00000000;
    rd_cycle[12071] = 1'b1;  wr_cycle[12071] = 1'b0;  addr_rom[12071]='h000004c0;  wr_data_rom[12071]='h00000000;
    rd_cycle[12072] = 1'b0;  wr_cycle[12072] = 1'b1;  addr_rom[12072]='h0000384c;  wr_data_rom[12072]='h00000706;
    rd_cycle[12073] = 1'b0;  wr_cycle[12073] = 1'b1;  addr_rom[12073]='h000036e0;  wr_data_rom[12073]='h00000c12;
    rd_cycle[12074] = 1'b0;  wr_cycle[12074] = 1'b1;  addr_rom[12074]='h000009ec;  wr_data_rom[12074]='h00003473;
    rd_cycle[12075] = 1'b1;  wr_cycle[12075] = 1'b0;  addr_rom[12075]='h0000077c;  wr_data_rom[12075]='h00000000;
    rd_cycle[12076] = 1'b0;  wr_cycle[12076] = 1'b1;  addr_rom[12076]='h00001dc0;  wr_data_rom[12076]='h00003ba6;
    rd_cycle[12077] = 1'b0;  wr_cycle[12077] = 1'b1;  addr_rom[12077]='h000006e0;  wr_data_rom[12077]='h0000022b;
    rd_cycle[12078] = 1'b0;  wr_cycle[12078] = 1'b1;  addr_rom[12078]='h00000bfc;  wr_data_rom[12078]='h00000c0d;
    rd_cycle[12079] = 1'b1;  wr_cycle[12079] = 1'b0;  addr_rom[12079]='h00003210;  wr_data_rom[12079]='h00000000;
    rd_cycle[12080] = 1'b1;  wr_cycle[12080] = 1'b0;  addr_rom[12080]='h00003180;  wr_data_rom[12080]='h00000000;
    rd_cycle[12081] = 1'b0;  wr_cycle[12081] = 1'b1;  addr_rom[12081]='h00001474;  wr_data_rom[12081]='h0000379f;
    rd_cycle[12082] = 1'b1;  wr_cycle[12082] = 1'b0;  addr_rom[12082]='h000010f4;  wr_data_rom[12082]='h00000000;
    rd_cycle[12083] = 1'b1;  wr_cycle[12083] = 1'b0;  addr_rom[12083]='h000018b0;  wr_data_rom[12083]='h00000000;
    rd_cycle[12084] = 1'b1;  wr_cycle[12084] = 1'b0;  addr_rom[12084]='h00002304;  wr_data_rom[12084]='h00000000;
    rd_cycle[12085] = 1'b0;  wr_cycle[12085] = 1'b1;  addr_rom[12085]='h0000296c;  wr_data_rom[12085]='h00001a87;
    rd_cycle[12086] = 1'b1;  wr_cycle[12086] = 1'b0;  addr_rom[12086]='h00001b74;  wr_data_rom[12086]='h00000000;
    rd_cycle[12087] = 1'b0;  wr_cycle[12087] = 1'b1;  addr_rom[12087]='h00003334;  wr_data_rom[12087]='h000026b1;
    rd_cycle[12088] = 1'b0;  wr_cycle[12088] = 1'b1;  addr_rom[12088]='h00000c50;  wr_data_rom[12088]='h00003af7;
    rd_cycle[12089] = 1'b1;  wr_cycle[12089] = 1'b0;  addr_rom[12089]='h00003f7c;  wr_data_rom[12089]='h00000000;
    rd_cycle[12090] = 1'b0;  wr_cycle[12090] = 1'b1;  addr_rom[12090]='h00003940;  wr_data_rom[12090]='h00000358;
    rd_cycle[12091] = 1'b1;  wr_cycle[12091] = 1'b0;  addr_rom[12091]='h000029b4;  wr_data_rom[12091]='h00000000;
    rd_cycle[12092] = 1'b1;  wr_cycle[12092] = 1'b0;  addr_rom[12092]='h00002494;  wr_data_rom[12092]='h00000000;
    rd_cycle[12093] = 1'b0;  wr_cycle[12093] = 1'b1;  addr_rom[12093]='h00000b94;  wr_data_rom[12093]='h000024ff;
    rd_cycle[12094] = 1'b0;  wr_cycle[12094] = 1'b1;  addr_rom[12094]='h00001d98;  wr_data_rom[12094]='h00000932;
    rd_cycle[12095] = 1'b0;  wr_cycle[12095] = 1'b1;  addr_rom[12095]='h00003d6c;  wr_data_rom[12095]='h00002126;
    rd_cycle[12096] = 1'b0;  wr_cycle[12096] = 1'b1;  addr_rom[12096]='h00002230;  wr_data_rom[12096]='h000039b9;
    rd_cycle[12097] = 1'b0;  wr_cycle[12097] = 1'b1;  addr_rom[12097]='h00000ad4;  wr_data_rom[12097]='h000025c2;
    rd_cycle[12098] = 1'b0;  wr_cycle[12098] = 1'b1;  addr_rom[12098]='h0000210c;  wr_data_rom[12098]='h00002b05;
    rd_cycle[12099] = 1'b1;  wr_cycle[12099] = 1'b0;  addr_rom[12099]='h00000658;  wr_data_rom[12099]='h00000000;
    rd_cycle[12100] = 1'b0;  wr_cycle[12100] = 1'b1;  addr_rom[12100]='h00003774;  wr_data_rom[12100]='h0000227f;
    rd_cycle[12101] = 1'b1;  wr_cycle[12101] = 1'b0;  addr_rom[12101]='h00000c80;  wr_data_rom[12101]='h00000000;
    rd_cycle[12102] = 1'b0;  wr_cycle[12102] = 1'b1;  addr_rom[12102]='h00002ab8;  wr_data_rom[12102]='h00000aa3;
    rd_cycle[12103] = 1'b1;  wr_cycle[12103] = 1'b0;  addr_rom[12103]='h00001c7c;  wr_data_rom[12103]='h00000000;
    rd_cycle[12104] = 1'b0;  wr_cycle[12104] = 1'b1;  addr_rom[12104]='h000031ac;  wr_data_rom[12104]='h000038f3;
    rd_cycle[12105] = 1'b1;  wr_cycle[12105] = 1'b0;  addr_rom[12105]='h000031f4;  wr_data_rom[12105]='h00000000;
    rd_cycle[12106] = 1'b1;  wr_cycle[12106] = 1'b0;  addr_rom[12106]='h00002f84;  wr_data_rom[12106]='h00000000;
    rd_cycle[12107] = 1'b0;  wr_cycle[12107] = 1'b1;  addr_rom[12107]='h00002b9c;  wr_data_rom[12107]='h00000264;
    rd_cycle[12108] = 1'b1;  wr_cycle[12108] = 1'b0;  addr_rom[12108]='h00000fa0;  wr_data_rom[12108]='h00000000;
    rd_cycle[12109] = 1'b1;  wr_cycle[12109] = 1'b0;  addr_rom[12109]='h00002234;  wr_data_rom[12109]='h00000000;
    rd_cycle[12110] = 1'b0;  wr_cycle[12110] = 1'b1;  addr_rom[12110]='h00003f10;  wr_data_rom[12110]='h00003ef7;
    rd_cycle[12111] = 1'b1;  wr_cycle[12111] = 1'b0;  addr_rom[12111]='h00002cec;  wr_data_rom[12111]='h00000000;
    rd_cycle[12112] = 1'b1;  wr_cycle[12112] = 1'b0;  addr_rom[12112]='h00001ee4;  wr_data_rom[12112]='h00000000;
    rd_cycle[12113] = 1'b0;  wr_cycle[12113] = 1'b1;  addr_rom[12113]='h000034b8;  wr_data_rom[12113]='h00002850;
    rd_cycle[12114] = 1'b1;  wr_cycle[12114] = 1'b0;  addr_rom[12114]='h00003d94;  wr_data_rom[12114]='h00000000;
    rd_cycle[12115] = 1'b0;  wr_cycle[12115] = 1'b1;  addr_rom[12115]='h00002ff0;  wr_data_rom[12115]='h000000d9;
    rd_cycle[12116] = 1'b1;  wr_cycle[12116] = 1'b0;  addr_rom[12116]='h00002cb0;  wr_data_rom[12116]='h00000000;
    rd_cycle[12117] = 1'b0;  wr_cycle[12117] = 1'b1;  addr_rom[12117]='h000005b8;  wr_data_rom[12117]='h00002581;
    rd_cycle[12118] = 1'b1;  wr_cycle[12118] = 1'b0;  addr_rom[12118]='h000037c0;  wr_data_rom[12118]='h00000000;
    rd_cycle[12119] = 1'b1;  wr_cycle[12119] = 1'b0;  addr_rom[12119]='h000025dc;  wr_data_rom[12119]='h00000000;
    rd_cycle[12120] = 1'b0;  wr_cycle[12120] = 1'b1;  addr_rom[12120]='h000035dc;  wr_data_rom[12120]='h000030d2;
    rd_cycle[12121] = 1'b0;  wr_cycle[12121] = 1'b1;  addr_rom[12121]='h00003230;  wr_data_rom[12121]='h00003bd7;
    rd_cycle[12122] = 1'b1;  wr_cycle[12122] = 1'b0;  addr_rom[12122]='h00003e14;  wr_data_rom[12122]='h00000000;
    rd_cycle[12123] = 1'b1;  wr_cycle[12123] = 1'b0;  addr_rom[12123]='h00003a14;  wr_data_rom[12123]='h00000000;
    rd_cycle[12124] = 1'b1;  wr_cycle[12124] = 1'b0;  addr_rom[12124]='h000033a8;  wr_data_rom[12124]='h00000000;
    rd_cycle[12125] = 1'b0;  wr_cycle[12125] = 1'b1;  addr_rom[12125]='h00002e50;  wr_data_rom[12125]='h00003f88;
    rd_cycle[12126] = 1'b1;  wr_cycle[12126] = 1'b0;  addr_rom[12126]='h00002518;  wr_data_rom[12126]='h00000000;
    rd_cycle[12127] = 1'b1;  wr_cycle[12127] = 1'b0;  addr_rom[12127]='h00003a90;  wr_data_rom[12127]='h00000000;
    rd_cycle[12128] = 1'b0;  wr_cycle[12128] = 1'b1;  addr_rom[12128]='h00003064;  wr_data_rom[12128]='h000028cc;
    rd_cycle[12129] = 1'b0;  wr_cycle[12129] = 1'b1;  addr_rom[12129]='h000018f0;  wr_data_rom[12129]='h00000523;
    rd_cycle[12130] = 1'b0;  wr_cycle[12130] = 1'b1;  addr_rom[12130]='h000026a4;  wr_data_rom[12130]='h00003096;
    rd_cycle[12131] = 1'b0;  wr_cycle[12131] = 1'b1;  addr_rom[12131]='h00000720;  wr_data_rom[12131]='h00002a1d;
    rd_cycle[12132] = 1'b1;  wr_cycle[12132] = 1'b0;  addr_rom[12132]='h00002454;  wr_data_rom[12132]='h00000000;
    rd_cycle[12133] = 1'b0;  wr_cycle[12133] = 1'b1;  addr_rom[12133]='h00003810;  wr_data_rom[12133]='h0000043b;
    rd_cycle[12134] = 1'b1;  wr_cycle[12134] = 1'b0;  addr_rom[12134]='h00001fac;  wr_data_rom[12134]='h00000000;
    rd_cycle[12135] = 1'b0;  wr_cycle[12135] = 1'b1;  addr_rom[12135]='h00003744;  wr_data_rom[12135]='h0000395b;
    rd_cycle[12136] = 1'b0;  wr_cycle[12136] = 1'b1;  addr_rom[12136]='h00001b58;  wr_data_rom[12136]='h00003ab2;
    rd_cycle[12137] = 1'b0;  wr_cycle[12137] = 1'b1;  addr_rom[12137]='h000000d4;  wr_data_rom[12137]='h00001eca;
    rd_cycle[12138] = 1'b1;  wr_cycle[12138] = 1'b0;  addr_rom[12138]='h00002680;  wr_data_rom[12138]='h00000000;
    rd_cycle[12139] = 1'b1;  wr_cycle[12139] = 1'b0;  addr_rom[12139]='h0000141c;  wr_data_rom[12139]='h00000000;
    rd_cycle[12140] = 1'b1;  wr_cycle[12140] = 1'b0;  addr_rom[12140]='h00001e54;  wr_data_rom[12140]='h00000000;
    rd_cycle[12141] = 1'b1;  wr_cycle[12141] = 1'b0;  addr_rom[12141]='h00003020;  wr_data_rom[12141]='h00000000;
    rd_cycle[12142] = 1'b0;  wr_cycle[12142] = 1'b1;  addr_rom[12142]='h00001028;  wr_data_rom[12142]='h00000c19;
    rd_cycle[12143] = 1'b1;  wr_cycle[12143] = 1'b0;  addr_rom[12143]='h00002014;  wr_data_rom[12143]='h00000000;
    rd_cycle[12144] = 1'b0;  wr_cycle[12144] = 1'b1;  addr_rom[12144]='h00003ca0;  wr_data_rom[12144]='h00003316;
    rd_cycle[12145] = 1'b1;  wr_cycle[12145] = 1'b0;  addr_rom[12145]='h00002dc8;  wr_data_rom[12145]='h00000000;
    rd_cycle[12146] = 1'b0;  wr_cycle[12146] = 1'b1;  addr_rom[12146]='h00001b90;  wr_data_rom[12146]='h000004b2;
    rd_cycle[12147] = 1'b1;  wr_cycle[12147] = 1'b0;  addr_rom[12147]='h00003714;  wr_data_rom[12147]='h00000000;
    rd_cycle[12148] = 1'b0;  wr_cycle[12148] = 1'b1;  addr_rom[12148]='h00000030;  wr_data_rom[12148]='h00003ab3;
    rd_cycle[12149] = 1'b1;  wr_cycle[12149] = 1'b0;  addr_rom[12149]='h000012fc;  wr_data_rom[12149]='h00000000;
    rd_cycle[12150] = 1'b0;  wr_cycle[12150] = 1'b1;  addr_rom[12150]='h00003a9c;  wr_data_rom[12150]='h00001a06;
    rd_cycle[12151] = 1'b1;  wr_cycle[12151] = 1'b0;  addr_rom[12151]='h000007e0;  wr_data_rom[12151]='h00000000;
    rd_cycle[12152] = 1'b1;  wr_cycle[12152] = 1'b0;  addr_rom[12152]='h00000b30;  wr_data_rom[12152]='h00000000;
    rd_cycle[12153] = 1'b1;  wr_cycle[12153] = 1'b0;  addr_rom[12153]='h00000a04;  wr_data_rom[12153]='h00000000;
    rd_cycle[12154] = 1'b1;  wr_cycle[12154] = 1'b0;  addr_rom[12154]='h00002a30;  wr_data_rom[12154]='h00000000;
    rd_cycle[12155] = 1'b1;  wr_cycle[12155] = 1'b0;  addr_rom[12155]='h00000640;  wr_data_rom[12155]='h00000000;
    rd_cycle[12156] = 1'b1;  wr_cycle[12156] = 1'b0;  addr_rom[12156]='h00002074;  wr_data_rom[12156]='h00000000;
    rd_cycle[12157] = 1'b0;  wr_cycle[12157] = 1'b1;  addr_rom[12157]='h00002dd0;  wr_data_rom[12157]='h00002b35;
    rd_cycle[12158] = 1'b1;  wr_cycle[12158] = 1'b0;  addr_rom[12158]='h00000c40;  wr_data_rom[12158]='h00000000;
    rd_cycle[12159] = 1'b1;  wr_cycle[12159] = 1'b0;  addr_rom[12159]='h00002844;  wr_data_rom[12159]='h00000000;
    rd_cycle[12160] = 1'b1;  wr_cycle[12160] = 1'b0;  addr_rom[12160]='h00000454;  wr_data_rom[12160]='h00000000;
    rd_cycle[12161] = 1'b0;  wr_cycle[12161] = 1'b1;  addr_rom[12161]='h00002344;  wr_data_rom[12161]='h0000381b;
    rd_cycle[12162] = 1'b1;  wr_cycle[12162] = 1'b0;  addr_rom[12162]='h00000948;  wr_data_rom[12162]='h00000000;
    rd_cycle[12163] = 1'b0;  wr_cycle[12163] = 1'b1;  addr_rom[12163]='h0000101c;  wr_data_rom[12163]='h0000202f;
    rd_cycle[12164] = 1'b1;  wr_cycle[12164] = 1'b0;  addr_rom[12164]='h000006d4;  wr_data_rom[12164]='h00000000;
    rd_cycle[12165] = 1'b0;  wr_cycle[12165] = 1'b1;  addr_rom[12165]='h000036fc;  wr_data_rom[12165]='h000023df;
    rd_cycle[12166] = 1'b1;  wr_cycle[12166] = 1'b0;  addr_rom[12166]='h00003544;  wr_data_rom[12166]='h00000000;
    rd_cycle[12167] = 1'b1;  wr_cycle[12167] = 1'b0;  addr_rom[12167]='h00003b84;  wr_data_rom[12167]='h00000000;
    rd_cycle[12168] = 1'b1;  wr_cycle[12168] = 1'b0;  addr_rom[12168]='h00002110;  wr_data_rom[12168]='h00000000;
    rd_cycle[12169] = 1'b0;  wr_cycle[12169] = 1'b1;  addr_rom[12169]='h00000cd0;  wr_data_rom[12169]='h00003677;
    rd_cycle[12170] = 1'b1;  wr_cycle[12170] = 1'b0;  addr_rom[12170]='h00002aa4;  wr_data_rom[12170]='h00000000;
    rd_cycle[12171] = 1'b1;  wr_cycle[12171] = 1'b0;  addr_rom[12171]='h00002a4c;  wr_data_rom[12171]='h00000000;
    rd_cycle[12172] = 1'b1;  wr_cycle[12172] = 1'b0;  addr_rom[12172]='h00003160;  wr_data_rom[12172]='h00000000;
    rd_cycle[12173] = 1'b1;  wr_cycle[12173] = 1'b0;  addr_rom[12173]='h00003538;  wr_data_rom[12173]='h00000000;
    rd_cycle[12174] = 1'b1;  wr_cycle[12174] = 1'b0;  addr_rom[12174]='h000033bc;  wr_data_rom[12174]='h00000000;
    rd_cycle[12175] = 1'b0;  wr_cycle[12175] = 1'b1;  addr_rom[12175]='h00002cc0;  wr_data_rom[12175]='h000025fe;
    rd_cycle[12176] = 1'b1;  wr_cycle[12176] = 1'b0;  addr_rom[12176]='h0000264c;  wr_data_rom[12176]='h00000000;
    rd_cycle[12177] = 1'b1;  wr_cycle[12177] = 1'b0;  addr_rom[12177]='h00003000;  wr_data_rom[12177]='h00000000;
    rd_cycle[12178] = 1'b1;  wr_cycle[12178] = 1'b0;  addr_rom[12178]='h0000080c;  wr_data_rom[12178]='h00000000;
    rd_cycle[12179] = 1'b1;  wr_cycle[12179] = 1'b0;  addr_rom[12179]='h000023f8;  wr_data_rom[12179]='h00000000;
    rd_cycle[12180] = 1'b1;  wr_cycle[12180] = 1'b0;  addr_rom[12180]='h0000299c;  wr_data_rom[12180]='h00000000;
    rd_cycle[12181] = 1'b1;  wr_cycle[12181] = 1'b0;  addr_rom[12181]='h000015dc;  wr_data_rom[12181]='h00000000;
    rd_cycle[12182] = 1'b1;  wr_cycle[12182] = 1'b0;  addr_rom[12182]='h000030a4;  wr_data_rom[12182]='h00000000;
    rd_cycle[12183] = 1'b1;  wr_cycle[12183] = 1'b0;  addr_rom[12183]='h00002454;  wr_data_rom[12183]='h00000000;
    rd_cycle[12184] = 1'b0;  wr_cycle[12184] = 1'b1;  addr_rom[12184]='h00002a1c;  wr_data_rom[12184]='h00000d65;
    rd_cycle[12185] = 1'b1;  wr_cycle[12185] = 1'b0;  addr_rom[12185]='h00002834;  wr_data_rom[12185]='h00000000;
    rd_cycle[12186] = 1'b0;  wr_cycle[12186] = 1'b1;  addr_rom[12186]='h00003ed8;  wr_data_rom[12186]='h000029b7;
    rd_cycle[12187] = 1'b0;  wr_cycle[12187] = 1'b1;  addr_rom[12187]='h000014e8;  wr_data_rom[12187]='h000003ae;
    rd_cycle[12188] = 1'b0;  wr_cycle[12188] = 1'b1;  addr_rom[12188]='h00002198;  wr_data_rom[12188]='h000013e7;
    rd_cycle[12189] = 1'b1;  wr_cycle[12189] = 1'b0;  addr_rom[12189]='h00000ebc;  wr_data_rom[12189]='h00000000;
    rd_cycle[12190] = 1'b1;  wr_cycle[12190] = 1'b0;  addr_rom[12190]='h00000f40;  wr_data_rom[12190]='h00000000;
    rd_cycle[12191] = 1'b0;  wr_cycle[12191] = 1'b1;  addr_rom[12191]='h00000a5c;  wr_data_rom[12191]='h000037c7;
    rd_cycle[12192] = 1'b1;  wr_cycle[12192] = 1'b0;  addr_rom[12192]='h00001f80;  wr_data_rom[12192]='h00000000;
    rd_cycle[12193] = 1'b1;  wr_cycle[12193] = 1'b0;  addr_rom[12193]='h00002008;  wr_data_rom[12193]='h00000000;
    rd_cycle[12194] = 1'b0;  wr_cycle[12194] = 1'b1;  addr_rom[12194]='h00003cbc;  wr_data_rom[12194]='h00000a25;
    rd_cycle[12195] = 1'b1;  wr_cycle[12195] = 1'b0;  addr_rom[12195]='h0000263c;  wr_data_rom[12195]='h00000000;
    rd_cycle[12196] = 1'b1;  wr_cycle[12196] = 1'b0;  addr_rom[12196]='h00000ce4;  wr_data_rom[12196]='h00000000;
    rd_cycle[12197] = 1'b0;  wr_cycle[12197] = 1'b1;  addr_rom[12197]='h00003238;  wr_data_rom[12197]='h000027b2;
    rd_cycle[12198] = 1'b1;  wr_cycle[12198] = 1'b0;  addr_rom[12198]='h00000c4c;  wr_data_rom[12198]='h00000000;
    rd_cycle[12199] = 1'b0;  wr_cycle[12199] = 1'b1;  addr_rom[12199]='h00003848;  wr_data_rom[12199]='h0000025d;
    rd_cycle[12200] = 1'b0;  wr_cycle[12200] = 1'b1;  addr_rom[12200]='h000003a0;  wr_data_rom[12200]='h00002b86;
    rd_cycle[12201] = 1'b1;  wr_cycle[12201] = 1'b0;  addr_rom[12201]='h000017c8;  wr_data_rom[12201]='h00000000;
    rd_cycle[12202] = 1'b1;  wr_cycle[12202] = 1'b0;  addr_rom[12202]='h00002344;  wr_data_rom[12202]='h00000000;
    rd_cycle[12203] = 1'b0;  wr_cycle[12203] = 1'b1;  addr_rom[12203]='h000032fc;  wr_data_rom[12203]='h00001fe7;
    rd_cycle[12204] = 1'b1;  wr_cycle[12204] = 1'b0;  addr_rom[12204]='h000011f0;  wr_data_rom[12204]='h00000000;
    rd_cycle[12205] = 1'b1;  wr_cycle[12205] = 1'b0;  addr_rom[12205]='h00003fac;  wr_data_rom[12205]='h00000000;
    rd_cycle[12206] = 1'b1;  wr_cycle[12206] = 1'b0;  addr_rom[12206]='h00001264;  wr_data_rom[12206]='h00000000;
    rd_cycle[12207] = 1'b1;  wr_cycle[12207] = 1'b0;  addr_rom[12207]='h00000f64;  wr_data_rom[12207]='h00000000;
    rd_cycle[12208] = 1'b1;  wr_cycle[12208] = 1'b0;  addr_rom[12208]='h000037e8;  wr_data_rom[12208]='h00000000;
    rd_cycle[12209] = 1'b0;  wr_cycle[12209] = 1'b1;  addr_rom[12209]='h000037f8;  wr_data_rom[12209]='h0000102c;
    rd_cycle[12210] = 1'b0;  wr_cycle[12210] = 1'b1;  addr_rom[12210]='h000018fc;  wr_data_rom[12210]='h00000d34;
    rd_cycle[12211] = 1'b1;  wr_cycle[12211] = 1'b0;  addr_rom[12211]='h000037c0;  wr_data_rom[12211]='h00000000;
    rd_cycle[12212] = 1'b1;  wr_cycle[12212] = 1'b0;  addr_rom[12212]='h00003dac;  wr_data_rom[12212]='h00000000;
    rd_cycle[12213] = 1'b0;  wr_cycle[12213] = 1'b1;  addr_rom[12213]='h00002ee8;  wr_data_rom[12213]='h00002b0a;
    rd_cycle[12214] = 1'b0;  wr_cycle[12214] = 1'b1;  addr_rom[12214]='h0000385c;  wr_data_rom[12214]='h0000206c;
    rd_cycle[12215] = 1'b1;  wr_cycle[12215] = 1'b0;  addr_rom[12215]='h00000304;  wr_data_rom[12215]='h00000000;
    rd_cycle[12216] = 1'b1;  wr_cycle[12216] = 1'b0;  addr_rom[12216]='h000012c8;  wr_data_rom[12216]='h00000000;
    rd_cycle[12217] = 1'b1;  wr_cycle[12217] = 1'b0;  addr_rom[12217]='h000013c0;  wr_data_rom[12217]='h00000000;
    rd_cycle[12218] = 1'b1;  wr_cycle[12218] = 1'b0;  addr_rom[12218]='h000016bc;  wr_data_rom[12218]='h00000000;
    rd_cycle[12219] = 1'b1;  wr_cycle[12219] = 1'b0;  addr_rom[12219]='h0000123c;  wr_data_rom[12219]='h00000000;
    rd_cycle[12220] = 1'b1;  wr_cycle[12220] = 1'b0;  addr_rom[12220]='h00002c6c;  wr_data_rom[12220]='h00000000;
    rd_cycle[12221] = 1'b0;  wr_cycle[12221] = 1'b1;  addr_rom[12221]='h00000018;  wr_data_rom[12221]='h00003a24;
    rd_cycle[12222] = 1'b0;  wr_cycle[12222] = 1'b1;  addr_rom[12222]='h00003f48;  wr_data_rom[12222]='h000027fe;
    rd_cycle[12223] = 1'b0;  wr_cycle[12223] = 1'b1;  addr_rom[12223]='h00003edc;  wr_data_rom[12223]='h00003008;
    rd_cycle[12224] = 1'b0;  wr_cycle[12224] = 1'b1;  addr_rom[12224]='h0000293c;  wr_data_rom[12224]='h00000a3e;
    rd_cycle[12225] = 1'b1;  wr_cycle[12225] = 1'b0;  addr_rom[12225]='h000021a0;  wr_data_rom[12225]='h00000000;
    rd_cycle[12226] = 1'b1;  wr_cycle[12226] = 1'b0;  addr_rom[12226]='h0000329c;  wr_data_rom[12226]='h00000000;
    rd_cycle[12227] = 1'b1;  wr_cycle[12227] = 1'b0;  addr_rom[12227]='h00003dfc;  wr_data_rom[12227]='h00000000;
    rd_cycle[12228] = 1'b1;  wr_cycle[12228] = 1'b0;  addr_rom[12228]='h000029d8;  wr_data_rom[12228]='h00000000;
    rd_cycle[12229] = 1'b0;  wr_cycle[12229] = 1'b1;  addr_rom[12229]='h00001374;  wr_data_rom[12229]='h00002ac4;
    rd_cycle[12230] = 1'b1;  wr_cycle[12230] = 1'b0;  addr_rom[12230]='h00003b38;  wr_data_rom[12230]='h00000000;
    rd_cycle[12231] = 1'b1;  wr_cycle[12231] = 1'b0;  addr_rom[12231]='h000026b0;  wr_data_rom[12231]='h00000000;
    rd_cycle[12232] = 1'b0;  wr_cycle[12232] = 1'b1;  addr_rom[12232]='h00000d74;  wr_data_rom[12232]='h00002862;
    rd_cycle[12233] = 1'b1;  wr_cycle[12233] = 1'b0;  addr_rom[12233]='h000039d8;  wr_data_rom[12233]='h00000000;
    rd_cycle[12234] = 1'b0;  wr_cycle[12234] = 1'b1;  addr_rom[12234]='h000014d8;  wr_data_rom[12234]='h0000034d;
    rd_cycle[12235] = 1'b1;  wr_cycle[12235] = 1'b0;  addr_rom[12235]='h0000030c;  wr_data_rom[12235]='h00000000;
    rd_cycle[12236] = 1'b1;  wr_cycle[12236] = 1'b0;  addr_rom[12236]='h00000100;  wr_data_rom[12236]='h00000000;
    rd_cycle[12237] = 1'b0;  wr_cycle[12237] = 1'b1;  addr_rom[12237]='h000024f4;  wr_data_rom[12237]='h00000163;
    rd_cycle[12238] = 1'b1;  wr_cycle[12238] = 1'b0;  addr_rom[12238]='h000008d0;  wr_data_rom[12238]='h00000000;
    rd_cycle[12239] = 1'b0;  wr_cycle[12239] = 1'b1;  addr_rom[12239]='h00002744;  wr_data_rom[12239]='h00000ce7;
    rd_cycle[12240] = 1'b0;  wr_cycle[12240] = 1'b1;  addr_rom[12240]='h00000d44;  wr_data_rom[12240]='h0000248d;
    rd_cycle[12241] = 1'b1;  wr_cycle[12241] = 1'b0;  addr_rom[12241]='h00003b08;  wr_data_rom[12241]='h00000000;
    rd_cycle[12242] = 1'b1;  wr_cycle[12242] = 1'b0;  addr_rom[12242]='h00003dcc;  wr_data_rom[12242]='h00000000;
    rd_cycle[12243] = 1'b0;  wr_cycle[12243] = 1'b1;  addr_rom[12243]='h000016ec;  wr_data_rom[12243]='h00002e65;
    rd_cycle[12244] = 1'b0;  wr_cycle[12244] = 1'b1;  addr_rom[12244]='h00003264;  wr_data_rom[12244]='h000003f7;
    rd_cycle[12245] = 1'b0;  wr_cycle[12245] = 1'b1;  addr_rom[12245]='h000016c0;  wr_data_rom[12245]='h0000374e;
    rd_cycle[12246] = 1'b1;  wr_cycle[12246] = 1'b0;  addr_rom[12246]='h00000a8c;  wr_data_rom[12246]='h00000000;
    rd_cycle[12247] = 1'b0;  wr_cycle[12247] = 1'b1;  addr_rom[12247]='h00000e0c;  wr_data_rom[12247]='h00002aa8;
    rd_cycle[12248] = 1'b1;  wr_cycle[12248] = 1'b0;  addr_rom[12248]='h00002580;  wr_data_rom[12248]='h00000000;
    rd_cycle[12249] = 1'b0;  wr_cycle[12249] = 1'b1;  addr_rom[12249]='h0000381c;  wr_data_rom[12249]='h000005ec;
    rd_cycle[12250] = 1'b1;  wr_cycle[12250] = 1'b0;  addr_rom[12250]='h00001708;  wr_data_rom[12250]='h00000000;
    rd_cycle[12251] = 1'b0;  wr_cycle[12251] = 1'b1;  addr_rom[12251]='h000016e4;  wr_data_rom[12251]='h000011c6;
    rd_cycle[12252] = 1'b0;  wr_cycle[12252] = 1'b1;  addr_rom[12252]='h000037d0;  wr_data_rom[12252]='h00002d5d;
    rd_cycle[12253] = 1'b1;  wr_cycle[12253] = 1'b0;  addr_rom[12253]='h00000d44;  wr_data_rom[12253]='h00000000;
    rd_cycle[12254] = 1'b0;  wr_cycle[12254] = 1'b1;  addr_rom[12254]='h000015f0;  wr_data_rom[12254]='h000011b5;
    rd_cycle[12255] = 1'b0;  wr_cycle[12255] = 1'b1;  addr_rom[12255]='h0000216c;  wr_data_rom[12255]='h000021ed;
    rd_cycle[12256] = 1'b1;  wr_cycle[12256] = 1'b0;  addr_rom[12256]='h0000048c;  wr_data_rom[12256]='h00000000;
    rd_cycle[12257] = 1'b1;  wr_cycle[12257] = 1'b0;  addr_rom[12257]='h00001a9c;  wr_data_rom[12257]='h00000000;
    rd_cycle[12258] = 1'b1;  wr_cycle[12258] = 1'b0;  addr_rom[12258]='h00002bd4;  wr_data_rom[12258]='h00000000;
    rd_cycle[12259] = 1'b1;  wr_cycle[12259] = 1'b0;  addr_rom[12259]='h0000134c;  wr_data_rom[12259]='h00000000;
    rd_cycle[12260] = 1'b1;  wr_cycle[12260] = 1'b0;  addr_rom[12260]='h00000474;  wr_data_rom[12260]='h00000000;
    rd_cycle[12261] = 1'b1;  wr_cycle[12261] = 1'b0;  addr_rom[12261]='h00001510;  wr_data_rom[12261]='h00000000;
    rd_cycle[12262] = 1'b1;  wr_cycle[12262] = 1'b0;  addr_rom[12262]='h00001ab0;  wr_data_rom[12262]='h00000000;
    rd_cycle[12263] = 1'b1;  wr_cycle[12263] = 1'b0;  addr_rom[12263]='h00000ff0;  wr_data_rom[12263]='h00000000;
    rd_cycle[12264] = 1'b0;  wr_cycle[12264] = 1'b1;  addr_rom[12264]='h00001540;  wr_data_rom[12264]='h0000261e;
    rd_cycle[12265] = 1'b0;  wr_cycle[12265] = 1'b1;  addr_rom[12265]='h00002bb0;  wr_data_rom[12265]='h000029bf;
    rd_cycle[12266] = 1'b1;  wr_cycle[12266] = 1'b0;  addr_rom[12266]='h000034bc;  wr_data_rom[12266]='h00000000;
    rd_cycle[12267] = 1'b1;  wr_cycle[12267] = 1'b0;  addr_rom[12267]='h00002b20;  wr_data_rom[12267]='h00000000;
    rd_cycle[12268] = 1'b0;  wr_cycle[12268] = 1'b1;  addr_rom[12268]='h0000326c;  wr_data_rom[12268]='h000007b2;
    rd_cycle[12269] = 1'b1;  wr_cycle[12269] = 1'b0;  addr_rom[12269]='h00000108;  wr_data_rom[12269]='h00000000;
    rd_cycle[12270] = 1'b0;  wr_cycle[12270] = 1'b1;  addr_rom[12270]='h00001008;  wr_data_rom[12270]='h0000340f;
    rd_cycle[12271] = 1'b1;  wr_cycle[12271] = 1'b0;  addr_rom[12271]='h0000249c;  wr_data_rom[12271]='h00000000;
    rd_cycle[12272] = 1'b1;  wr_cycle[12272] = 1'b0;  addr_rom[12272]='h000024f4;  wr_data_rom[12272]='h00000000;
    rd_cycle[12273] = 1'b0;  wr_cycle[12273] = 1'b1;  addr_rom[12273]='h00002e70;  wr_data_rom[12273]='h000000fc;
    rd_cycle[12274] = 1'b0;  wr_cycle[12274] = 1'b1;  addr_rom[12274]='h000002ec;  wr_data_rom[12274]='h00002bd1;
    rd_cycle[12275] = 1'b0;  wr_cycle[12275] = 1'b1;  addr_rom[12275]='h00001b68;  wr_data_rom[12275]='h00002081;
    rd_cycle[12276] = 1'b1;  wr_cycle[12276] = 1'b0;  addr_rom[12276]='h000006a4;  wr_data_rom[12276]='h00000000;
    rd_cycle[12277] = 1'b0;  wr_cycle[12277] = 1'b1;  addr_rom[12277]='h000028dc;  wr_data_rom[12277]='h000015a2;
    rd_cycle[12278] = 1'b1;  wr_cycle[12278] = 1'b0;  addr_rom[12278]='h00000090;  wr_data_rom[12278]='h00000000;
    rd_cycle[12279] = 1'b0;  wr_cycle[12279] = 1'b1;  addr_rom[12279]='h00003580;  wr_data_rom[12279]='h00003752;
    rd_cycle[12280] = 1'b0;  wr_cycle[12280] = 1'b1;  addr_rom[12280]='h00002398;  wr_data_rom[12280]='h000000a3;
    rd_cycle[12281] = 1'b0;  wr_cycle[12281] = 1'b1;  addr_rom[12281]='h000028b0;  wr_data_rom[12281]='h0000151b;
    rd_cycle[12282] = 1'b0;  wr_cycle[12282] = 1'b1;  addr_rom[12282]='h00003e28;  wr_data_rom[12282]='h00003731;
    rd_cycle[12283] = 1'b1;  wr_cycle[12283] = 1'b0;  addr_rom[12283]='h00000b80;  wr_data_rom[12283]='h00000000;
    rd_cycle[12284] = 1'b1;  wr_cycle[12284] = 1'b0;  addr_rom[12284]='h00001e44;  wr_data_rom[12284]='h00000000;
    rd_cycle[12285] = 1'b0;  wr_cycle[12285] = 1'b1;  addr_rom[12285]='h00002638;  wr_data_rom[12285]='h000006ff;
    rd_cycle[12286] = 1'b0;  wr_cycle[12286] = 1'b1;  addr_rom[12286]='h0000233c;  wr_data_rom[12286]='h000037b1;
    rd_cycle[12287] = 1'b1;  wr_cycle[12287] = 1'b0;  addr_rom[12287]='h00003c94;  wr_data_rom[12287]='h00000000;
    rd_cycle[12288] = 1'b1;  wr_cycle[12288] = 1'b0;  addr_rom[12288]='h00001d50;  wr_data_rom[12288]='h00000000;
    rd_cycle[12289] = 1'b0;  wr_cycle[12289] = 1'b1;  addr_rom[12289]='h00001bac;  wr_data_rom[12289]='h00003476;
    rd_cycle[12290] = 1'b1;  wr_cycle[12290] = 1'b0;  addr_rom[12290]='h00003db4;  wr_data_rom[12290]='h00000000;
    rd_cycle[12291] = 1'b0;  wr_cycle[12291] = 1'b1;  addr_rom[12291]='h00001c38;  wr_data_rom[12291]='h00002e80;
    rd_cycle[12292] = 1'b0;  wr_cycle[12292] = 1'b1;  addr_rom[12292]='h000014dc;  wr_data_rom[12292]='h000016b1;
    rd_cycle[12293] = 1'b1;  wr_cycle[12293] = 1'b0;  addr_rom[12293]='h00001634;  wr_data_rom[12293]='h00000000;
    rd_cycle[12294] = 1'b0;  wr_cycle[12294] = 1'b1;  addr_rom[12294]='h00001984;  wr_data_rom[12294]='h00001d4b;
    rd_cycle[12295] = 1'b0;  wr_cycle[12295] = 1'b1;  addr_rom[12295]='h00003c40;  wr_data_rom[12295]='h00003f5f;
    rd_cycle[12296] = 1'b0;  wr_cycle[12296] = 1'b1;  addr_rom[12296]='h000011c4;  wr_data_rom[12296]='h000004b9;
    rd_cycle[12297] = 1'b1;  wr_cycle[12297] = 1'b0;  addr_rom[12297]='h00001a60;  wr_data_rom[12297]='h00000000;
    rd_cycle[12298] = 1'b0;  wr_cycle[12298] = 1'b1;  addr_rom[12298]='h00000764;  wr_data_rom[12298]='h00002aed;
    rd_cycle[12299] = 1'b0;  wr_cycle[12299] = 1'b1;  addr_rom[12299]='h00003180;  wr_data_rom[12299]='h00002a70;
    rd_cycle[12300] = 1'b1;  wr_cycle[12300] = 1'b0;  addr_rom[12300]='h00003180;  wr_data_rom[12300]='h00000000;
    rd_cycle[12301] = 1'b0;  wr_cycle[12301] = 1'b1;  addr_rom[12301]='h0000373c;  wr_data_rom[12301]='h00002b56;
    rd_cycle[12302] = 1'b1;  wr_cycle[12302] = 1'b0;  addr_rom[12302]='h00003e48;  wr_data_rom[12302]='h00000000;
    rd_cycle[12303] = 1'b1;  wr_cycle[12303] = 1'b0;  addr_rom[12303]='h00003e10;  wr_data_rom[12303]='h00000000;
    rd_cycle[12304] = 1'b0;  wr_cycle[12304] = 1'b1;  addr_rom[12304]='h00002e20;  wr_data_rom[12304]='h000031cb;
    rd_cycle[12305] = 1'b0;  wr_cycle[12305] = 1'b1;  addr_rom[12305]='h000032e8;  wr_data_rom[12305]='h0000352e;
    rd_cycle[12306] = 1'b1;  wr_cycle[12306] = 1'b0;  addr_rom[12306]='h00002280;  wr_data_rom[12306]='h00000000;
    rd_cycle[12307] = 1'b0;  wr_cycle[12307] = 1'b1;  addr_rom[12307]='h00003d08;  wr_data_rom[12307]='h000010ad;
    rd_cycle[12308] = 1'b0;  wr_cycle[12308] = 1'b1;  addr_rom[12308]='h00000244;  wr_data_rom[12308]='h00002685;
    rd_cycle[12309] = 1'b1;  wr_cycle[12309] = 1'b0;  addr_rom[12309]='h000010b4;  wr_data_rom[12309]='h00000000;
    rd_cycle[12310] = 1'b0;  wr_cycle[12310] = 1'b1;  addr_rom[12310]='h00001324;  wr_data_rom[12310]='h00000c8c;
    rd_cycle[12311] = 1'b1;  wr_cycle[12311] = 1'b0;  addr_rom[12311]='h00001c60;  wr_data_rom[12311]='h00000000;
    rd_cycle[12312] = 1'b0;  wr_cycle[12312] = 1'b1;  addr_rom[12312]='h000037ec;  wr_data_rom[12312]='h0000212a;
    rd_cycle[12313] = 1'b0;  wr_cycle[12313] = 1'b1;  addr_rom[12313]='h00000d9c;  wr_data_rom[12313]='h00002468;
    rd_cycle[12314] = 1'b0;  wr_cycle[12314] = 1'b1;  addr_rom[12314]='h00002014;  wr_data_rom[12314]='h000018a7;
    rd_cycle[12315] = 1'b1;  wr_cycle[12315] = 1'b0;  addr_rom[12315]='h0000395c;  wr_data_rom[12315]='h00000000;
    rd_cycle[12316] = 1'b0;  wr_cycle[12316] = 1'b1;  addr_rom[12316]='h00003980;  wr_data_rom[12316]='h000028bb;
    rd_cycle[12317] = 1'b0;  wr_cycle[12317] = 1'b1;  addr_rom[12317]='h0000256c;  wr_data_rom[12317]='h00002223;
    rd_cycle[12318] = 1'b1;  wr_cycle[12318] = 1'b0;  addr_rom[12318]='h00003758;  wr_data_rom[12318]='h00000000;
    rd_cycle[12319] = 1'b0;  wr_cycle[12319] = 1'b1;  addr_rom[12319]='h00001b24;  wr_data_rom[12319]='h00000408;
    rd_cycle[12320] = 1'b1;  wr_cycle[12320] = 1'b0;  addr_rom[12320]='h000029b4;  wr_data_rom[12320]='h00000000;
    rd_cycle[12321] = 1'b1;  wr_cycle[12321] = 1'b0;  addr_rom[12321]='h00000cc4;  wr_data_rom[12321]='h00000000;
    rd_cycle[12322] = 1'b0;  wr_cycle[12322] = 1'b1;  addr_rom[12322]='h00003008;  wr_data_rom[12322]='h000006f9;
    rd_cycle[12323] = 1'b0;  wr_cycle[12323] = 1'b1;  addr_rom[12323]='h00000b34;  wr_data_rom[12323]='h000011d4;
    rd_cycle[12324] = 1'b0;  wr_cycle[12324] = 1'b1;  addr_rom[12324]='h000000fc;  wr_data_rom[12324]='h00000fe5;
    rd_cycle[12325] = 1'b1;  wr_cycle[12325] = 1'b0;  addr_rom[12325]='h00001660;  wr_data_rom[12325]='h00000000;
    rd_cycle[12326] = 1'b1;  wr_cycle[12326] = 1'b0;  addr_rom[12326]='h000016e0;  wr_data_rom[12326]='h00000000;
    rd_cycle[12327] = 1'b0;  wr_cycle[12327] = 1'b1;  addr_rom[12327]='h00001830;  wr_data_rom[12327]='h00000b5a;
    rd_cycle[12328] = 1'b0;  wr_cycle[12328] = 1'b1;  addr_rom[12328]='h00003a74;  wr_data_rom[12328]='h00001c91;
    rd_cycle[12329] = 1'b1;  wr_cycle[12329] = 1'b0;  addr_rom[12329]='h00000eec;  wr_data_rom[12329]='h00000000;
    rd_cycle[12330] = 1'b0;  wr_cycle[12330] = 1'b1;  addr_rom[12330]='h00001628;  wr_data_rom[12330]='h00002909;
    rd_cycle[12331] = 1'b0;  wr_cycle[12331] = 1'b1;  addr_rom[12331]='h00002f38;  wr_data_rom[12331]='h00003854;
    rd_cycle[12332] = 1'b0;  wr_cycle[12332] = 1'b1;  addr_rom[12332]='h0000006c;  wr_data_rom[12332]='h000033e3;
    rd_cycle[12333] = 1'b1;  wr_cycle[12333] = 1'b0;  addr_rom[12333]='h00002d5c;  wr_data_rom[12333]='h00000000;
    rd_cycle[12334] = 1'b1;  wr_cycle[12334] = 1'b0;  addr_rom[12334]='h00002d60;  wr_data_rom[12334]='h00000000;
    rd_cycle[12335] = 1'b1;  wr_cycle[12335] = 1'b0;  addr_rom[12335]='h00002a54;  wr_data_rom[12335]='h00000000;
    rd_cycle[12336] = 1'b1;  wr_cycle[12336] = 1'b0;  addr_rom[12336]='h000031b4;  wr_data_rom[12336]='h00000000;
    rd_cycle[12337] = 1'b1;  wr_cycle[12337] = 1'b0;  addr_rom[12337]='h00000c14;  wr_data_rom[12337]='h00000000;
    rd_cycle[12338] = 1'b1;  wr_cycle[12338] = 1'b0;  addr_rom[12338]='h0000216c;  wr_data_rom[12338]='h00000000;
    rd_cycle[12339] = 1'b0;  wr_cycle[12339] = 1'b1;  addr_rom[12339]='h0000339c;  wr_data_rom[12339]='h00003d68;
    rd_cycle[12340] = 1'b0;  wr_cycle[12340] = 1'b1;  addr_rom[12340]='h0000309c;  wr_data_rom[12340]='h00003a6e;
    rd_cycle[12341] = 1'b1;  wr_cycle[12341] = 1'b0;  addr_rom[12341]='h000027ec;  wr_data_rom[12341]='h00000000;
    rd_cycle[12342] = 1'b0;  wr_cycle[12342] = 1'b1;  addr_rom[12342]='h000038c4;  wr_data_rom[12342]='h0000291b;
    rd_cycle[12343] = 1'b1;  wr_cycle[12343] = 1'b0;  addr_rom[12343]='h000031d0;  wr_data_rom[12343]='h00000000;
    rd_cycle[12344] = 1'b1;  wr_cycle[12344] = 1'b0;  addr_rom[12344]='h00002240;  wr_data_rom[12344]='h00000000;
    rd_cycle[12345] = 1'b0;  wr_cycle[12345] = 1'b1;  addr_rom[12345]='h00003f68;  wr_data_rom[12345]='h0000146d;
    rd_cycle[12346] = 1'b0;  wr_cycle[12346] = 1'b1;  addr_rom[12346]='h00003290;  wr_data_rom[12346]='h00003790;
    rd_cycle[12347] = 1'b1;  wr_cycle[12347] = 1'b0;  addr_rom[12347]='h00002678;  wr_data_rom[12347]='h00000000;
    rd_cycle[12348] = 1'b0;  wr_cycle[12348] = 1'b1;  addr_rom[12348]='h00003324;  wr_data_rom[12348]='h000009fc;
    rd_cycle[12349] = 1'b0;  wr_cycle[12349] = 1'b1;  addr_rom[12349]='h000020cc;  wr_data_rom[12349]='h0000156c;
    rd_cycle[12350] = 1'b0;  wr_cycle[12350] = 1'b1;  addr_rom[12350]='h000039a0;  wr_data_rom[12350]='h00002ab6;
    rd_cycle[12351] = 1'b0;  wr_cycle[12351] = 1'b1;  addr_rom[12351]='h000003c8;  wr_data_rom[12351]='h0000183c;
    rd_cycle[12352] = 1'b1;  wr_cycle[12352] = 1'b0;  addr_rom[12352]='h0000219c;  wr_data_rom[12352]='h00000000;
    rd_cycle[12353] = 1'b0;  wr_cycle[12353] = 1'b1;  addr_rom[12353]='h00001ad0;  wr_data_rom[12353]='h000014e9;
    rd_cycle[12354] = 1'b1;  wr_cycle[12354] = 1'b0;  addr_rom[12354]='h000018a8;  wr_data_rom[12354]='h00000000;
    rd_cycle[12355] = 1'b1;  wr_cycle[12355] = 1'b0;  addr_rom[12355]='h000037d8;  wr_data_rom[12355]='h00000000;
    rd_cycle[12356] = 1'b1;  wr_cycle[12356] = 1'b0;  addr_rom[12356]='h00001348;  wr_data_rom[12356]='h00000000;
    rd_cycle[12357] = 1'b1;  wr_cycle[12357] = 1'b0;  addr_rom[12357]='h00000828;  wr_data_rom[12357]='h00000000;
    rd_cycle[12358] = 1'b0;  wr_cycle[12358] = 1'b1;  addr_rom[12358]='h00002714;  wr_data_rom[12358]='h000008d4;
    rd_cycle[12359] = 1'b0;  wr_cycle[12359] = 1'b1;  addr_rom[12359]='h00000c10;  wr_data_rom[12359]='h00000b46;
    rd_cycle[12360] = 1'b1;  wr_cycle[12360] = 1'b0;  addr_rom[12360]='h00003740;  wr_data_rom[12360]='h00000000;
    rd_cycle[12361] = 1'b1;  wr_cycle[12361] = 1'b0;  addr_rom[12361]='h000023e4;  wr_data_rom[12361]='h00000000;
    rd_cycle[12362] = 1'b1;  wr_cycle[12362] = 1'b0;  addr_rom[12362]='h00001a50;  wr_data_rom[12362]='h00000000;
    rd_cycle[12363] = 1'b1;  wr_cycle[12363] = 1'b0;  addr_rom[12363]='h00000908;  wr_data_rom[12363]='h00000000;
    rd_cycle[12364] = 1'b0;  wr_cycle[12364] = 1'b1;  addr_rom[12364]='h000015e0;  wr_data_rom[12364]='h000015e4;
    rd_cycle[12365] = 1'b1;  wr_cycle[12365] = 1'b0;  addr_rom[12365]='h00003ff0;  wr_data_rom[12365]='h00000000;
    rd_cycle[12366] = 1'b1;  wr_cycle[12366] = 1'b0;  addr_rom[12366]='h000009f4;  wr_data_rom[12366]='h00000000;
    rd_cycle[12367] = 1'b0;  wr_cycle[12367] = 1'b1;  addr_rom[12367]='h00000278;  wr_data_rom[12367]='h00001803;
    rd_cycle[12368] = 1'b0;  wr_cycle[12368] = 1'b1;  addr_rom[12368]='h00003284;  wr_data_rom[12368]='h00000373;
    rd_cycle[12369] = 1'b0;  wr_cycle[12369] = 1'b1;  addr_rom[12369]='h00002060;  wr_data_rom[12369]='h0000192e;
    rd_cycle[12370] = 1'b0;  wr_cycle[12370] = 1'b1;  addr_rom[12370]='h00001d74;  wr_data_rom[12370]='h0000070b;
    rd_cycle[12371] = 1'b0;  wr_cycle[12371] = 1'b1;  addr_rom[12371]='h00001ce4;  wr_data_rom[12371]='h000009e4;
    rd_cycle[12372] = 1'b0;  wr_cycle[12372] = 1'b1;  addr_rom[12372]='h00002db4;  wr_data_rom[12372]='h00000b06;
    rd_cycle[12373] = 1'b0;  wr_cycle[12373] = 1'b1;  addr_rom[12373]='h000038dc;  wr_data_rom[12373]='h000004ff;
    rd_cycle[12374] = 1'b1;  wr_cycle[12374] = 1'b0;  addr_rom[12374]='h000003d0;  wr_data_rom[12374]='h00000000;
    rd_cycle[12375] = 1'b0;  wr_cycle[12375] = 1'b1;  addr_rom[12375]='h00002d74;  wr_data_rom[12375]='h0000351f;
    rd_cycle[12376] = 1'b0;  wr_cycle[12376] = 1'b1;  addr_rom[12376]='h00002768;  wr_data_rom[12376]='h000023de;
    rd_cycle[12377] = 1'b1;  wr_cycle[12377] = 1'b0;  addr_rom[12377]='h00001de0;  wr_data_rom[12377]='h00000000;
    rd_cycle[12378] = 1'b1;  wr_cycle[12378] = 1'b0;  addr_rom[12378]='h00000b78;  wr_data_rom[12378]='h00000000;
    rd_cycle[12379] = 1'b1;  wr_cycle[12379] = 1'b0;  addr_rom[12379]='h000000fc;  wr_data_rom[12379]='h00000000;
    rd_cycle[12380] = 1'b0;  wr_cycle[12380] = 1'b1;  addr_rom[12380]='h00001668;  wr_data_rom[12380]='h00000431;
    rd_cycle[12381] = 1'b0;  wr_cycle[12381] = 1'b1;  addr_rom[12381]='h00000aa8;  wr_data_rom[12381]='h0000316b;
    rd_cycle[12382] = 1'b0;  wr_cycle[12382] = 1'b1;  addr_rom[12382]='h00001a74;  wr_data_rom[12382]='h000003c1;
    rd_cycle[12383] = 1'b0;  wr_cycle[12383] = 1'b1;  addr_rom[12383]='h00003888;  wr_data_rom[12383]='h0000396c;
    rd_cycle[12384] = 1'b1;  wr_cycle[12384] = 1'b0;  addr_rom[12384]='h00000268;  wr_data_rom[12384]='h00000000;
    rd_cycle[12385] = 1'b0;  wr_cycle[12385] = 1'b1;  addr_rom[12385]='h00001770;  wr_data_rom[12385]='h00002233;
    rd_cycle[12386] = 1'b1;  wr_cycle[12386] = 1'b0;  addr_rom[12386]='h000036c8;  wr_data_rom[12386]='h00000000;
    rd_cycle[12387] = 1'b0;  wr_cycle[12387] = 1'b1;  addr_rom[12387]='h00003e7c;  wr_data_rom[12387]='h00001fe6;
    rd_cycle[12388] = 1'b1;  wr_cycle[12388] = 1'b0;  addr_rom[12388]='h00003f00;  wr_data_rom[12388]='h00000000;
    rd_cycle[12389] = 1'b1;  wr_cycle[12389] = 1'b0;  addr_rom[12389]='h00003898;  wr_data_rom[12389]='h00000000;
    rd_cycle[12390] = 1'b0;  wr_cycle[12390] = 1'b1;  addr_rom[12390]='h000009c8;  wr_data_rom[12390]='h0000034c;
    rd_cycle[12391] = 1'b1;  wr_cycle[12391] = 1'b0;  addr_rom[12391]='h00002fd0;  wr_data_rom[12391]='h00000000;
    rd_cycle[12392] = 1'b0;  wr_cycle[12392] = 1'b1;  addr_rom[12392]='h00000a34;  wr_data_rom[12392]='h0000151a;
    rd_cycle[12393] = 1'b0;  wr_cycle[12393] = 1'b1;  addr_rom[12393]='h00002f1c;  wr_data_rom[12393]='h00001df7;
    rd_cycle[12394] = 1'b0;  wr_cycle[12394] = 1'b1;  addr_rom[12394]='h00001a58;  wr_data_rom[12394]='h0000347f;
    rd_cycle[12395] = 1'b1;  wr_cycle[12395] = 1'b0;  addr_rom[12395]='h00001b1c;  wr_data_rom[12395]='h00000000;
    rd_cycle[12396] = 1'b1;  wr_cycle[12396] = 1'b0;  addr_rom[12396]='h00001bb8;  wr_data_rom[12396]='h00000000;
    rd_cycle[12397] = 1'b0;  wr_cycle[12397] = 1'b1;  addr_rom[12397]='h000000bc;  wr_data_rom[12397]='h000012c4;
    rd_cycle[12398] = 1'b0;  wr_cycle[12398] = 1'b1;  addr_rom[12398]='h000009fc;  wr_data_rom[12398]='h000010a4;
    rd_cycle[12399] = 1'b0;  wr_cycle[12399] = 1'b1;  addr_rom[12399]='h00003c68;  wr_data_rom[12399]='h00001389;
    rd_cycle[12400] = 1'b0;  wr_cycle[12400] = 1'b1;  addr_rom[12400]='h00000544;  wr_data_rom[12400]='h0000195b;
    rd_cycle[12401] = 1'b0;  wr_cycle[12401] = 1'b1;  addr_rom[12401]='h00003820;  wr_data_rom[12401]='h000016e0;
    rd_cycle[12402] = 1'b0;  wr_cycle[12402] = 1'b1;  addr_rom[12402]='h00002014;  wr_data_rom[12402]='h0000207b;
    rd_cycle[12403] = 1'b0;  wr_cycle[12403] = 1'b1;  addr_rom[12403]='h0000252c;  wr_data_rom[12403]='h00001461;
    rd_cycle[12404] = 1'b0;  wr_cycle[12404] = 1'b1;  addr_rom[12404]='h00001a98;  wr_data_rom[12404]='h00003fe1;
    rd_cycle[12405] = 1'b1;  wr_cycle[12405] = 1'b0;  addr_rom[12405]='h00003f1c;  wr_data_rom[12405]='h00000000;
    rd_cycle[12406] = 1'b1;  wr_cycle[12406] = 1'b0;  addr_rom[12406]='h00000e08;  wr_data_rom[12406]='h00000000;
    rd_cycle[12407] = 1'b1;  wr_cycle[12407] = 1'b0;  addr_rom[12407]='h00001038;  wr_data_rom[12407]='h00000000;
    rd_cycle[12408] = 1'b0;  wr_cycle[12408] = 1'b1;  addr_rom[12408]='h00003dd0;  wr_data_rom[12408]='h00001f7b;
    rd_cycle[12409] = 1'b1;  wr_cycle[12409] = 1'b0;  addr_rom[12409]='h00002a20;  wr_data_rom[12409]='h00000000;
    rd_cycle[12410] = 1'b0;  wr_cycle[12410] = 1'b1;  addr_rom[12410]='h00002c80;  wr_data_rom[12410]='h0000261e;
    rd_cycle[12411] = 1'b0;  wr_cycle[12411] = 1'b1;  addr_rom[12411]='h00003130;  wr_data_rom[12411]='h00003373;
    rd_cycle[12412] = 1'b0;  wr_cycle[12412] = 1'b1;  addr_rom[12412]='h0000099c;  wr_data_rom[12412]='h00002cb9;
    rd_cycle[12413] = 1'b1;  wr_cycle[12413] = 1'b0;  addr_rom[12413]='h00000d28;  wr_data_rom[12413]='h00000000;
    rd_cycle[12414] = 1'b1;  wr_cycle[12414] = 1'b0;  addr_rom[12414]='h00003b04;  wr_data_rom[12414]='h00000000;
    rd_cycle[12415] = 1'b1;  wr_cycle[12415] = 1'b0;  addr_rom[12415]='h000015c4;  wr_data_rom[12415]='h00000000;
    rd_cycle[12416] = 1'b0;  wr_cycle[12416] = 1'b1;  addr_rom[12416]='h0000136c;  wr_data_rom[12416]='h000031bb;
    rd_cycle[12417] = 1'b1;  wr_cycle[12417] = 1'b0;  addr_rom[12417]='h00003428;  wr_data_rom[12417]='h00000000;
    rd_cycle[12418] = 1'b0;  wr_cycle[12418] = 1'b1;  addr_rom[12418]='h000008f4;  wr_data_rom[12418]='h00002bf5;
    rd_cycle[12419] = 1'b1;  wr_cycle[12419] = 1'b0;  addr_rom[12419]='h00001dd0;  wr_data_rom[12419]='h00000000;
    rd_cycle[12420] = 1'b1;  wr_cycle[12420] = 1'b0;  addr_rom[12420]='h000010b0;  wr_data_rom[12420]='h00000000;
    rd_cycle[12421] = 1'b0;  wr_cycle[12421] = 1'b1;  addr_rom[12421]='h000018c8;  wr_data_rom[12421]='h00000813;
    rd_cycle[12422] = 1'b1;  wr_cycle[12422] = 1'b0;  addr_rom[12422]='h00003db4;  wr_data_rom[12422]='h00000000;
    rd_cycle[12423] = 1'b0;  wr_cycle[12423] = 1'b1;  addr_rom[12423]='h00001e00;  wr_data_rom[12423]='h0000317c;
    rd_cycle[12424] = 1'b1;  wr_cycle[12424] = 1'b0;  addr_rom[12424]='h00001a54;  wr_data_rom[12424]='h00000000;
    rd_cycle[12425] = 1'b1;  wr_cycle[12425] = 1'b0;  addr_rom[12425]='h000000ac;  wr_data_rom[12425]='h00000000;
    rd_cycle[12426] = 1'b1;  wr_cycle[12426] = 1'b0;  addr_rom[12426]='h00003988;  wr_data_rom[12426]='h00000000;
    rd_cycle[12427] = 1'b1;  wr_cycle[12427] = 1'b0;  addr_rom[12427]='h000002e4;  wr_data_rom[12427]='h00000000;
    rd_cycle[12428] = 1'b0;  wr_cycle[12428] = 1'b1;  addr_rom[12428]='h0000150c;  wr_data_rom[12428]='h00002100;
    rd_cycle[12429] = 1'b0;  wr_cycle[12429] = 1'b1;  addr_rom[12429]='h00001fc0;  wr_data_rom[12429]='h00000621;
    rd_cycle[12430] = 1'b0;  wr_cycle[12430] = 1'b1;  addr_rom[12430]='h00001ae0;  wr_data_rom[12430]='h0000093f;
    rd_cycle[12431] = 1'b1;  wr_cycle[12431] = 1'b0;  addr_rom[12431]='h00003c4c;  wr_data_rom[12431]='h00000000;
    rd_cycle[12432] = 1'b1;  wr_cycle[12432] = 1'b0;  addr_rom[12432]='h00000e8c;  wr_data_rom[12432]='h00000000;
    rd_cycle[12433] = 1'b1;  wr_cycle[12433] = 1'b0;  addr_rom[12433]='h00003b48;  wr_data_rom[12433]='h00000000;
    rd_cycle[12434] = 1'b0;  wr_cycle[12434] = 1'b1;  addr_rom[12434]='h00003354;  wr_data_rom[12434]='h000036a8;
    rd_cycle[12435] = 1'b0;  wr_cycle[12435] = 1'b1;  addr_rom[12435]='h00003e14;  wr_data_rom[12435]='h00001f6b;
    rd_cycle[12436] = 1'b0;  wr_cycle[12436] = 1'b1;  addr_rom[12436]='h00002f70;  wr_data_rom[12436]='h00002b68;
    rd_cycle[12437] = 1'b0;  wr_cycle[12437] = 1'b1;  addr_rom[12437]='h00002030;  wr_data_rom[12437]='h0000307c;
    rd_cycle[12438] = 1'b0;  wr_cycle[12438] = 1'b1;  addr_rom[12438]='h00000430;  wr_data_rom[12438]='h00001ac4;
    rd_cycle[12439] = 1'b1;  wr_cycle[12439] = 1'b0;  addr_rom[12439]='h000039ac;  wr_data_rom[12439]='h00000000;
    rd_cycle[12440] = 1'b1;  wr_cycle[12440] = 1'b0;  addr_rom[12440]='h00002d34;  wr_data_rom[12440]='h00000000;
    rd_cycle[12441] = 1'b1;  wr_cycle[12441] = 1'b0;  addr_rom[12441]='h00003264;  wr_data_rom[12441]='h00000000;
    rd_cycle[12442] = 1'b1;  wr_cycle[12442] = 1'b0;  addr_rom[12442]='h000003e4;  wr_data_rom[12442]='h00000000;
    rd_cycle[12443] = 1'b1;  wr_cycle[12443] = 1'b0;  addr_rom[12443]='h00001140;  wr_data_rom[12443]='h00000000;
    rd_cycle[12444] = 1'b0;  wr_cycle[12444] = 1'b1;  addr_rom[12444]='h0000022c;  wr_data_rom[12444]='h000006af;
    rd_cycle[12445] = 1'b1;  wr_cycle[12445] = 1'b0;  addr_rom[12445]='h00001608;  wr_data_rom[12445]='h00000000;
    rd_cycle[12446] = 1'b1;  wr_cycle[12446] = 1'b0;  addr_rom[12446]='h0000061c;  wr_data_rom[12446]='h00000000;
    rd_cycle[12447] = 1'b0;  wr_cycle[12447] = 1'b1;  addr_rom[12447]='h00001ef0;  wr_data_rom[12447]='h000036fb;
    rd_cycle[12448] = 1'b1;  wr_cycle[12448] = 1'b0;  addr_rom[12448]='h000001ac;  wr_data_rom[12448]='h00000000;
    rd_cycle[12449] = 1'b0;  wr_cycle[12449] = 1'b1;  addr_rom[12449]='h00001dd0;  wr_data_rom[12449]='h00001340;
    rd_cycle[12450] = 1'b1;  wr_cycle[12450] = 1'b0;  addr_rom[12450]='h000030a0;  wr_data_rom[12450]='h00000000;
    rd_cycle[12451] = 1'b1;  wr_cycle[12451] = 1'b0;  addr_rom[12451]='h0000391c;  wr_data_rom[12451]='h00000000;
    rd_cycle[12452] = 1'b0;  wr_cycle[12452] = 1'b1;  addr_rom[12452]='h00003ce4;  wr_data_rom[12452]='h000000cc;
    rd_cycle[12453] = 1'b0;  wr_cycle[12453] = 1'b1;  addr_rom[12453]='h000010c8;  wr_data_rom[12453]='h00003738;
    rd_cycle[12454] = 1'b1;  wr_cycle[12454] = 1'b0;  addr_rom[12454]='h000023c0;  wr_data_rom[12454]='h00000000;
    rd_cycle[12455] = 1'b0;  wr_cycle[12455] = 1'b1;  addr_rom[12455]='h00002970;  wr_data_rom[12455]='h00000e61;
    rd_cycle[12456] = 1'b1;  wr_cycle[12456] = 1'b0;  addr_rom[12456]='h0000347c;  wr_data_rom[12456]='h00000000;
    rd_cycle[12457] = 1'b1;  wr_cycle[12457] = 1'b0;  addr_rom[12457]='h00003658;  wr_data_rom[12457]='h00000000;
    rd_cycle[12458] = 1'b0;  wr_cycle[12458] = 1'b1;  addr_rom[12458]='h00000adc;  wr_data_rom[12458]='h0000257e;
    rd_cycle[12459] = 1'b0;  wr_cycle[12459] = 1'b1;  addr_rom[12459]='h00000434;  wr_data_rom[12459]='h00002c03;
    rd_cycle[12460] = 1'b1;  wr_cycle[12460] = 1'b0;  addr_rom[12460]='h000018d8;  wr_data_rom[12460]='h00000000;
    rd_cycle[12461] = 1'b1;  wr_cycle[12461] = 1'b0;  addr_rom[12461]='h00003a70;  wr_data_rom[12461]='h00000000;
    rd_cycle[12462] = 1'b1;  wr_cycle[12462] = 1'b0;  addr_rom[12462]='h00001e98;  wr_data_rom[12462]='h00000000;
    rd_cycle[12463] = 1'b1;  wr_cycle[12463] = 1'b0;  addr_rom[12463]='h00002e38;  wr_data_rom[12463]='h00000000;
    rd_cycle[12464] = 1'b1;  wr_cycle[12464] = 1'b0;  addr_rom[12464]='h00001984;  wr_data_rom[12464]='h00000000;
    rd_cycle[12465] = 1'b0;  wr_cycle[12465] = 1'b1;  addr_rom[12465]='h00003ad8;  wr_data_rom[12465]='h000016aa;
    rd_cycle[12466] = 1'b0;  wr_cycle[12466] = 1'b1;  addr_rom[12466]='h00000eb8;  wr_data_rom[12466]='h0000034a;
    rd_cycle[12467] = 1'b1;  wr_cycle[12467] = 1'b0;  addr_rom[12467]='h00000044;  wr_data_rom[12467]='h00000000;
    rd_cycle[12468] = 1'b0;  wr_cycle[12468] = 1'b1;  addr_rom[12468]='h00000b44;  wr_data_rom[12468]='h000012f7;
    rd_cycle[12469] = 1'b0;  wr_cycle[12469] = 1'b1;  addr_rom[12469]='h00000c20;  wr_data_rom[12469]='h0000035a;
    rd_cycle[12470] = 1'b0;  wr_cycle[12470] = 1'b1;  addr_rom[12470]='h0000170c;  wr_data_rom[12470]='h000032b9;
    rd_cycle[12471] = 1'b0;  wr_cycle[12471] = 1'b1;  addr_rom[12471]='h00002abc;  wr_data_rom[12471]='h0000181d;
    rd_cycle[12472] = 1'b0;  wr_cycle[12472] = 1'b1;  addr_rom[12472]='h00002b38;  wr_data_rom[12472]='h00002cf5;
    rd_cycle[12473] = 1'b0;  wr_cycle[12473] = 1'b1;  addr_rom[12473]='h00003978;  wr_data_rom[12473]='h00003d51;
    rd_cycle[12474] = 1'b0;  wr_cycle[12474] = 1'b1;  addr_rom[12474]='h00001cc0;  wr_data_rom[12474]='h00001243;
    rd_cycle[12475] = 1'b0;  wr_cycle[12475] = 1'b1;  addr_rom[12475]='h00003320;  wr_data_rom[12475]='h00002026;
    rd_cycle[12476] = 1'b1;  wr_cycle[12476] = 1'b0;  addr_rom[12476]='h00003138;  wr_data_rom[12476]='h00000000;
    rd_cycle[12477] = 1'b1;  wr_cycle[12477] = 1'b0;  addr_rom[12477]='h000022d8;  wr_data_rom[12477]='h00000000;
    rd_cycle[12478] = 1'b0;  wr_cycle[12478] = 1'b1;  addr_rom[12478]='h0000350c;  wr_data_rom[12478]='h00003557;
    rd_cycle[12479] = 1'b1;  wr_cycle[12479] = 1'b0;  addr_rom[12479]='h00000f54;  wr_data_rom[12479]='h00000000;
    rd_cycle[12480] = 1'b1;  wr_cycle[12480] = 1'b0;  addr_rom[12480]='h0000378c;  wr_data_rom[12480]='h00000000;
    rd_cycle[12481] = 1'b1;  wr_cycle[12481] = 1'b0;  addr_rom[12481]='h000015b0;  wr_data_rom[12481]='h00000000;
    rd_cycle[12482] = 1'b1;  wr_cycle[12482] = 1'b0;  addr_rom[12482]='h00002050;  wr_data_rom[12482]='h00000000;
    rd_cycle[12483] = 1'b0;  wr_cycle[12483] = 1'b1;  addr_rom[12483]='h00002538;  wr_data_rom[12483]='h0000167f;
    rd_cycle[12484] = 1'b1;  wr_cycle[12484] = 1'b0;  addr_rom[12484]='h00002298;  wr_data_rom[12484]='h00000000;
    rd_cycle[12485] = 1'b0;  wr_cycle[12485] = 1'b1;  addr_rom[12485]='h000015a8;  wr_data_rom[12485]='h000001e9;
    rd_cycle[12486] = 1'b1;  wr_cycle[12486] = 1'b0;  addr_rom[12486]='h00003624;  wr_data_rom[12486]='h00000000;
    rd_cycle[12487] = 1'b0;  wr_cycle[12487] = 1'b1;  addr_rom[12487]='h000004f8;  wr_data_rom[12487]='h000010f4;
    rd_cycle[12488] = 1'b1;  wr_cycle[12488] = 1'b0;  addr_rom[12488]='h000034c8;  wr_data_rom[12488]='h00000000;
    rd_cycle[12489] = 1'b1;  wr_cycle[12489] = 1'b0;  addr_rom[12489]='h000003fc;  wr_data_rom[12489]='h00000000;
    rd_cycle[12490] = 1'b0;  wr_cycle[12490] = 1'b1;  addr_rom[12490]='h00001924;  wr_data_rom[12490]='h000009ed;
    rd_cycle[12491] = 1'b1;  wr_cycle[12491] = 1'b0;  addr_rom[12491]='h00003b70;  wr_data_rom[12491]='h00000000;
    rd_cycle[12492] = 1'b1;  wr_cycle[12492] = 1'b0;  addr_rom[12492]='h000008cc;  wr_data_rom[12492]='h00000000;
    rd_cycle[12493] = 1'b0;  wr_cycle[12493] = 1'b1;  addr_rom[12493]='h00003b48;  wr_data_rom[12493]='h000005fc;
    rd_cycle[12494] = 1'b1;  wr_cycle[12494] = 1'b0;  addr_rom[12494]='h00001ba4;  wr_data_rom[12494]='h00000000;
    rd_cycle[12495] = 1'b0;  wr_cycle[12495] = 1'b1;  addr_rom[12495]='h00002ce0;  wr_data_rom[12495]='h00001939;
    rd_cycle[12496] = 1'b0;  wr_cycle[12496] = 1'b1;  addr_rom[12496]='h00001b40;  wr_data_rom[12496]='h0000000c;
    rd_cycle[12497] = 1'b1;  wr_cycle[12497] = 1'b0;  addr_rom[12497]='h0000248c;  wr_data_rom[12497]='h00000000;
    rd_cycle[12498] = 1'b1;  wr_cycle[12498] = 1'b0;  addr_rom[12498]='h00000530;  wr_data_rom[12498]='h00000000;
    rd_cycle[12499] = 1'b0;  wr_cycle[12499] = 1'b1;  addr_rom[12499]='h0000285c;  wr_data_rom[12499]='h00003586;
    rd_cycle[12500] = 1'b0;  wr_cycle[12500] = 1'b1;  addr_rom[12500]='h00003760;  wr_data_rom[12500]='h0000246a;
    rd_cycle[12501] = 1'b1;  wr_cycle[12501] = 1'b0;  addr_rom[12501]='h000024e4;  wr_data_rom[12501]='h00000000;
    rd_cycle[12502] = 1'b0;  wr_cycle[12502] = 1'b1;  addr_rom[12502]='h00000da4;  wr_data_rom[12502]='h00002ee8;
    rd_cycle[12503] = 1'b0;  wr_cycle[12503] = 1'b1;  addr_rom[12503]='h000023a8;  wr_data_rom[12503]='h00001075;
    rd_cycle[12504] = 1'b1;  wr_cycle[12504] = 1'b0;  addr_rom[12504]='h000029ac;  wr_data_rom[12504]='h00000000;
    rd_cycle[12505] = 1'b1;  wr_cycle[12505] = 1'b0;  addr_rom[12505]='h000029a8;  wr_data_rom[12505]='h00000000;
    rd_cycle[12506] = 1'b1;  wr_cycle[12506] = 1'b0;  addr_rom[12506]='h000011a0;  wr_data_rom[12506]='h00000000;
    rd_cycle[12507] = 1'b1;  wr_cycle[12507] = 1'b0;  addr_rom[12507]='h000031c0;  wr_data_rom[12507]='h00000000;
    rd_cycle[12508] = 1'b0;  wr_cycle[12508] = 1'b1;  addr_rom[12508]='h00001050;  wr_data_rom[12508]='h000038aa;
    rd_cycle[12509] = 1'b1;  wr_cycle[12509] = 1'b0;  addr_rom[12509]='h000006f8;  wr_data_rom[12509]='h00000000;
    rd_cycle[12510] = 1'b0;  wr_cycle[12510] = 1'b1;  addr_rom[12510]='h000007fc;  wr_data_rom[12510]='h00003599;
    rd_cycle[12511] = 1'b0;  wr_cycle[12511] = 1'b1;  addr_rom[12511]='h00002c00;  wr_data_rom[12511]='h00002f31;
    rd_cycle[12512] = 1'b0;  wr_cycle[12512] = 1'b1;  addr_rom[12512]='h00000578;  wr_data_rom[12512]='h00003bf0;
    rd_cycle[12513] = 1'b1;  wr_cycle[12513] = 1'b0;  addr_rom[12513]='h00000544;  wr_data_rom[12513]='h00000000;
    rd_cycle[12514] = 1'b1;  wr_cycle[12514] = 1'b0;  addr_rom[12514]='h000034d0;  wr_data_rom[12514]='h00000000;
    rd_cycle[12515] = 1'b0;  wr_cycle[12515] = 1'b1;  addr_rom[12515]='h00000df0;  wr_data_rom[12515]='h00000133;
    rd_cycle[12516] = 1'b0;  wr_cycle[12516] = 1'b1;  addr_rom[12516]='h00003994;  wr_data_rom[12516]='h000031e8;
    rd_cycle[12517] = 1'b1;  wr_cycle[12517] = 1'b0;  addr_rom[12517]='h00001ce8;  wr_data_rom[12517]='h00000000;
    rd_cycle[12518] = 1'b0;  wr_cycle[12518] = 1'b1;  addr_rom[12518]='h00001658;  wr_data_rom[12518]='h00001ded;
    rd_cycle[12519] = 1'b0;  wr_cycle[12519] = 1'b1;  addr_rom[12519]='h00000e2c;  wr_data_rom[12519]='h0000071e;
    rd_cycle[12520] = 1'b0;  wr_cycle[12520] = 1'b1;  addr_rom[12520]='h000018e0;  wr_data_rom[12520]='h00001af3;
    rd_cycle[12521] = 1'b0;  wr_cycle[12521] = 1'b1;  addr_rom[12521]='h00002400;  wr_data_rom[12521]='h00000d16;
    rd_cycle[12522] = 1'b1;  wr_cycle[12522] = 1'b0;  addr_rom[12522]='h000032b8;  wr_data_rom[12522]='h00000000;
    rd_cycle[12523] = 1'b0;  wr_cycle[12523] = 1'b1;  addr_rom[12523]='h00001554;  wr_data_rom[12523]='h00003a7a;
    rd_cycle[12524] = 1'b1;  wr_cycle[12524] = 1'b0;  addr_rom[12524]='h000012cc;  wr_data_rom[12524]='h00000000;
    rd_cycle[12525] = 1'b1;  wr_cycle[12525] = 1'b0;  addr_rom[12525]='h0000030c;  wr_data_rom[12525]='h00000000;
    rd_cycle[12526] = 1'b0;  wr_cycle[12526] = 1'b1;  addr_rom[12526]='h000025cc;  wr_data_rom[12526]='h00000dd0;
    rd_cycle[12527] = 1'b1;  wr_cycle[12527] = 1'b0;  addr_rom[12527]='h00000a98;  wr_data_rom[12527]='h00000000;
    rd_cycle[12528] = 1'b0;  wr_cycle[12528] = 1'b1;  addr_rom[12528]='h0000199c;  wr_data_rom[12528]='h000003cb;
    rd_cycle[12529] = 1'b0;  wr_cycle[12529] = 1'b1;  addr_rom[12529]='h00000514;  wr_data_rom[12529]='h000021d0;
    rd_cycle[12530] = 1'b0;  wr_cycle[12530] = 1'b1;  addr_rom[12530]='h00000840;  wr_data_rom[12530]='h00000cf9;
    rd_cycle[12531] = 1'b0;  wr_cycle[12531] = 1'b1;  addr_rom[12531]='h000023d4;  wr_data_rom[12531]='h00003f8e;
    rd_cycle[12532] = 1'b0;  wr_cycle[12532] = 1'b1;  addr_rom[12532]='h0000089c;  wr_data_rom[12532]='h00000c1a;
    rd_cycle[12533] = 1'b1;  wr_cycle[12533] = 1'b0;  addr_rom[12533]='h000031a0;  wr_data_rom[12533]='h00000000;
    rd_cycle[12534] = 1'b1;  wr_cycle[12534] = 1'b0;  addr_rom[12534]='h0000209c;  wr_data_rom[12534]='h00000000;
    rd_cycle[12535] = 1'b0;  wr_cycle[12535] = 1'b1;  addr_rom[12535]='h00003244;  wr_data_rom[12535]='h00002c53;
    rd_cycle[12536] = 1'b1;  wr_cycle[12536] = 1'b0;  addr_rom[12536]='h00001b90;  wr_data_rom[12536]='h00000000;
    rd_cycle[12537] = 1'b1;  wr_cycle[12537] = 1'b0;  addr_rom[12537]='h00002724;  wr_data_rom[12537]='h00000000;
    rd_cycle[12538] = 1'b1;  wr_cycle[12538] = 1'b0;  addr_rom[12538]='h00001688;  wr_data_rom[12538]='h00000000;
    rd_cycle[12539] = 1'b1;  wr_cycle[12539] = 1'b0;  addr_rom[12539]='h0000214c;  wr_data_rom[12539]='h00000000;
    rd_cycle[12540] = 1'b1;  wr_cycle[12540] = 1'b0;  addr_rom[12540]='h000003d8;  wr_data_rom[12540]='h00000000;
    rd_cycle[12541] = 1'b0;  wr_cycle[12541] = 1'b1;  addr_rom[12541]='h00001634;  wr_data_rom[12541]='h00000550;
    rd_cycle[12542] = 1'b0;  wr_cycle[12542] = 1'b1;  addr_rom[12542]='h0000005c;  wr_data_rom[12542]='h00001274;
    rd_cycle[12543] = 1'b0;  wr_cycle[12543] = 1'b1;  addr_rom[12543]='h000013a8;  wr_data_rom[12543]='h00001448;
    rd_cycle[12544] = 1'b0;  wr_cycle[12544] = 1'b1;  addr_rom[12544]='h000007b8;  wr_data_rom[12544]='h00002439;
    rd_cycle[12545] = 1'b1;  wr_cycle[12545] = 1'b0;  addr_rom[12545]='h00002730;  wr_data_rom[12545]='h00000000;
    rd_cycle[12546] = 1'b1;  wr_cycle[12546] = 1'b0;  addr_rom[12546]='h00001688;  wr_data_rom[12546]='h00000000;
    rd_cycle[12547] = 1'b1;  wr_cycle[12547] = 1'b0;  addr_rom[12547]='h00001d34;  wr_data_rom[12547]='h00000000;
    rd_cycle[12548] = 1'b1;  wr_cycle[12548] = 1'b0;  addr_rom[12548]='h0000049c;  wr_data_rom[12548]='h00000000;
    rd_cycle[12549] = 1'b1;  wr_cycle[12549] = 1'b0;  addr_rom[12549]='h00003b30;  wr_data_rom[12549]='h00000000;
    rd_cycle[12550] = 1'b0;  wr_cycle[12550] = 1'b1;  addr_rom[12550]='h00003350;  wr_data_rom[12550]='h00000ce0;
    rd_cycle[12551] = 1'b1;  wr_cycle[12551] = 1'b0;  addr_rom[12551]='h00001774;  wr_data_rom[12551]='h00000000;
    rd_cycle[12552] = 1'b1;  wr_cycle[12552] = 1'b0;  addr_rom[12552]='h00000d00;  wr_data_rom[12552]='h00000000;
    rd_cycle[12553] = 1'b0;  wr_cycle[12553] = 1'b1;  addr_rom[12553]='h00002328;  wr_data_rom[12553]='h000018a1;
    rd_cycle[12554] = 1'b1;  wr_cycle[12554] = 1'b0;  addr_rom[12554]='h0000364c;  wr_data_rom[12554]='h00000000;
    rd_cycle[12555] = 1'b0;  wr_cycle[12555] = 1'b1;  addr_rom[12555]='h00000558;  wr_data_rom[12555]='h00001153;
    rd_cycle[12556] = 1'b1;  wr_cycle[12556] = 1'b0;  addr_rom[12556]='h00003fd4;  wr_data_rom[12556]='h00000000;
    rd_cycle[12557] = 1'b0;  wr_cycle[12557] = 1'b1;  addr_rom[12557]='h0000111c;  wr_data_rom[12557]='h00000813;
    rd_cycle[12558] = 1'b0;  wr_cycle[12558] = 1'b1;  addr_rom[12558]='h00003fbc;  wr_data_rom[12558]='h00003706;
    rd_cycle[12559] = 1'b0;  wr_cycle[12559] = 1'b1;  addr_rom[12559]='h00003f3c;  wr_data_rom[12559]='h0000321e;
    rd_cycle[12560] = 1'b1;  wr_cycle[12560] = 1'b0;  addr_rom[12560]='h00001068;  wr_data_rom[12560]='h00000000;
    rd_cycle[12561] = 1'b0;  wr_cycle[12561] = 1'b1;  addr_rom[12561]='h00003028;  wr_data_rom[12561]='h000013be;
    rd_cycle[12562] = 1'b0;  wr_cycle[12562] = 1'b1;  addr_rom[12562]='h00003570;  wr_data_rom[12562]='h00002e69;
    rd_cycle[12563] = 1'b0;  wr_cycle[12563] = 1'b1;  addr_rom[12563]='h00003648;  wr_data_rom[12563]='h00002d84;
    rd_cycle[12564] = 1'b1;  wr_cycle[12564] = 1'b0;  addr_rom[12564]='h00000c2c;  wr_data_rom[12564]='h00000000;
    rd_cycle[12565] = 1'b0;  wr_cycle[12565] = 1'b1;  addr_rom[12565]='h00003dfc;  wr_data_rom[12565]='h00003321;
    rd_cycle[12566] = 1'b0;  wr_cycle[12566] = 1'b1;  addr_rom[12566]='h00003850;  wr_data_rom[12566]='h00002218;
    rd_cycle[12567] = 1'b1;  wr_cycle[12567] = 1'b0;  addr_rom[12567]='h00003708;  wr_data_rom[12567]='h00000000;
    rd_cycle[12568] = 1'b1;  wr_cycle[12568] = 1'b0;  addr_rom[12568]='h00003aa4;  wr_data_rom[12568]='h00000000;
    rd_cycle[12569] = 1'b0;  wr_cycle[12569] = 1'b1;  addr_rom[12569]='h00002df4;  wr_data_rom[12569]='h00002f6e;
    rd_cycle[12570] = 1'b0;  wr_cycle[12570] = 1'b1;  addr_rom[12570]='h000033f0;  wr_data_rom[12570]='h00003fbc;
    rd_cycle[12571] = 1'b0;  wr_cycle[12571] = 1'b1;  addr_rom[12571]='h00000a04;  wr_data_rom[12571]='h000012de;
    rd_cycle[12572] = 1'b1;  wr_cycle[12572] = 1'b0;  addr_rom[12572]='h00000380;  wr_data_rom[12572]='h00000000;
    rd_cycle[12573] = 1'b0;  wr_cycle[12573] = 1'b1;  addr_rom[12573]='h000023ec;  wr_data_rom[12573]='h00001115;
    rd_cycle[12574] = 1'b0;  wr_cycle[12574] = 1'b1;  addr_rom[12574]='h00000c88;  wr_data_rom[12574]='h00003767;
    rd_cycle[12575] = 1'b0;  wr_cycle[12575] = 1'b1;  addr_rom[12575]='h00002c20;  wr_data_rom[12575]='h00003d65;
    rd_cycle[12576] = 1'b1;  wr_cycle[12576] = 1'b0;  addr_rom[12576]='h000025b4;  wr_data_rom[12576]='h00000000;
    rd_cycle[12577] = 1'b0;  wr_cycle[12577] = 1'b1;  addr_rom[12577]='h00002bd4;  wr_data_rom[12577]='h00003778;
    rd_cycle[12578] = 1'b0;  wr_cycle[12578] = 1'b1;  addr_rom[12578]='h00002364;  wr_data_rom[12578]='h000021f5;
    rd_cycle[12579] = 1'b1;  wr_cycle[12579] = 1'b0;  addr_rom[12579]='h000027ac;  wr_data_rom[12579]='h00000000;
    rd_cycle[12580] = 1'b0;  wr_cycle[12580] = 1'b1;  addr_rom[12580]='h00001d0c;  wr_data_rom[12580]='h000020a9;
    rd_cycle[12581] = 1'b0;  wr_cycle[12581] = 1'b1;  addr_rom[12581]='h00001120;  wr_data_rom[12581]='h00000a21;
    rd_cycle[12582] = 1'b1;  wr_cycle[12582] = 1'b0;  addr_rom[12582]='h00001920;  wr_data_rom[12582]='h00000000;
    rd_cycle[12583] = 1'b0;  wr_cycle[12583] = 1'b1;  addr_rom[12583]='h00002cf8;  wr_data_rom[12583]='h0000080e;
    rd_cycle[12584] = 1'b1;  wr_cycle[12584] = 1'b0;  addr_rom[12584]='h000025ec;  wr_data_rom[12584]='h00000000;
    rd_cycle[12585] = 1'b1;  wr_cycle[12585] = 1'b0;  addr_rom[12585]='h00002768;  wr_data_rom[12585]='h00000000;
    rd_cycle[12586] = 1'b0;  wr_cycle[12586] = 1'b1;  addr_rom[12586]='h000035dc;  wr_data_rom[12586]='h00001891;
    rd_cycle[12587] = 1'b1;  wr_cycle[12587] = 1'b0;  addr_rom[12587]='h000008ec;  wr_data_rom[12587]='h00000000;
    rd_cycle[12588] = 1'b1;  wr_cycle[12588] = 1'b0;  addr_rom[12588]='h000002cc;  wr_data_rom[12588]='h00000000;
    rd_cycle[12589] = 1'b1;  wr_cycle[12589] = 1'b0;  addr_rom[12589]='h0000101c;  wr_data_rom[12589]='h00000000;
    rd_cycle[12590] = 1'b1;  wr_cycle[12590] = 1'b0;  addr_rom[12590]='h00003cfc;  wr_data_rom[12590]='h00000000;
    rd_cycle[12591] = 1'b1;  wr_cycle[12591] = 1'b0;  addr_rom[12591]='h000033cc;  wr_data_rom[12591]='h00000000;
    rd_cycle[12592] = 1'b1;  wr_cycle[12592] = 1'b0;  addr_rom[12592]='h000026c0;  wr_data_rom[12592]='h00000000;
    rd_cycle[12593] = 1'b0;  wr_cycle[12593] = 1'b1;  addr_rom[12593]='h00002cbc;  wr_data_rom[12593]='h000001c2;
    rd_cycle[12594] = 1'b0;  wr_cycle[12594] = 1'b1;  addr_rom[12594]='h00003bbc;  wr_data_rom[12594]='h00001e82;
    rd_cycle[12595] = 1'b1;  wr_cycle[12595] = 1'b0;  addr_rom[12595]='h000023c4;  wr_data_rom[12595]='h00000000;
    rd_cycle[12596] = 1'b0;  wr_cycle[12596] = 1'b1;  addr_rom[12596]='h000030d8;  wr_data_rom[12596]='h00001f4b;
    rd_cycle[12597] = 1'b1;  wr_cycle[12597] = 1'b0;  addr_rom[12597]='h00001cb4;  wr_data_rom[12597]='h00000000;
    rd_cycle[12598] = 1'b0;  wr_cycle[12598] = 1'b1;  addr_rom[12598]='h00000550;  wr_data_rom[12598]='h00001527;
    rd_cycle[12599] = 1'b1;  wr_cycle[12599] = 1'b0;  addr_rom[12599]='h00003018;  wr_data_rom[12599]='h00000000;
    rd_cycle[12600] = 1'b0;  wr_cycle[12600] = 1'b1;  addr_rom[12600]='h00001400;  wr_data_rom[12600]='h00000598;
    rd_cycle[12601] = 1'b1;  wr_cycle[12601] = 1'b0;  addr_rom[12601]='h00001fc8;  wr_data_rom[12601]='h00000000;
    rd_cycle[12602] = 1'b0;  wr_cycle[12602] = 1'b1;  addr_rom[12602]='h000035f8;  wr_data_rom[12602]='h00003311;
    rd_cycle[12603] = 1'b0;  wr_cycle[12603] = 1'b1;  addr_rom[12603]='h000033a4;  wr_data_rom[12603]='h00001d0e;
    rd_cycle[12604] = 1'b1;  wr_cycle[12604] = 1'b0;  addr_rom[12604]='h000020c8;  wr_data_rom[12604]='h00000000;
    rd_cycle[12605] = 1'b0;  wr_cycle[12605] = 1'b1;  addr_rom[12605]='h00000a00;  wr_data_rom[12605]='h0000069a;
    rd_cycle[12606] = 1'b1;  wr_cycle[12606] = 1'b0;  addr_rom[12606]='h00000790;  wr_data_rom[12606]='h00000000;
    rd_cycle[12607] = 1'b0;  wr_cycle[12607] = 1'b1;  addr_rom[12607]='h0000343c;  wr_data_rom[12607]='h00002db1;
    rd_cycle[12608] = 1'b0;  wr_cycle[12608] = 1'b1;  addr_rom[12608]='h00002160;  wr_data_rom[12608]='h00003777;
    rd_cycle[12609] = 1'b1;  wr_cycle[12609] = 1'b0;  addr_rom[12609]='h00002574;  wr_data_rom[12609]='h00000000;
    rd_cycle[12610] = 1'b1;  wr_cycle[12610] = 1'b0;  addr_rom[12610]='h000010f4;  wr_data_rom[12610]='h00000000;
    rd_cycle[12611] = 1'b1;  wr_cycle[12611] = 1'b0;  addr_rom[12611]='h000024d4;  wr_data_rom[12611]='h00000000;
    rd_cycle[12612] = 1'b1;  wr_cycle[12612] = 1'b0;  addr_rom[12612]='h00000af0;  wr_data_rom[12612]='h00000000;
    rd_cycle[12613] = 1'b0;  wr_cycle[12613] = 1'b1;  addr_rom[12613]='h00000e34;  wr_data_rom[12613]='h00002881;
    rd_cycle[12614] = 1'b1;  wr_cycle[12614] = 1'b0;  addr_rom[12614]='h00000b24;  wr_data_rom[12614]='h00000000;
    rd_cycle[12615] = 1'b1;  wr_cycle[12615] = 1'b0;  addr_rom[12615]='h000018ac;  wr_data_rom[12615]='h00000000;
    rd_cycle[12616] = 1'b0;  wr_cycle[12616] = 1'b1;  addr_rom[12616]='h0000080c;  wr_data_rom[12616]='h00000ada;
    rd_cycle[12617] = 1'b1;  wr_cycle[12617] = 1'b0;  addr_rom[12617]='h00003834;  wr_data_rom[12617]='h00000000;
    rd_cycle[12618] = 1'b1;  wr_cycle[12618] = 1'b0;  addr_rom[12618]='h00001f98;  wr_data_rom[12618]='h00000000;
    rd_cycle[12619] = 1'b0;  wr_cycle[12619] = 1'b1;  addr_rom[12619]='h00000f20;  wr_data_rom[12619]='h00000773;
    rd_cycle[12620] = 1'b0;  wr_cycle[12620] = 1'b1;  addr_rom[12620]='h00001d20;  wr_data_rom[12620]='h00001378;
    rd_cycle[12621] = 1'b0;  wr_cycle[12621] = 1'b1;  addr_rom[12621]='h00000508;  wr_data_rom[12621]='h0000160b;
    rd_cycle[12622] = 1'b1;  wr_cycle[12622] = 1'b0;  addr_rom[12622]='h00002cc8;  wr_data_rom[12622]='h00000000;
    rd_cycle[12623] = 1'b0;  wr_cycle[12623] = 1'b1;  addr_rom[12623]='h00000928;  wr_data_rom[12623]='h00003f08;
    rd_cycle[12624] = 1'b1;  wr_cycle[12624] = 1'b0;  addr_rom[12624]='h00003690;  wr_data_rom[12624]='h00000000;
    rd_cycle[12625] = 1'b1;  wr_cycle[12625] = 1'b0;  addr_rom[12625]='h0000385c;  wr_data_rom[12625]='h00000000;
    rd_cycle[12626] = 1'b0;  wr_cycle[12626] = 1'b1;  addr_rom[12626]='h00001380;  wr_data_rom[12626]='h00001127;
    rd_cycle[12627] = 1'b0;  wr_cycle[12627] = 1'b1;  addr_rom[12627]='h00003258;  wr_data_rom[12627]='h00003302;
    rd_cycle[12628] = 1'b0;  wr_cycle[12628] = 1'b1;  addr_rom[12628]='h00002f60;  wr_data_rom[12628]='h0000377c;
    rd_cycle[12629] = 1'b0;  wr_cycle[12629] = 1'b1;  addr_rom[12629]='h00002020;  wr_data_rom[12629]='h00000fde;
    rd_cycle[12630] = 1'b1;  wr_cycle[12630] = 1'b0;  addr_rom[12630]='h00000330;  wr_data_rom[12630]='h00000000;
    rd_cycle[12631] = 1'b0;  wr_cycle[12631] = 1'b1;  addr_rom[12631]='h000025f4;  wr_data_rom[12631]='h000036e8;
    rd_cycle[12632] = 1'b0;  wr_cycle[12632] = 1'b1;  addr_rom[12632]='h000036f0;  wr_data_rom[12632]='h00000f1b;
    rd_cycle[12633] = 1'b0;  wr_cycle[12633] = 1'b1;  addr_rom[12633]='h0000235c;  wr_data_rom[12633]='h0000064f;
    rd_cycle[12634] = 1'b0;  wr_cycle[12634] = 1'b1;  addr_rom[12634]='h0000364c;  wr_data_rom[12634]='h00002fcb;
    rd_cycle[12635] = 1'b1;  wr_cycle[12635] = 1'b0;  addr_rom[12635]='h00003b78;  wr_data_rom[12635]='h00000000;
    rd_cycle[12636] = 1'b1;  wr_cycle[12636] = 1'b0;  addr_rom[12636]='h0000285c;  wr_data_rom[12636]='h00000000;
    rd_cycle[12637] = 1'b1;  wr_cycle[12637] = 1'b0;  addr_rom[12637]='h00003708;  wr_data_rom[12637]='h00000000;
    rd_cycle[12638] = 1'b0;  wr_cycle[12638] = 1'b1;  addr_rom[12638]='h00001aa0;  wr_data_rom[12638]='h00000680;
    rd_cycle[12639] = 1'b1;  wr_cycle[12639] = 1'b0;  addr_rom[12639]='h00002764;  wr_data_rom[12639]='h00000000;
    rd_cycle[12640] = 1'b0;  wr_cycle[12640] = 1'b1;  addr_rom[12640]='h00003960;  wr_data_rom[12640]='h00000942;
    rd_cycle[12641] = 1'b0;  wr_cycle[12641] = 1'b1;  addr_rom[12641]='h00000a4c;  wr_data_rom[12641]='h000027eb;
    rd_cycle[12642] = 1'b0;  wr_cycle[12642] = 1'b1;  addr_rom[12642]='h000023bc;  wr_data_rom[12642]='h00000a80;
    rd_cycle[12643] = 1'b0;  wr_cycle[12643] = 1'b1;  addr_rom[12643]='h000018ec;  wr_data_rom[12643]='h00002fce;
    rd_cycle[12644] = 1'b0;  wr_cycle[12644] = 1'b1;  addr_rom[12644]='h000004a0;  wr_data_rom[12644]='h0000272c;
    rd_cycle[12645] = 1'b1;  wr_cycle[12645] = 1'b0;  addr_rom[12645]='h0000085c;  wr_data_rom[12645]='h00000000;
    rd_cycle[12646] = 1'b0;  wr_cycle[12646] = 1'b1;  addr_rom[12646]='h00000a50;  wr_data_rom[12646]='h000024bd;
    rd_cycle[12647] = 1'b1;  wr_cycle[12647] = 1'b0;  addr_rom[12647]='h00003a48;  wr_data_rom[12647]='h00000000;
    rd_cycle[12648] = 1'b1;  wr_cycle[12648] = 1'b0;  addr_rom[12648]='h00002d50;  wr_data_rom[12648]='h00000000;
    rd_cycle[12649] = 1'b1;  wr_cycle[12649] = 1'b0;  addr_rom[12649]='h000022b4;  wr_data_rom[12649]='h00000000;
    rd_cycle[12650] = 1'b0;  wr_cycle[12650] = 1'b1;  addr_rom[12650]='h00000c4c;  wr_data_rom[12650]='h000003e9;
    rd_cycle[12651] = 1'b1;  wr_cycle[12651] = 1'b0;  addr_rom[12651]='h0000067c;  wr_data_rom[12651]='h00000000;
    rd_cycle[12652] = 1'b1;  wr_cycle[12652] = 1'b0;  addr_rom[12652]='h000032c0;  wr_data_rom[12652]='h00000000;
    rd_cycle[12653] = 1'b1;  wr_cycle[12653] = 1'b0;  addr_rom[12653]='h000000a4;  wr_data_rom[12653]='h00000000;
    rd_cycle[12654] = 1'b0;  wr_cycle[12654] = 1'b1;  addr_rom[12654]='h000001cc;  wr_data_rom[12654]='h000039f8;
    rd_cycle[12655] = 1'b1;  wr_cycle[12655] = 1'b0;  addr_rom[12655]='h000005a4;  wr_data_rom[12655]='h00000000;
    rd_cycle[12656] = 1'b1;  wr_cycle[12656] = 1'b0;  addr_rom[12656]='h000025d0;  wr_data_rom[12656]='h00000000;
    rd_cycle[12657] = 1'b0;  wr_cycle[12657] = 1'b1;  addr_rom[12657]='h00000c04;  wr_data_rom[12657]='h00001540;
    rd_cycle[12658] = 1'b1;  wr_cycle[12658] = 1'b0;  addr_rom[12658]='h00000294;  wr_data_rom[12658]='h00000000;
    rd_cycle[12659] = 1'b1;  wr_cycle[12659] = 1'b0;  addr_rom[12659]='h00000c14;  wr_data_rom[12659]='h00000000;
    rd_cycle[12660] = 1'b0;  wr_cycle[12660] = 1'b1;  addr_rom[12660]='h00003bc4;  wr_data_rom[12660]='h00002218;
    rd_cycle[12661] = 1'b1;  wr_cycle[12661] = 1'b0;  addr_rom[12661]='h00001a48;  wr_data_rom[12661]='h00000000;
    rd_cycle[12662] = 1'b0;  wr_cycle[12662] = 1'b1;  addr_rom[12662]='h000002fc;  wr_data_rom[12662]='h000029bf;
    rd_cycle[12663] = 1'b1;  wr_cycle[12663] = 1'b0;  addr_rom[12663]='h00000c88;  wr_data_rom[12663]='h00000000;
    rd_cycle[12664] = 1'b1;  wr_cycle[12664] = 1'b0;  addr_rom[12664]='h00002c60;  wr_data_rom[12664]='h00000000;
    rd_cycle[12665] = 1'b0;  wr_cycle[12665] = 1'b1;  addr_rom[12665]='h0000073c;  wr_data_rom[12665]='h0000227d;
    rd_cycle[12666] = 1'b1;  wr_cycle[12666] = 1'b0;  addr_rom[12666]='h000025ec;  wr_data_rom[12666]='h00000000;
    rd_cycle[12667] = 1'b1;  wr_cycle[12667] = 1'b0;  addr_rom[12667]='h000004b4;  wr_data_rom[12667]='h00000000;
    rd_cycle[12668] = 1'b1;  wr_cycle[12668] = 1'b0;  addr_rom[12668]='h000039a0;  wr_data_rom[12668]='h00000000;
    rd_cycle[12669] = 1'b1;  wr_cycle[12669] = 1'b0;  addr_rom[12669]='h00002130;  wr_data_rom[12669]='h00000000;
    rd_cycle[12670] = 1'b0;  wr_cycle[12670] = 1'b1;  addr_rom[12670]='h00000c54;  wr_data_rom[12670]='h00000666;
    rd_cycle[12671] = 1'b0;  wr_cycle[12671] = 1'b1;  addr_rom[12671]='h00000940;  wr_data_rom[12671]='h00001e07;
    rd_cycle[12672] = 1'b1;  wr_cycle[12672] = 1'b0;  addr_rom[12672]='h00002bfc;  wr_data_rom[12672]='h00000000;
    rd_cycle[12673] = 1'b0;  wr_cycle[12673] = 1'b1;  addr_rom[12673]='h000036e4;  wr_data_rom[12673]='h00003ebc;
    rd_cycle[12674] = 1'b0;  wr_cycle[12674] = 1'b1;  addr_rom[12674]='h000032ec;  wr_data_rom[12674]='h000034aa;
    rd_cycle[12675] = 1'b1;  wr_cycle[12675] = 1'b0;  addr_rom[12675]='h00001154;  wr_data_rom[12675]='h00000000;
    rd_cycle[12676] = 1'b0;  wr_cycle[12676] = 1'b1;  addr_rom[12676]='h00003314;  wr_data_rom[12676]='h00000ddd;
    rd_cycle[12677] = 1'b0;  wr_cycle[12677] = 1'b1;  addr_rom[12677]='h000031e4;  wr_data_rom[12677]='h00001051;
    rd_cycle[12678] = 1'b0;  wr_cycle[12678] = 1'b1;  addr_rom[12678]='h00001590;  wr_data_rom[12678]='h00003d06;
    rd_cycle[12679] = 1'b1;  wr_cycle[12679] = 1'b0;  addr_rom[12679]='h000020dc;  wr_data_rom[12679]='h00000000;
    rd_cycle[12680] = 1'b0;  wr_cycle[12680] = 1'b1;  addr_rom[12680]='h00003648;  wr_data_rom[12680]='h00000ff5;
    rd_cycle[12681] = 1'b1;  wr_cycle[12681] = 1'b0;  addr_rom[12681]='h00001704;  wr_data_rom[12681]='h00000000;
    rd_cycle[12682] = 1'b1;  wr_cycle[12682] = 1'b0;  addr_rom[12682]='h00003e90;  wr_data_rom[12682]='h00000000;
    rd_cycle[12683] = 1'b0;  wr_cycle[12683] = 1'b1;  addr_rom[12683]='h0000260c;  wr_data_rom[12683]='h000032ff;
    rd_cycle[12684] = 1'b0;  wr_cycle[12684] = 1'b1;  addr_rom[12684]='h00002df4;  wr_data_rom[12684]='h0000399c;
    rd_cycle[12685] = 1'b1;  wr_cycle[12685] = 1'b0;  addr_rom[12685]='h000006cc;  wr_data_rom[12685]='h00000000;
    rd_cycle[12686] = 1'b0;  wr_cycle[12686] = 1'b1;  addr_rom[12686]='h000008b4;  wr_data_rom[12686]='h000020bd;
    rd_cycle[12687] = 1'b0;  wr_cycle[12687] = 1'b1;  addr_rom[12687]='h00003e00;  wr_data_rom[12687]='h0000021b;
    rd_cycle[12688] = 1'b0;  wr_cycle[12688] = 1'b1;  addr_rom[12688]='h00001de4;  wr_data_rom[12688]='h00001b0d;
    rd_cycle[12689] = 1'b0;  wr_cycle[12689] = 1'b1;  addr_rom[12689]='h00000ac4;  wr_data_rom[12689]='h00003ca1;
    rd_cycle[12690] = 1'b1;  wr_cycle[12690] = 1'b0;  addr_rom[12690]='h00002118;  wr_data_rom[12690]='h00000000;
    rd_cycle[12691] = 1'b1;  wr_cycle[12691] = 1'b0;  addr_rom[12691]='h00000cd4;  wr_data_rom[12691]='h00000000;
    rd_cycle[12692] = 1'b0;  wr_cycle[12692] = 1'b1;  addr_rom[12692]='h00000f30;  wr_data_rom[12692]='h00003fea;
    rd_cycle[12693] = 1'b1;  wr_cycle[12693] = 1'b0;  addr_rom[12693]='h00003a84;  wr_data_rom[12693]='h00000000;
    rd_cycle[12694] = 1'b1;  wr_cycle[12694] = 1'b0;  addr_rom[12694]='h000004f8;  wr_data_rom[12694]='h00000000;
    rd_cycle[12695] = 1'b1;  wr_cycle[12695] = 1'b0;  addr_rom[12695]='h0000090c;  wr_data_rom[12695]='h00000000;
    rd_cycle[12696] = 1'b1;  wr_cycle[12696] = 1'b0;  addr_rom[12696]='h000039b0;  wr_data_rom[12696]='h00000000;
    rd_cycle[12697] = 1'b0;  wr_cycle[12697] = 1'b1;  addr_rom[12697]='h0000131c;  wr_data_rom[12697]='h00001f7d;
    rd_cycle[12698] = 1'b0;  wr_cycle[12698] = 1'b1;  addr_rom[12698]='h00002d8c;  wr_data_rom[12698]='h000018f4;
    rd_cycle[12699] = 1'b0;  wr_cycle[12699] = 1'b1;  addr_rom[12699]='h00000e20;  wr_data_rom[12699]='h00002685;
    rd_cycle[12700] = 1'b1;  wr_cycle[12700] = 1'b0;  addr_rom[12700]='h00000324;  wr_data_rom[12700]='h00000000;
    rd_cycle[12701] = 1'b1;  wr_cycle[12701] = 1'b0;  addr_rom[12701]='h00001a6c;  wr_data_rom[12701]='h00000000;
    rd_cycle[12702] = 1'b0;  wr_cycle[12702] = 1'b1;  addr_rom[12702]='h00002340;  wr_data_rom[12702]='h00000d48;
    rd_cycle[12703] = 1'b1;  wr_cycle[12703] = 1'b0;  addr_rom[12703]='h00003b04;  wr_data_rom[12703]='h00000000;
    rd_cycle[12704] = 1'b1;  wr_cycle[12704] = 1'b0;  addr_rom[12704]='h00000db4;  wr_data_rom[12704]='h00000000;
    rd_cycle[12705] = 1'b1;  wr_cycle[12705] = 1'b0;  addr_rom[12705]='h000016d0;  wr_data_rom[12705]='h00000000;
    rd_cycle[12706] = 1'b1;  wr_cycle[12706] = 1'b0;  addr_rom[12706]='h00001df0;  wr_data_rom[12706]='h00000000;
    rd_cycle[12707] = 1'b0;  wr_cycle[12707] = 1'b1;  addr_rom[12707]='h00003844;  wr_data_rom[12707]='h00000120;
    rd_cycle[12708] = 1'b0;  wr_cycle[12708] = 1'b1;  addr_rom[12708]='h000035b0;  wr_data_rom[12708]='h000003f5;
    rd_cycle[12709] = 1'b0;  wr_cycle[12709] = 1'b1;  addr_rom[12709]='h000021e8;  wr_data_rom[12709]='h00000584;
    rd_cycle[12710] = 1'b0;  wr_cycle[12710] = 1'b1;  addr_rom[12710]='h00002e5c;  wr_data_rom[12710]='h00001a1b;
    rd_cycle[12711] = 1'b1;  wr_cycle[12711] = 1'b0;  addr_rom[12711]='h000002d0;  wr_data_rom[12711]='h00000000;
    rd_cycle[12712] = 1'b1;  wr_cycle[12712] = 1'b0;  addr_rom[12712]='h000020b8;  wr_data_rom[12712]='h00000000;
    rd_cycle[12713] = 1'b1;  wr_cycle[12713] = 1'b0;  addr_rom[12713]='h0000029c;  wr_data_rom[12713]='h00000000;
    rd_cycle[12714] = 1'b0;  wr_cycle[12714] = 1'b1;  addr_rom[12714]='h00000fc4;  wr_data_rom[12714]='h00003817;
    rd_cycle[12715] = 1'b0;  wr_cycle[12715] = 1'b1;  addr_rom[12715]='h00001738;  wr_data_rom[12715]='h00003ac5;
    rd_cycle[12716] = 1'b1;  wr_cycle[12716] = 1'b0;  addr_rom[12716]='h00002fb4;  wr_data_rom[12716]='h00000000;
    rd_cycle[12717] = 1'b1;  wr_cycle[12717] = 1'b0;  addr_rom[12717]='h00002090;  wr_data_rom[12717]='h00000000;
    rd_cycle[12718] = 1'b0;  wr_cycle[12718] = 1'b1;  addr_rom[12718]='h000018b8;  wr_data_rom[12718]='h00002cc7;
    rd_cycle[12719] = 1'b0;  wr_cycle[12719] = 1'b1;  addr_rom[12719]='h00000a7c;  wr_data_rom[12719]='h00003fb6;
    rd_cycle[12720] = 1'b0;  wr_cycle[12720] = 1'b1;  addr_rom[12720]='h00000490;  wr_data_rom[12720]='h00003020;
    rd_cycle[12721] = 1'b0;  wr_cycle[12721] = 1'b1;  addr_rom[12721]='h00002614;  wr_data_rom[12721]='h0000076e;
    rd_cycle[12722] = 1'b0;  wr_cycle[12722] = 1'b1;  addr_rom[12722]='h00003ed0;  wr_data_rom[12722]='h00001eb0;
    rd_cycle[12723] = 1'b1;  wr_cycle[12723] = 1'b0;  addr_rom[12723]='h00001ef8;  wr_data_rom[12723]='h00000000;
    rd_cycle[12724] = 1'b0;  wr_cycle[12724] = 1'b1;  addr_rom[12724]='h0000248c;  wr_data_rom[12724]='h00002b18;
    rd_cycle[12725] = 1'b0;  wr_cycle[12725] = 1'b1;  addr_rom[12725]='h00001198;  wr_data_rom[12725]='h00003f5a;
    rd_cycle[12726] = 1'b1;  wr_cycle[12726] = 1'b0;  addr_rom[12726]='h00000474;  wr_data_rom[12726]='h00000000;
    rd_cycle[12727] = 1'b0;  wr_cycle[12727] = 1'b1;  addr_rom[12727]='h00000eac;  wr_data_rom[12727]='h00000a6f;
    rd_cycle[12728] = 1'b1;  wr_cycle[12728] = 1'b0;  addr_rom[12728]='h0000272c;  wr_data_rom[12728]='h00000000;
    rd_cycle[12729] = 1'b1;  wr_cycle[12729] = 1'b0;  addr_rom[12729]='h0000321c;  wr_data_rom[12729]='h00000000;
    rd_cycle[12730] = 1'b1;  wr_cycle[12730] = 1'b0;  addr_rom[12730]='h00002544;  wr_data_rom[12730]='h00000000;
    rd_cycle[12731] = 1'b1;  wr_cycle[12731] = 1'b0;  addr_rom[12731]='h00003184;  wr_data_rom[12731]='h00000000;
    rd_cycle[12732] = 1'b1;  wr_cycle[12732] = 1'b0;  addr_rom[12732]='h00001aa4;  wr_data_rom[12732]='h00000000;
    rd_cycle[12733] = 1'b0;  wr_cycle[12733] = 1'b1;  addr_rom[12733]='h00003e50;  wr_data_rom[12733]='h00000e46;
    rd_cycle[12734] = 1'b1;  wr_cycle[12734] = 1'b0;  addr_rom[12734]='h00000b90;  wr_data_rom[12734]='h00000000;
    rd_cycle[12735] = 1'b1;  wr_cycle[12735] = 1'b0;  addr_rom[12735]='h00002dd4;  wr_data_rom[12735]='h00000000;
    rd_cycle[12736] = 1'b1;  wr_cycle[12736] = 1'b0;  addr_rom[12736]='h00002fcc;  wr_data_rom[12736]='h00000000;
    rd_cycle[12737] = 1'b1;  wr_cycle[12737] = 1'b0;  addr_rom[12737]='h00001d70;  wr_data_rom[12737]='h00000000;
    rd_cycle[12738] = 1'b0;  wr_cycle[12738] = 1'b1;  addr_rom[12738]='h00003bd4;  wr_data_rom[12738]='h000012a5;
    rd_cycle[12739] = 1'b0;  wr_cycle[12739] = 1'b1;  addr_rom[12739]='h00003464;  wr_data_rom[12739]='h00001abf;
    rd_cycle[12740] = 1'b0;  wr_cycle[12740] = 1'b1;  addr_rom[12740]='h000010e0;  wr_data_rom[12740]='h00003df5;
    rd_cycle[12741] = 1'b0;  wr_cycle[12741] = 1'b1;  addr_rom[12741]='h00002248;  wr_data_rom[12741]='h00002797;
    rd_cycle[12742] = 1'b1;  wr_cycle[12742] = 1'b0;  addr_rom[12742]='h00000158;  wr_data_rom[12742]='h00000000;
    rd_cycle[12743] = 1'b0;  wr_cycle[12743] = 1'b1;  addr_rom[12743]='h00002900;  wr_data_rom[12743]='h00003e59;
    rd_cycle[12744] = 1'b0;  wr_cycle[12744] = 1'b1;  addr_rom[12744]='h00000d64;  wr_data_rom[12744]='h00002426;
    rd_cycle[12745] = 1'b1;  wr_cycle[12745] = 1'b0;  addr_rom[12745]='h000038f0;  wr_data_rom[12745]='h00000000;
    rd_cycle[12746] = 1'b0;  wr_cycle[12746] = 1'b1;  addr_rom[12746]='h00001f50;  wr_data_rom[12746]='h00003060;
    rd_cycle[12747] = 1'b1;  wr_cycle[12747] = 1'b0;  addr_rom[12747]='h0000311c;  wr_data_rom[12747]='h00000000;
    rd_cycle[12748] = 1'b0;  wr_cycle[12748] = 1'b1;  addr_rom[12748]='h00000838;  wr_data_rom[12748]='h00002b8d;
    rd_cycle[12749] = 1'b0;  wr_cycle[12749] = 1'b1;  addr_rom[12749]='h00000840;  wr_data_rom[12749]='h000008ba;
    rd_cycle[12750] = 1'b1;  wr_cycle[12750] = 1'b0;  addr_rom[12750]='h0000061c;  wr_data_rom[12750]='h00000000;
    rd_cycle[12751] = 1'b1;  wr_cycle[12751] = 1'b0;  addr_rom[12751]='h00003a84;  wr_data_rom[12751]='h00000000;
    rd_cycle[12752] = 1'b1;  wr_cycle[12752] = 1'b0;  addr_rom[12752]='h00000f8c;  wr_data_rom[12752]='h00000000;
    rd_cycle[12753] = 1'b0;  wr_cycle[12753] = 1'b1;  addr_rom[12753]='h000017f8;  wr_data_rom[12753]='h0000101b;
    rd_cycle[12754] = 1'b1;  wr_cycle[12754] = 1'b0;  addr_rom[12754]='h00002d04;  wr_data_rom[12754]='h00000000;
    rd_cycle[12755] = 1'b1;  wr_cycle[12755] = 1'b0;  addr_rom[12755]='h00000b78;  wr_data_rom[12755]='h00000000;
    rd_cycle[12756] = 1'b1;  wr_cycle[12756] = 1'b0;  addr_rom[12756]='h000018e8;  wr_data_rom[12756]='h00000000;
    rd_cycle[12757] = 1'b0;  wr_cycle[12757] = 1'b1;  addr_rom[12757]='h0000243c;  wr_data_rom[12757]='h000019a5;
    rd_cycle[12758] = 1'b1;  wr_cycle[12758] = 1'b0;  addr_rom[12758]='h0000121c;  wr_data_rom[12758]='h00000000;
    rd_cycle[12759] = 1'b0;  wr_cycle[12759] = 1'b1;  addr_rom[12759]='h00000bb0;  wr_data_rom[12759]='h000036f8;
    rd_cycle[12760] = 1'b1;  wr_cycle[12760] = 1'b0;  addr_rom[12760]='h000019c0;  wr_data_rom[12760]='h00000000;
    rd_cycle[12761] = 1'b0;  wr_cycle[12761] = 1'b1;  addr_rom[12761]='h00002c78;  wr_data_rom[12761]='h0000074b;
    rd_cycle[12762] = 1'b1;  wr_cycle[12762] = 1'b0;  addr_rom[12762]='h00000538;  wr_data_rom[12762]='h00000000;
    rd_cycle[12763] = 1'b0;  wr_cycle[12763] = 1'b1;  addr_rom[12763]='h00000b44;  wr_data_rom[12763]='h00002314;
    rd_cycle[12764] = 1'b0;  wr_cycle[12764] = 1'b1;  addr_rom[12764]='h00003120;  wr_data_rom[12764]='h000012fe;
    rd_cycle[12765] = 1'b1;  wr_cycle[12765] = 1'b0;  addr_rom[12765]='h00000ad4;  wr_data_rom[12765]='h00000000;
    rd_cycle[12766] = 1'b0;  wr_cycle[12766] = 1'b1;  addr_rom[12766]='h0000050c;  wr_data_rom[12766]='h00000f98;
    rd_cycle[12767] = 1'b1;  wr_cycle[12767] = 1'b0;  addr_rom[12767]='h000007f4;  wr_data_rom[12767]='h00000000;
    rd_cycle[12768] = 1'b0;  wr_cycle[12768] = 1'b1;  addr_rom[12768]='h00003c18;  wr_data_rom[12768]='h0000012a;
    rd_cycle[12769] = 1'b0;  wr_cycle[12769] = 1'b1;  addr_rom[12769]='h00003c44;  wr_data_rom[12769]='h00000bd3;
    rd_cycle[12770] = 1'b0;  wr_cycle[12770] = 1'b1;  addr_rom[12770]='h00001084;  wr_data_rom[12770]='h00003b52;
    rd_cycle[12771] = 1'b0;  wr_cycle[12771] = 1'b1;  addr_rom[12771]='h0000202c;  wr_data_rom[12771]='h00002494;
    rd_cycle[12772] = 1'b0;  wr_cycle[12772] = 1'b1;  addr_rom[12772]='h00001f24;  wr_data_rom[12772]='h00002b28;
    rd_cycle[12773] = 1'b0;  wr_cycle[12773] = 1'b1;  addr_rom[12773]='h000020d0;  wr_data_rom[12773]='h00002993;
    rd_cycle[12774] = 1'b0;  wr_cycle[12774] = 1'b1;  addr_rom[12774]='h00002920;  wr_data_rom[12774]='h00002381;
    rd_cycle[12775] = 1'b0;  wr_cycle[12775] = 1'b1;  addr_rom[12775]='h000020fc;  wr_data_rom[12775]='h00002d8a;
    rd_cycle[12776] = 1'b1;  wr_cycle[12776] = 1'b0;  addr_rom[12776]='h00002988;  wr_data_rom[12776]='h00000000;
    rd_cycle[12777] = 1'b0;  wr_cycle[12777] = 1'b1;  addr_rom[12777]='h00001614;  wr_data_rom[12777]='h00000e43;
    rd_cycle[12778] = 1'b0;  wr_cycle[12778] = 1'b1;  addr_rom[12778]='h00000fc4;  wr_data_rom[12778]='h00003fd9;
    rd_cycle[12779] = 1'b0;  wr_cycle[12779] = 1'b1;  addr_rom[12779]='h00000e2c;  wr_data_rom[12779]='h000021cd;
    rd_cycle[12780] = 1'b0;  wr_cycle[12780] = 1'b1;  addr_rom[12780]='h0000357c;  wr_data_rom[12780]='h00002128;
    rd_cycle[12781] = 1'b0;  wr_cycle[12781] = 1'b1;  addr_rom[12781]='h000017f8;  wr_data_rom[12781]='h00001cc9;
    rd_cycle[12782] = 1'b1;  wr_cycle[12782] = 1'b0;  addr_rom[12782]='h00000ee0;  wr_data_rom[12782]='h00000000;
    rd_cycle[12783] = 1'b1;  wr_cycle[12783] = 1'b0;  addr_rom[12783]='h00002be4;  wr_data_rom[12783]='h00000000;
    rd_cycle[12784] = 1'b0;  wr_cycle[12784] = 1'b1;  addr_rom[12784]='h0000135c;  wr_data_rom[12784]='h00000d84;
    rd_cycle[12785] = 1'b1;  wr_cycle[12785] = 1'b0;  addr_rom[12785]='h0000234c;  wr_data_rom[12785]='h00000000;
    rd_cycle[12786] = 1'b0;  wr_cycle[12786] = 1'b1;  addr_rom[12786]='h00001b74;  wr_data_rom[12786]='h00001288;
    rd_cycle[12787] = 1'b1;  wr_cycle[12787] = 1'b0;  addr_rom[12787]='h000023f0;  wr_data_rom[12787]='h00000000;
    rd_cycle[12788] = 1'b0;  wr_cycle[12788] = 1'b1;  addr_rom[12788]='h00002e48;  wr_data_rom[12788]='h00001513;
    rd_cycle[12789] = 1'b0;  wr_cycle[12789] = 1'b1;  addr_rom[12789]='h000028f0;  wr_data_rom[12789]='h0000262c;
    rd_cycle[12790] = 1'b0;  wr_cycle[12790] = 1'b1;  addr_rom[12790]='h00001f48;  wr_data_rom[12790]='h00003f74;
    rd_cycle[12791] = 1'b0;  wr_cycle[12791] = 1'b1;  addr_rom[12791]='h000021b4;  wr_data_rom[12791]='h000031ad;
    rd_cycle[12792] = 1'b1;  wr_cycle[12792] = 1'b0;  addr_rom[12792]='h00000fec;  wr_data_rom[12792]='h00000000;
    rd_cycle[12793] = 1'b0;  wr_cycle[12793] = 1'b1;  addr_rom[12793]='h00003ed4;  wr_data_rom[12793]='h0000380e;
    rd_cycle[12794] = 1'b0;  wr_cycle[12794] = 1'b1;  addr_rom[12794]='h00000d68;  wr_data_rom[12794]='h00000971;
    rd_cycle[12795] = 1'b1;  wr_cycle[12795] = 1'b0;  addr_rom[12795]='h00003504;  wr_data_rom[12795]='h00000000;
    rd_cycle[12796] = 1'b0;  wr_cycle[12796] = 1'b1;  addr_rom[12796]='h0000143c;  wr_data_rom[12796]='h00003f9d;
    rd_cycle[12797] = 1'b0;  wr_cycle[12797] = 1'b1;  addr_rom[12797]='h00002030;  wr_data_rom[12797]='h00003f02;
    rd_cycle[12798] = 1'b0;  wr_cycle[12798] = 1'b1;  addr_rom[12798]='h00002b40;  wr_data_rom[12798]='h00002b29;
    rd_cycle[12799] = 1'b0;  wr_cycle[12799] = 1'b1;  addr_rom[12799]='h000033f8;  wr_data_rom[12799]='h0000094c;
    rd_cycle[12800] = 1'b1;  wr_cycle[12800] = 1'b0;  addr_rom[12800]='h00002050;  wr_data_rom[12800]='h00000000;
    rd_cycle[12801] = 1'b0;  wr_cycle[12801] = 1'b1;  addr_rom[12801]='h00003a80;  wr_data_rom[12801]='h00002607;
    rd_cycle[12802] = 1'b1;  wr_cycle[12802] = 1'b0;  addr_rom[12802]='h00003674;  wr_data_rom[12802]='h00000000;
    rd_cycle[12803] = 1'b0;  wr_cycle[12803] = 1'b1;  addr_rom[12803]='h00002eb0;  wr_data_rom[12803]='h000006b8;
    rd_cycle[12804] = 1'b1;  wr_cycle[12804] = 1'b0;  addr_rom[12804]='h000035b4;  wr_data_rom[12804]='h00000000;
    rd_cycle[12805] = 1'b0;  wr_cycle[12805] = 1'b1;  addr_rom[12805]='h00000ba8;  wr_data_rom[12805]='h0000273c;
    rd_cycle[12806] = 1'b0;  wr_cycle[12806] = 1'b1;  addr_rom[12806]='h00003f74;  wr_data_rom[12806]='h000001a6;
    rd_cycle[12807] = 1'b1;  wr_cycle[12807] = 1'b0;  addr_rom[12807]='h00002a50;  wr_data_rom[12807]='h00000000;
    rd_cycle[12808] = 1'b1;  wr_cycle[12808] = 1'b0;  addr_rom[12808]='h0000144c;  wr_data_rom[12808]='h00000000;
    rd_cycle[12809] = 1'b0;  wr_cycle[12809] = 1'b1;  addr_rom[12809]='h00003550;  wr_data_rom[12809]='h00003df5;
    rd_cycle[12810] = 1'b1;  wr_cycle[12810] = 1'b0;  addr_rom[12810]='h00001dfc;  wr_data_rom[12810]='h00000000;
    rd_cycle[12811] = 1'b1;  wr_cycle[12811] = 1'b0;  addr_rom[12811]='h000008b4;  wr_data_rom[12811]='h00000000;
    rd_cycle[12812] = 1'b1;  wr_cycle[12812] = 1'b0;  addr_rom[12812]='h0000338c;  wr_data_rom[12812]='h00000000;
    rd_cycle[12813] = 1'b0;  wr_cycle[12813] = 1'b1;  addr_rom[12813]='h00002ac8;  wr_data_rom[12813]='h00000809;
    rd_cycle[12814] = 1'b0;  wr_cycle[12814] = 1'b1;  addr_rom[12814]='h00000e80;  wr_data_rom[12814]='h0000348c;
    rd_cycle[12815] = 1'b0;  wr_cycle[12815] = 1'b1;  addr_rom[12815]='h000017d8;  wr_data_rom[12815]='h00000988;
    rd_cycle[12816] = 1'b0;  wr_cycle[12816] = 1'b1;  addr_rom[12816]='h00003bb8;  wr_data_rom[12816]='h000030b1;
    rd_cycle[12817] = 1'b1;  wr_cycle[12817] = 1'b0;  addr_rom[12817]='h00000678;  wr_data_rom[12817]='h00000000;
    rd_cycle[12818] = 1'b1;  wr_cycle[12818] = 1'b0;  addr_rom[12818]='h00002858;  wr_data_rom[12818]='h00000000;
    rd_cycle[12819] = 1'b0;  wr_cycle[12819] = 1'b1;  addr_rom[12819]='h00000cb4;  wr_data_rom[12819]='h00003c28;
    rd_cycle[12820] = 1'b0;  wr_cycle[12820] = 1'b1;  addr_rom[12820]='h000004fc;  wr_data_rom[12820]='h00001e0e;
    rd_cycle[12821] = 1'b1;  wr_cycle[12821] = 1'b0;  addr_rom[12821]='h00000f60;  wr_data_rom[12821]='h00000000;
    rd_cycle[12822] = 1'b1;  wr_cycle[12822] = 1'b0;  addr_rom[12822]='h0000188c;  wr_data_rom[12822]='h00000000;
    rd_cycle[12823] = 1'b0;  wr_cycle[12823] = 1'b1;  addr_rom[12823]='h000028b4;  wr_data_rom[12823]='h00000e95;
    rd_cycle[12824] = 1'b0;  wr_cycle[12824] = 1'b1;  addr_rom[12824]='h00000260;  wr_data_rom[12824]='h0000028b;
    rd_cycle[12825] = 1'b0;  wr_cycle[12825] = 1'b1;  addr_rom[12825]='h00003e14;  wr_data_rom[12825]='h00002594;
    rd_cycle[12826] = 1'b1;  wr_cycle[12826] = 1'b0;  addr_rom[12826]='h00002098;  wr_data_rom[12826]='h00000000;
    rd_cycle[12827] = 1'b1;  wr_cycle[12827] = 1'b0;  addr_rom[12827]='h00003054;  wr_data_rom[12827]='h00000000;
    rd_cycle[12828] = 1'b0;  wr_cycle[12828] = 1'b1;  addr_rom[12828]='h00003e6c;  wr_data_rom[12828]='h00000bcc;
    rd_cycle[12829] = 1'b0;  wr_cycle[12829] = 1'b1;  addr_rom[12829]='h00002bb0;  wr_data_rom[12829]='h00003b16;
    rd_cycle[12830] = 1'b0;  wr_cycle[12830] = 1'b1;  addr_rom[12830]='h0000123c;  wr_data_rom[12830]='h00001dc7;
    rd_cycle[12831] = 1'b1;  wr_cycle[12831] = 1'b0;  addr_rom[12831]='h00002514;  wr_data_rom[12831]='h00000000;
    rd_cycle[12832] = 1'b1;  wr_cycle[12832] = 1'b0;  addr_rom[12832]='h00000d10;  wr_data_rom[12832]='h00000000;
    rd_cycle[12833] = 1'b0;  wr_cycle[12833] = 1'b1;  addr_rom[12833]='h00003d04;  wr_data_rom[12833]='h000016c9;
    rd_cycle[12834] = 1'b1;  wr_cycle[12834] = 1'b0;  addr_rom[12834]='h0000266c;  wr_data_rom[12834]='h00000000;
    rd_cycle[12835] = 1'b1;  wr_cycle[12835] = 1'b0;  addr_rom[12835]='h000007f4;  wr_data_rom[12835]='h00000000;
    rd_cycle[12836] = 1'b1;  wr_cycle[12836] = 1'b0;  addr_rom[12836]='h00000530;  wr_data_rom[12836]='h00000000;
    rd_cycle[12837] = 1'b0;  wr_cycle[12837] = 1'b1;  addr_rom[12837]='h00002f30;  wr_data_rom[12837]='h00002a17;
    rd_cycle[12838] = 1'b0;  wr_cycle[12838] = 1'b1;  addr_rom[12838]='h00001df0;  wr_data_rom[12838]='h00003a19;
    rd_cycle[12839] = 1'b1;  wr_cycle[12839] = 1'b0;  addr_rom[12839]='h000029c0;  wr_data_rom[12839]='h00000000;
    rd_cycle[12840] = 1'b1;  wr_cycle[12840] = 1'b0;  addr_rom[12840]='h00003cc4;  wr_data_rom[12840]='h00000000;
    rd_cycle[12841] = 1'b0;  wr_cycle[12841] = 1'b1;  addr_rom[12841]='h00003d2c;  wr_data_rom[12841]='h00002b97;
    rd_cycle[12842] = 1'b1;  wr_cycle[12842] = 1'b0;  addr_rom[12842]='h0000340c;  wr_data_rom[12842]='h00000000;
    rd_cycle[12843] = 1'b1;  wr_cycle[12843] = 1'b0;  addr_rom[12843]='h00001c5c;  wr_data_rom[12843]='h00000000;
    rd_cycle[12844] = 1'b1;  wr_cycle[12844] = 1'b0;  addr_rom[12844]='h00002968;  wr_data_rom[12844]='h00000000;
    rd_cycle[12845] = 1'b1;  wr_cycle[12845] = 1'b0;  addr_rom[12845]='h00000618;  wr_data_rom[12845]='h00000000;
    rd_cycle[12846] = 1'b1;  wr_cycle[12846] = 1'b0;  addr_rom[12846]='h00001268;  wr_data_rom[12846]='h00000000;
    rd_cycle[12847] = 1'b0;  wr_cycle[12847] = 1'b1;  addr_rom[12847]='h00003e80;  wr_data_rom[12847]='h00001712;
    rd_cycle[12848] = 1'b1;  wr_cycle[12848] = 1'b0;  addr_rom[12848]='h000014ec;  wr_data_rom[12848]='h00000000;
    rd_cycle[12849] = 1'b1;  wr_cycle[12849] = 1'b0;  addr_rom[12849]='h0000242c;  wr_data_rom[12849]='h00000000;
    rd_cycle[12850] = 1'b1;  wr_cycle[12850] = 1'b0;  addr_rom[12850]='h000027e0;  wr_data_rom[12850]='h00000000;
    rd_cycle[12851] = 1'b0;  wr_cycle[12851] = 1'b1;  addr_rom[12851]='h00002da8;  wr_data_rom[12851]='h000015b6;
    rd_cycle[12852] = 1'b1;  wr_cycle[12852] = 1'b0;  addr_rom[12852]='h000000c0;  wr_data_rom[12852]='h00000000;
    rd_cycle[12853] = 1'b1;  wr_cycle[12853] = 1'b0;  addr_rom[12853]='h0000371c;  wr_data_rom[12853]='h00000000;
    rd_cycle[12854] = 1'b0;  wr_cycle[12854] = 1'b1;  addr_rom[12854]='h00000fd4;  wr_data_rom[12854]='h000025f6;
    rd_cycle[12855] = 1'b0;  wr_cycle[12855] = 1'b1;  addr_rom[12855]='h00003184;  wr_data_rom[12855]='h000026ff;
    rd_cycle[12856] = 1'b1;  wr_cycle[12856] = 1'b0;  addr_rom[12856]='h000015e0;  wr_data_rom[12856]='h00000000;
    rd_cycle[12857] = 1'b1;  wr_cycle[12857] = 1'b0;  addr_rom[12857]='h00000c8c;  wr_data_rom[12857]='h00000000;
    rd_cycle[12858] = 1'b1;  wr_cycle[12858] = 1'b0;  addr_rom[12858]='h00001a7c;  wr_data_rom[12858]='h00000000;
    rd_cycle[12859] = 1'b0;  wr_cycle[12859] = 1'b1;  addr_rom[12859]='h00003130;  wr_data_rom[12859]='h00002a48;
    rd_cycle[12860] = 1'b0;  wr_cycle[12860] = 1'b1;  addr_rom[12860]='h00001810;  wr_data_rom[12860]='h00000c3f;
    rd_cycle[12861] = 1'b1;  wr_cycle[12861] = 1'b0;  addr_rom[12861]='h00000994;  wr_data_rom[12861]='h00000000;
    rd_cycle[12862] = 1'b0;  wr_cycle[12862] = 1'b1;  addr_rom[12862]='h00000c98;  wr_data_rom[12862]='h000022b3;
    rd_cycle[12863] = 1'b0;  wr_cycle[12863] = 1'b1;  addr_rom[12863]='h00000770;  wr_data_rom[12863]='h000032ad;
    rd_cycle[12864] = 1'b1;  wr_cycle[12864] = 1'b0;  addr_rom[12864]='h00000900;  wr_data_rom[12864]='h00000000;
    rd_cycle[12865] = 1'b0;  wr_cycle[12865] = 1'b1;  addr_rom[12865]='h00001058;  wr_data_rom[12865]='h0000203e;
    rd_cycle[12866] = 1'b0;  wr_cycle[12866] = 1'b1;  addr_rom[12866]='h00001388;  wr_data_rom[12866]='h00001581;
    rd_cycle[12867] = 1'b0;  wr_cycle[12867] = 1'b1;  addr_rom[12867]='h00000770;  wr_data_rom[12867]='h00000c01;
    rd_cycle[12868] = 1'b1;  wr_cycle[12868] = 1'b0;  addr_rom[12868]='h000020a0;  wr_data_rom[12868]='h00000000;
    rd_cycle[12869] = 1'b1;  wr_cycle[12869] = 1'b0;  addr_rom[12869]='h00000cc0;  wr_data_rom[12869]='h00000000;
    rd_cycle[12870] = 1'b0;  wr_cycle[12870] = 1'b1;  addr_rom[12870]='h00000a70;  wr_data_rom[12870]='h00001030;
    rd_cycle[12871] = 1'b1;  wr_cycle[12871] = 1'b0;  addr_rom[12871]='h00000734;  wr_data_rom[12871]='h00000000;
    rd_cycle[12872] = 1'b0;  wr_cycle[12872] = 1'b1;  addr_rom[12872]='h000038b0;  wr_data_rom[12872]='h00002769;
    rd_cycle[12873] = 1'b0;  wr_cycle[12873] = 1'b1;  addr_rom[12873]='h00001ff8;  wr_data_rom[12873]='h00000939;
    rd_cycle[12874] = 1'b0;  wr_cycle[12874] = 1'b1;  addr_rom[12874]='h00002d2c;  wr_data_rom[12874]='h00000c9e;
    rd_cycle[12875] = 1'b1;  wr_cycle[12875] = 1'b0;  addr_rom[12875]='h00000a54;  wr_data_rom[12875]='h00000000;
    rd_cycle[12876] = 1'b1;  wr_cycle[12876] = 1'b0;  addr_rom[12876]='h00000478;  wr_data_rom[12876]='h00000000;
    rd_cycle[12877] = 1'b1;  wr_cycle[12877] = 1'b0;  addr_rom[12877]='h00001258;  wr_data_rom[12877]='h00000000;
    rd_cycle[12878] = 1'b1;  wr_cycle[12878] = 1'b0;  addr_rom[12878]='h00002c10;  wr_data_rom[12878]='h00000000;
    rd_cycle[12879] = 1'b0;  wr_cycle[12879] = 1'b1;  addr_rom[12879]='h000030a0;  wr_data_rom[12879]='h00001789;
    rd_cycle[12880] = 1'b1;  wr_cycle[12880] = 1'b0;  addr_rom[12880]='h00001154;  wr_data_rom[12880]='h00000000;
    rd_cycle[12881] = 1'b0;  wr_cycle[12881] = 1'b1;  addr_rom[12881]='h000021f8;  wr_data_rom[12881]='h00001f6f;
    rd_cycle[12882] = 1'b0;  wr_cycle[12882] = 1'b1;  addr_rom[12882]='h000004e8;  wr_data_rom[12882]='h000027c3;
    rd_cycle[12883] = 1'b1;  wr_cycle[12883] = 1'b0;  addr_rom[12883]='h00002550;  wr_data_rom[12883]='h00000000;
    rd_cycle[12884] = 1'b1;  wr_cycle[12884] = 1'b0;  addr_rom[12884]='h00001f78;  wr_data_rom[12884]='h00000000;
    rd_cycle[12885] = 1'b0;  wr_cycle[12885] = 1'b1;  addr_rom[12885]='h00000c54;  wr_data_rom[12885]='h000017cb;
    rd_cycle[12886] = 1'b0;  wr_cycle[12886] = 1'b1;  addr_rom[12886]='h00000a1c;  wr_data_rom[12886]='h0000120c;
    rd_cycle[12887] = 1'b0;  wr_cycle[12887] = 1'b1;  addr_rom[12887]='h00001fa0;  wr_data_rom[12887]='h000010d5;
    rd_cycle[12888] = 1'b1;  wr_cycle[12888] = 1'b0;  addr_rom[12888]='h00001fc8;  wr_data_rom[12888]='h00000000;
    rd_cycle[12889] = 1'b1;  wr_cycle[12889] = 1'b0;  addr_rom[12889]='h00002614;  wr_data_rom[12889]='h00000000;
    rd_cycle[12890] = 1'b0;  wr_cycle[12890] = 1'b1;  addr_rom[12890]='h00002368;  wr_data_rom[12890]='h0000372d;
    rd_cycle[12891] = 1'b1;  wr_cycle[12891] = 1'b0;  addr_rom[12891]='h00002cd4;  wr_data_rom[12891]='h00000000;
    rd_cycle[12892] = 1'b0;  wr_cycle[12892] = 1'b1;  addr_rom[12892]='h00000398;  wr_data_rom[12892]='h000014a4;
    rd_cycle[12893] = 1'b0;  wr_cycle[12893] = 1'b1;  addr_rom[12893]='h00001578;  wr_data_rom[12893]='h0000255e;
    rd_cycle[12894] = 1'b0;  wr_cycle[12894] = 1'b1;  addr_rom[12894]='h00002a5c;  wr_data_rom[12894]='h00003a50;
    rd_cycle[12895] = 1'b0;  wr_cycle[12895] = 1'b1;  addr_rom[12895]='h0000110c;  wr_data_rom[12895]='h0000248a;
    rd_cycle[12896] = 1'b1;  wr_cycle[12896] = 1'b0;  addr_rom[12896]='h00002604;  wr_data_rom[12896]='h00000000;
    rd_cycle[12897] = 1'b1;  wr_cycle[12897] = 1'b0;  addr_rom[12897]='h0000392c;  wr_data_rom[12897]='h00000000;
    rd_cycle[12898] = 1'b0;  wr_cycle[12898] = 1'b1;  addr_rom[12898]='h00002388;  wr_data_rom[12898]='h000023f7;
    rd_cycle[12899] = 1'b0;  wr_cycle[12899] = 1'b1;  addr_rom[12899]='h00001334;  wr_data_rom[12899]='h000017df;
    rd_cycle[12900] = 1'b0;  wr_cycle[12900] = 1'b1;  addr_rom[12900]='h00000338;  wr_data_rom[12900]='h000010d4;
    rd_cycle[12901] = 1'b1;  wr_cycle[12901] = 1'b0;  addr_rom[12901]='h0000388c;  wr_data_rom[12901]='h00000000;
    rd_cycle[12902] = 1'b0;  wr_cycle[12902] = 1'b1;  addr_rom[12902]='h000034cc;  wr_data_rom[12902]='h00001b0e;
    rd_cycle[12903] = 1'b1;  wr_cycle[12903] = 1'b0;  addr_rom[12903]='h0000130c;  wr_data_rom[12903]='h00000000;
    rd_cycle[12904] = 1'b0;  wr_cycle[12904] = 1'b1;  addr_rom[12904]='h00000428;  wr_data_rom[12904]='h00000769;
    rd_cycle[12905] = 1'b0;  wr_cycle[12905] = 1'b1;  addr_rom[12905]='h00000e4c;  wr_data_rom[12905]='h000033ac;
    rd_cycle[12906] = 1'b0;  wr_cycle[12906] = 1'b1;  addr_rom[12906]='h00001c14;  wr_data_rom[12906]='h00000e26;
    rd_cycle[12907] = 1'b0;  wr_cycle[12907] = 1'b1;  addr_rom[12907]='h00001770;  wr_data_rom[12907]='h00003d32;
    rd_cycle[12908] = 1'b0;  wr_cycle[12908] = 1'b1;  addr_rom[12908]='h000006e0;  wr_data_rom[12908]='h0000137e;
    rd_cycle[12909] = 1'b1;  wr_cycle[12909] = 1'b0;  addr_rom[12909]='h00002590;  wr_data_rom[12909]='h00000000;
    rd_cycle[12910] = 1'b1;  wr_cycle[12910] = 1'b0;  addr_rom[12910]='h00002a84;  wr_data_rom[12910]='h00000000;
    rd_cycle[12911] = 1'b0;  wr_cycle[12911] = 1'b1;  addr_rom[12911]='h00002e04;  wr_data_rom[12911]='h00003d6d;
    rd_cycle[12912] = 1'b0;  wr_cycle[12912] = 1'b1;  addr_rom[12912]='h000039d0;  wr_data_rom[12912]='h00001fe7;
    rd_cycle[12913] = 1'b1;  wr_cycle[12913] = 1'b0;  addr_rom[12913]='h0000313c;  wr_data_rom[12913]='h00000000;
    rd_cycle[12914] = 1'b1;  wr_cycle[12914] = 1'b0;  addr_rom[12914]='h000031b0;  wr_data_rom[12914]='h00000000;
    rd_cycle[12915] = 1'b0;  wr_cycle[12915] = 1'b1;  addr_rom[12915]='h00002a20;  wr_data_rom[12915]='h00000f39;
    rd_cycle[12916] = 1'b1;  wr_cycle[12916] = 1'b0;  addr_rom[12916]='h00002424;  wr_data_rom[12916]='h00000000;
    rd_cycle[12917] = 1'b0;  wr_cycle[12917] = 1'b1;  addr_rom[12917]='h00003960;  wr_data_rom[12917]='h000028be;
    rd_cycle[12918] = 1'b0;  wr_cycle[12918] = 1'b1;  addr_rom[12918]='h00002904;  wr_data_rom[12918]='h000036b2;
    rd_cycle[12919] = 1'b0;  wr_cycle[12919] = 1'b1;  addr_rom[12919]='h00002c30;  wr_data_rom[12919]='h0000008e;
    rd_cycle[12920] = 1'b0;  wr_cycle[12920] = 1'b1;  addr_rom[12920]='h0000115c;  wr_data_rom[12920]='h00001fbf;
    rd_cycle[12921] = 1'b0;  wr_cycle[12921] = 1'b1;  addr_rom[12921]='h00002968;  wr_data_rom[12921]='h0000310e;
    rd_cycle[12922] = 1'b1;  wr_cycle[12922] = 1'b0;  addr_rom[12922]='h000036cc;  wr_data_rom[12922]='h00000000;
    rd_cycle[12923] = 1'b1;  wr_cycle[12923] = 1'b0;  addr_rom[12923]='h00000918;  wr_data_rom[12923]='h00000000;
    rd_cycle[12924] = 1'b1;  wr_cycle[12924] = 1'b0;  addr_rom[12924]='h000018dc;  wr_data_rom[12924]='h00000000;
    rd_cycle[12925] = 1'b0;  wr_cycle[12925] = 1'b1;  addr_rom[12925]='h00003040;  wr_data_rom[12925]='h0000156a;
    rd_cycle[12926] = 1'b0;  wr_cycle[12926] = 1'b1;  addr_rom[12926]='h0000015c;  wr_data_rom[12926]='h00003b4e;
    rd_cycle[12927] = 1'b1;  wr_cycle[12927] = 1'b0;  addr_rom[12927]='h00003188;  wr_data_rom[12927]='h00000000;
    rd_cycle[12928] = 1'b1;  wr_cycle[12928] = 1'b0;  addr_rom[12928]='h00002a2c;  wr_data_rom[12928]='h00000000;
    rd_cycle[12929] = 1'b1;  wr_cycle[12929] = 1'b0;  addr_rom[12929]='h00002d54;  wr_data_rom[12929]='h00000000;
    rd_cycle[12930] = 1'b1;  wr_cycle[12930] = 1'b0;  addr_rom[12930]='h00002fcc;  wr_data_rom[12930]='h00000000;
    rd_cycle[12931] = 1'b1;  wr_cycle[12931] = 1'b0;  addr_rom[12931]='h00001d10;  wr_data_rom[12931]='h00000000;
    rd_cycle[12932] = 1'b0;  wr_cycle[12932] = 1'b1;  addr_rom[12932]='h00003d7c;  wr_data_rom[12932]='h00003995;
    rd_cycle[12933] = 1'b0;  wr_cycle[12933] = 1'b1;  addr_rom[12933]='h00003f18;  wr_data_rom[12933]='h00002913;
    rd_cycle[12934] = 1'b0;  wr_cycle[12934] = 1'b1;  addr_rom[12934]='h00003378;  wr_data_rom[12934]='h00001a0a;
    rd_cycle[12935] = 1'b0;  wr_cycle[12935] = 1'b1;  addr_rom[12935]='h00000ef0;  wr_data_rom[12935]='h00001eec;
    rd_cycle[12936] = 1'b0;  wr_cycle[12936] = 1'b1;  addr_rom[12936]='h00000b04;  wr_data_rom[12936]='h00003ebf;
    rd_cycle[12937] = 1'b1;  wr_cycle[12937] = 1'b0;  addr_rom[12937]='h00000604;  wr_data_rom[12937]='h00000000;
    rd_cycle[12938] = 1'b0;  wr_cycle[12938] = 1'b1;  addr_rom[12938]='h000036f4;  wr_data_rom[12938]='h0000080f;
    rd_cycle[12939] = 1'b0;  wr_cycle[12939] = 1'b1;  addr_rom[12939]='h00003f60;  wr_data_rom[12939]='h00003904;
    rd_cycle[12940] = 1'b0;  wr_cycle[12940] = 1'b1;  addr_rom[12940]='h00003a1c;  wr_data_rom[12940]='h000029b7;
    rd_cycle[12941] = 1'b1;  wr_cycle[12941] = 1'b0;  addr_rom[12941]='h00002a5c;  wr_data_rom[12941]='h00000000;
    rd_cycle[12942] = 1'b0;  wr_cycle[12942] = 1'b1;  addr_rom[12942]='h0000230c;  wr_data_rom[12942]='h000001dd;
    rd_cycle[12943] = 1'b1;  wr_cycle[12943] = 1'b0;  addr_rom[12943]='h00003314;  wr_data_rom[12943]='h00000000;
    rd_cycle[12944] = 1'b0;  wr_cycle[12944] = 1'b1;  addr_rom[12944]='h00001ee4;  wr_data_rom[12944]='h0000032f;
    rd_cycle[12945] = 1'b1;  wr_cycle[12945] = 1'b0;  addr_rom[12945]='h000011c8;  wr_data_rom[12945]='h00000000;
    rd_cycle[12946] = 1'b1;  wr_cycle[12946] = 1'b0;  addr_rom[12946]='h00003fa8;  wr_data_rom[12946]='h00000000;
    rd_cycle[12947] = 1'b1;  wr_cycle[12947] = 1'b0;  addr_rom[12947]='h000025f8;  wr_data_rom[12947]='h00000000;
    rd_cycle[12948] = 1'b1;  wr_cycle[12948] = 1'b0;  addr_rom[12948]='h000036a8;  wr_data_rom[12948]='h00000000;
    rd_cycle[12949] = 1'b1;  wr_cycle[12949] = 1'b0;  addr_rom[12949]='h000001cc;  wr_data_rom[12949]='h00000000;
    rd_cycle[12950] = 1'b1;  wr_cycle[12950] = 1'b0;  addr_rom[12950]='h00001cb8;  wr_data_rom[12950]='h00000000;
    rd_cycle[12951] = 1'b1;  wr_cycle[12951] = 1'b0;  addr_rom[12951]='h00003394;  wr_data_rom[12951]='h00000000;
    rd_cycle[12952] = 1'b1;  wr_cycle[12952] = 1'b0;  addr_rom[12952]='h00001604;  wr_data_rom[12952]='h00000000;
    rd_cycle[12953] = 1'b0;  wr_cycle[12953] = 1'b1;  addr_rom[12953]='h000009e4;  wr_data_rom[12953]='h000027ea;
    rd_cycle[12954] = 1'b1;  wr_cycle[12954] = 1'b0;  addr_rom[12954]='h00002008;  wr_data_rom[12954]='h00000000;
    rd_cycle[12955] = 1'b1;  wr_cycle[12955] = 1'b0;  addr_rom[12955]='h000032dc;  wr_data_rom[12955]='h00000000;
    rd_cycle[12956] = 1'b1;  wr_cycle[12956] = 1'b0;  addr_rom[12956]='h00003d2c;  wr_data_rom[12956]='h00000000;
    rd_cycle[12957] = 1'b0;  wr_cycle[12957] = 1'b1;  addr_rom[12957]='h000037ac;  wr_data_rom[12957]='h000021c4;
    rd_cycle[12958] = 1'b1;  wr_cycle[12958] = 1'b0;  addr_rom[12958]='h00000598;  wr_data_rom[12958]='h00000000;
    rd_cycle[12959] = 1'b1;  wr_cycle[12959] = 1'b0;  addr_rom[12959]='h00003968;  wr_data_rom[12959]='h00000000;
    rd_cycle[12960] = 1'b0;  wr_cycle[12960] = 1'b1;  addr_rom[12960]='h000011e0;  wr_data_rom[12960]='h00001709;
    rd_cycle[12961] = 1'b0;  wr_cycle[12961] = 1'b1;  addr_rom[12961]='h000023f4;  wr_data_rom[12961]='h00002d32;
    rd_cycle[12962] = 1'b0;  wr_cycle[12962] = 1'b1;  addr_rom[12962]='h00000b00;  wr_data_rom[12962]='h00002446;
    rd_cycle[12963] = 1'b1;  wr_cycle[12963] = 1'b0;  addr_rom[12963]='h00002cb0;  wr_data_rom[12963]='h00000000;
    rd_cycle[12964] = 1'b0;  wr_cycle[12964] = 1'b1;  addr_rom[12964]='h00003a3c;  wr_data_rom[12964]='h00000394;
    rd_cycle[12965] = 1'b0;  wr_cycle[12965] = 1'b1;  addr_rom[12965]='h00000844;  wr_data_rom[12965]='h00001f3e;
    rd_cycle[12966] = 1'b1;  wr_cycle[12966] = 1'b0;  addr_rom[12966]='h00001ee0;  wr_data_rom[12966]='h00000000;
    rd_cycle[12967] = 1'b1;  wr_cycle[12967] = 1'b0;  addr_rom[12967]='h00003e34;  wr_data_rom[12967]='h00000000;
    rd_cycle[12968] = 1'b0;  wr_cycle[12968] = 1'b1;  addr_rom[12968]='h000011c0;  wr_data_rom[12968]='h00002366;
    rd_cycle[12969] = 1'b1;  wr_cycle[12969] = 1'b0;  addr_rom[12969]='h00002198;  wr_data_rom[12969]='h00000000;
    rd_cycle[12970] = 1'b1;  wr_cycle[12970] = 1'b0;  addr_rom[12970]='h00003aac;  wr_data_rom[12970]='h00000000;
    rd_cycle[12971] = 1'b0;  wr_cycle[12971] = 1'b1;  addr_rom[12971]='h00001b6c;  wr_data_rom[12971]='h00000085;
    rd_cycle[12972] = 1'b0;  wr_cycle[12972] = 1'b1;  addr_rom[12972]='h000000ec;  wr_data_rom[12972]='h0000130e;
    rd_cycle[12973] = 1'b1;  wr_cycle[12973] = 1'b0;  addr_rom[12973]='h00001e1c;  wr_data_rom[12973]='h00000000;
    rd_cycle[12974] = 1'b0;  wr_cycle[12974] = 1'b1;  addr_rom[12974]='h00003140;  wr_data_rom[12974]='h00000a56;
    rd_cycle[12975] = 1'b0;  wr_cycle[12975] = 1'b1;  addr_rom[12975]='h0000174c;  wr_data_rom[12975]='h000006b1;
    rd_cycle[12976] = 1'b0;  wr_cycle[12976] = 1'b1;  addr_rom[12976]='h00003440;  wr_data_rom[12976]='h00002cde;
    rd_cycle[12977] = 1'b1;  wr_cycle[12977] = 1'b0;  addr_rom[12977]='h00003534;  wr_data_rom[12977]='h00000000;
    rd_cycle[12978] = 1'b0;  wr_cycle[12978] = 1'b1;  addr_rom[12978]='h000030f4;  wr_data_rom[12978]='h00002b5d;
    rd_cycle[12979] = 1'b1;  wr_cycle[12979] = 1'b0;  addr_rom[12979]='h00001e20;  wr_data_rom[12979]='h00000000;
    rd_cycle[12980] = 1'b1;  wr_cycle[12980] = 1'b0;  addr_rom[12980]='h0000229c;  wr_data_rom[12980]='h00000000;
    rd_cycle[12981] = 1'b1;  wr_cycle[12981] = 1'b0;  addr_rom[12981]='h00002d08;  wr_data_rom[12981]='h00000000;
    rd_cycle[12982] = 1'b0;  wr_cycle[12982] = 1'b1;  addr_rom[12982]='h00003780;  wr_data_rom[12982]='h0000328a;
    rd_cycle[12983] = 1'b1;  wr_cycle[12983] = 1'b0;  addr_rom[12983]='h00003b68;  wr_data_rom[12983]='h00000000;
    rd_cycle[12984] = 1'b0;  wr_cycle[12984] = 1'b1;  addr_rom[12984]='h00001a08;  wr_data_rom[12984]='h00003d6b;
    rd_cycle[12985] = 1'b1;  wr_cycle[12985] = 1'b0;  addr_rom[12985]='h00000900;  wr_data_rom[12985]='h00000000;
    rd_cycle[12986] = 1'b1;  wr_cycle[12986] = 1'b0;  addr_rom[12986]='h00002c98;  wr_data_rom[12986]='h00000000;
    rd_cycle[12987] = 1'b0;  wr_cycle[12987] = 1'b1;  addr_rom[12987]='h0000068c;  wr_data_rom[12987]='h00002f28;
    rd_cycle[12988] = 1'b0;  wr_cycle[12988] = 1'b1;  addr_rom[12988]='h00002510;  wr_data_rom[12988]='h00000503;
    rd_cycle[12989] = 1'b1;  wr_cycle[12989] = 1'b0;  addr_rom[12989]='h00003cdc;  wr_data_rom[12989]='h00000000;
    rd_cycle[12990] = 1'b0;  wr_cycle[12990] = 1'b1;  addr_rom[12990]='h00001704;  wr_data_rom[12990]='h00000cb9;
    rd_cycle[12991] = 1'b0;  wr_cycle[12991] = 1'b1;  addr_rom[12991]='h00003d9c;  wr_data_rom[12991]='h0000388a;
    rd_cycle[12992] = 1'b1;  wr_cycle[12992] = 1'b0;  addr_rom[12992]='h00001d74;  wr_data_rom[12992]='h00000000;
    rd_cycle[12993] = 1'b0;  wr_cycle[12993] = 1'b1;  addr_rom[12993]='h000032dc;  wr_data_rom[12993]='h00003832;
    rd_cycle[12994] = 1'b1;  wr_cycle[12994] = 1'b0;  addr_rom[12994]='h00002424;  wr_data_rom[12994]='h00000000;
    rd_cycle[12995] = 1'b0;  wr_cycle[12995] = 1'b1;  addr_rom[12995]='h0000000c;  wr_data_rom[12995]='h000033d8;
    rd_cycle[12996] = 1'b1;  wr_cycle[12996] = 1'b0;  addr_rom[12996]='h00000794;  wr_data_rom[12996]='h00000000;
    rd_cycle[12997] = 1'b0;  wr_cycle[12997] = 1'b1;  addr_rom[12997]='h000033f4;  wr_data_rom[12997]='h0000373a;
    rd_cycle[12998] = 1'b1;  wr_cycle[12998] = 1'b0;  addr_rom[12998]='h000037f0;  wr_data_rom[12998]='h00000000;
    rd_cycle[12999] = 1'b1;  wr_cycle[12999] = 1'b0;  addr_rom[12999]='h00001d08;  wr_data_rom[12999]='h00000000;
    rd_cycle[13000] = 1'b0;  wr_cycle[13000] = 1'b1;  addr_rom[13000]='h00002a6c;  wr_data_rom[13000]='h00001673;
    rd_cycle[13001] = 1'b0;  wr_cycle[13001] = 1'b1;  addr_rom[13001]='h000020d8;  wr_data_rom[13001]='h000007bd;
    rd_cycle[13002] = 1'b0;  wr_cycle[13002] = 1'b1;  addr_rom[13002]='h000028ec;  wr_data_rom[13002]='h00003fa6;
    rd_cycle[13003] = 1'b1;  wr_cycle[13003] = 1'b0;  addr_rom[13003]='h00001658;  wr_data_rom[13003]='h00000000;
    rd_cycle[13004] = 1'b1;  wr_cycle[13004] = 1'b0;  addr_rom[13004]='h00003520;  wr_data_rom[13004]='h00000000;
    rd_cycle[13005] = 1'b0;  wr_cycle[13005] = 1'b1;  addr_rom[13005]='h000003d8;  wr_data_rom[13005]='h0000056a;
    rd_cycle[13006] = 1'b1;  wr_cycle[13006] = 1'b0;  addr_rom[13006]='h00000a34;  wr_data_rom[13006]='h00000000;
    rd_cycle[13007] = 1'b1;  wr_cycle[13007] = 1'b0;  addr_rom[13007]='h000011d8;  wr_data_rom[13007]='h00000000;
    rd_cycle[13008] = 1'b0;  wr_cycle[13008] = 1'b1;  addr_rom[13008]='h00000acc;  wr_data_rom[13008]='h0000189d;
    rd_cycle[13009] = 1'b1;  wr_cycle[13009] = 1'b0;  addr_rom[13009]='h00003700;  wr_data_rom[13009]='h00000000;
    rd_cycle[13010] = 1'b1;  wr_cycle[13010] = 1'b0;  addr_rom[13010]='h00001368;  wr_data_rom[13010]='h00000000;
    rd_cycle[13011] = 1'b1;  wr_cycle[13011] = 1'b0;  addr_rom[13011]='h000031f0;  wr_data_rom[13011]='h00000000;
    rd_cycle[13012] = 1'b1;  wr_cycle[13012] = 1'b0;  addr_rom[13012]='h00000c18;  wr_data_rom[13012]='h00000000;
    rd_cycle[13013] = 1'b0;  wr_cycle[13013] = 1'b1;  addr_rom[13013]='h000010ac;  wr_data_rom[13013]='h00003e20;
    rd_cycle[13014] = 1'b0;  wr_cycle[13014] = 1'b1;  addr_rom[13014]='h00003224;  wr_data_rom[13014]='h00000775;
    rd_cycle[13015] = 1'b0;  wr_cycle[13015] = 1'b1;  addr_rom[13015]='h00002734;  wr_data_rom[13015]='h00001f6b;
    rd_cycle[13016] = 1'b0;  wr_cycle[13016] = 1'b1;  addr_rom[13016]='h0000326c;  wr_data_rom[13016]='h00000e08;
    rd_cycle[13017] = 1'b1;  wr_cycle[13017] = 1'b0;  addr_rom[13017]='h00002474;  wr_data_rom[13017]='h00000000;
    rd_cycle[13018] = 1'b1;  wr_cycle[13018] = 1'b0;  addr_rom[13018]='h00001cbc;  wr_data_rom[13018]='h00000000;
    rd_cycle[13019] = 1'b0;  wr_cycle[13019] = 1'b1;  addr_rom[13019]='h00001220;  wr_data_rom[13019]='h00001255;
    rd_cycle[13020] = 1'b0;  wr_cycle[13020] = 1'b1;  addr_rom[13020]='h000034c0;  wr_data_rom[13020]='h00000bba;
    rd_cycle[13021] = 1'b1;  wr_cycle[13021] = 1'b0;  addr_rom[13021]='h00003538;  wr_data_rom[13021]='h00000000;
    rd_cycle[13022] = 1'b1;  wr_cycle[13022] = 1'b0;  addr_rom[13022]='h00000af0;  wr_data_rom[13022]='h00000000;
    rd_cycle[13023] = 1'b0;  wr_cycle[13023] = 1'b1;  addr_rom[13023]='h000021b0;  wr_data_rom[13023]='h00000f8b;
    rd_cycle[13024] = 1'b0;  wr_cycle[13024] = 1'b1;  addr_rom[13024]='h00003734;  wr_data_rom[13024]='h00000799;
    rd_cycle[13025] = 1'b1;  wr_cycle[13025] = 1'b0;  addr_rom[13025]='h00000610;  wr_data_rom[13025]='h00000000;
    rd_cycle[13026] = 1'b1;  wr_cycle[13026] = 1'b0;  addr_rom[13026]='h000026c4;  wr_data_rom[13026]='h00000000;
    rd_cycle[13027] = 1'b1;  wr_cycle[13027] = 1'b0;  addr_rom[13027]='h000018c0;  wr_data_rom[13027]='h00000000;
    rd_cycle[13028] = 1'b1;  wr_cycle[13028] = 1'b0;  addr_rom[13028]='h00002900;  wr_data_rom[13028]='h00000000;
    rd_cycle[13029] = 1'b1;  wr_cycle[13029] = 1'b0;  addr_rom[13029]='h0000322c;  wr_data_rom[13029]='h00000000;
    rd_cycle[13030] = 1'b1;  wr_cycle[13030] = 1'b0;  addr_rom[13030]='h00000414;  wr_data_rom[13030]='h00000000;
    rd_cycle[13031] = 1'b1;  wr_cycle[13031] = 1'b0;  addr_rom[13031]='h00003aec;  wr_data_rom[13031]='h00000000;
    rd_cycle[13032] = 1'b1;  wr_cycle[13032] = 1'b0;  addr_rom[13032]='h0000226c;  wr_data_rom[13032]='h00000000;
    rd_cycle[13033] = 1'b0;  wr_cycle[13033] = 1'b1;  addr_rom[13033]='h00003a58;  wr_data_rom[13033]='h0000311a;
    rd_cycle[13034] = 1'b0;  wr_cycle[13034] = 1'b1;  addr_rom[13034]='h00001870;  wr_data_rom[13034]='h000025a4;
    rd_cycle[13035] = 1'b0;  wr_cycle[13035] = 1'b1;  addr_rom[13035]='h000006e8;  wr_data_rom[13035]='h000030d7;
    rd_cycle[13036] = 1'b0;  wr_cycle[13036] = 1'b1;  addr_rom[13036]='h000035b8;  wr_data_rom[13036]='h00001147;
    rd_cycle[13037] = 1'b0;  wr_cycle[13037] = 1'b1;  addr_rom[13037]='h00002b1c;  wr_data_rom[13037]='h00001d92;
    rd_cycle[13038] = 1'b1;  wr_cycle[13038] = 1'b0;  addr_rom[13038]='h000015cc;  wr_data_rom[13038]='h00000000;
    rd_cycle[13039] = 1'b1;  wr_cycle[13039] = 1'b0;  addr_rom[13039]='h00002a80;  wr_data_rom[13039]='h00000000;
    rd_cycle[13040] = 1'b0;  wr_cycle[13040] = 1'b1;  addr_rom[13040]='h00002dbc;  wr_data_rom[13040]='h00002e40;
    rd_cycle[13041] = 1'b0;  wr_cycle[13041] = 1'b1;  addr_rom[13041]='h00003f90;  wr_data_rom[13041]='h00002e4d;
    rd_cycle[13042] = 1'b0;  wr_cycle[13042] = 1'b1;  addr_rom[13042]='h00002588;  wr_data_rom[13042]='h00000217;
    rd_cycle[13043] = 1'b1;  wr_cycle[13043] = 1'b0;  addr_rom[13043]='h0000328c;  wr_data_rom[13043]='h00000000;
    rd_cycle[13044] = 1'b1;  wr_cycle[13044] = 1'b0;  addr_rom[13044]='h00000c24;  wr_data_rom[13044]='h00000000;
    rd_cycle[13045] = 1'b0;  wr_cycle[13045] = 1'b1;  addr_rom[13045]='h00000a04;  wr_data_rom[13045]='h00001541;
    rd_cycle[13046] = 1'b0;  wr_cycle[13046] = 1'b1;  addr_rom[13046]='h00001ff8;  wr_data_rom[13046]='h00001981;
    rd_cycle[13047] = 1'b0;  wr_cycle[13047] = 1'b1;  addr_rom[13047]='h00001f28;  wr_data_rom[13047]='h0000232d;
    rd_cycle[13048] = 1'b1;  wr_cycle[13048] = 1'b0;  addr_rom[13048]='h00002968;  wr_data_rom[13048]='h00000000;
    rd_cycle[13049] = 1'b0;  wr_cycle[13049] = 1'b1;  addr_rom[13049]='h00000f18;  wr_data_rom[13049]='h000025c7;
    rd_cycle[13050] = 1'b0;  wr_cycle[13050] = 1'b1;  addr_rom[13050]='h00001a9c;  wr_data_rom[13050]='h00000129;
    rd_cycle[13051] = 1'b1;  wr_cycle[13051] = 1'b0;  addr_rom[13051]='h00003518;  wr_data_rom[13051]='h00000000;
    rd_cycle[13052] = 1'b1;  wr_cycle[13052] = 1'b0;  addr_rom[13052]='h0000148c;  wr_data_rom[13052]='h00000000;
    rd_cycle[13053] = 1'b0;  wr_cycle[13053] = 1'b1;  addr_rom[13053]='h00001b38;  wr_data_rom[13053]='h000029d5;
    rd_cycle[13054] = 1'b0;  wr_cycle[13054] = 1'b1;  addr_rom[13054]='h00000a64;  wr_data_rom[13054]='h0000122e;
    rd_cycle[13055] = 1'b1;  wr_cycle[13055] = 1'b0;  addr_rom[13055]='h000016e4;  wr_data_rom[13055]='h00000000;
    rd_cycle[13056] = 1'b1;  wr_cycle[13056] = 1'b0;  addr_rom[13056]='h00002aa0;  wr_data_rom[13056]='h00000000;
    rd_cycle[13057] = 1'b1;  wr_cycle[13057] = 1'b0;  addr_rom[13057]='h000018d4;  wr_data_rom[13057]='h00000000;
    rd_cycle[13058] = 1'b0;  wr_cycle[13058] = 1'b1;  addr_rom[13058]='h00001328;  wr_data_rom[13058]='h000014ea;
    rd_cycle[13059] = 1'b0;  wr_cycle[13059] = 1'b1;  addr_rom[13059]='h0000314c;  wr_data_rom[13059]='h000004e2;
    rd_cycle[13060] = 1'b0;  wr_cycle[13060] = 1'b1;  addr_rom[13060]='h00000264;  wr_data_rom[13060]='h0000308c;
    rd_cycle[13061] = 1'b1;  wr_cycle[13061] = 1'b0;  addr_rom[13061]='h00003410;  wr_data_rom[13061]='h00000000;
    rd_cycle[13062] = 1'b1;  wr_cycle[13062] = 1'b0;  addr_rom[13062]='h00001e20;  wr_data_rom[13062]='h00000000;
    rd_cycle[13063] = 1'b1;  wr_cycle[13063] = 1'b0;  addr_rom[13063]='h000015ec;  wr_data_rom[13063]='h00000000;
    rd_cycle[13064] = 1'b1;  wr_cycle[13064] = 1'b0;  addr_rom[13064]='h000025e0;  wr_data_rom[13064]='h00000000;
    rd_cycle[13065] = 1'b1;  wr_cycle[13065] = 1'b0;  addr_rom[13065]='h00003f30;  wr_data_rom[13065]='h00000000;
    rd_cycle[13066] = 1'b0;  wr_cycle[13066] = 1'b1;  addr_rom[13066]='h000003e8;  wr_data_rom[13066]='h0000083a;
    rd_cycle[13067] = 1'b1;  wr_cycle[13067] = 1'b0;  addr_rom[13067]='h00001464;  wr_data_rom[13067]='h00000000;
    rd_cycle[13068] = 1'b1;  wr_cycle[13068] = 1'b0;  addr_rom[13068]='h00003ad8;  wr_data_rom[13068]='h00000000;
    rd_cycle[13069] = 1'b0;  wr_cycle[13069] = 1'b1;  addr_rom[13069]='h00001408;  wr_data_rom[13069]='h00001d8a;
    rd_cycle[13070] = 1'b0;  wr_cycle[13070] = 1'b1;  addr_rom[13070]='h00001c7c;  wr_data_rom[13070]='h0000027f;
    rd_cycle[13071] = 1'b1;  wr_cycle[13071] = 1'b0;  addr_rom[13071]='h00002f48;  wr_data_rom[13071]='h00000000;
    rd_cycle[13072] = 1'b1;  wr_cycle[13072] = 1'b0;  addr_rom[13072]='h00002848;  wr_data_rom[13072]='h00000000;
    rd_cycle[13073] = 1'b0;  wr_cycle[13073] = 1'b1;  addr_rom[13073]='h000038c8;  wr_data_rom[13073]='h000024c2;
    rd_cycle[13074] = 1'b0;  wr_cycle[13074] = 1'b1;  addr_rom[13074]='h000020a8;  wr_data_rom[13074]='h00003831;
    rd_cycle[13075] = 1'b0;  wr_cycle[13075] = 1'b1;  addr_rom[13075]='h000037b8;  wr_data_rom[13075]='h00003baf;
    rd_cycle[13076] = 1'b1;  wr_cycle[13076] = 1'b0;  addr_rom[13076]='h000013b0;  wr_data_rom[13076]='h00000000;
    rd_cycle[13077] = 1'b0;  wr_cycle[13077] = 1'b1;  addr_rom[13077]='h00000460;  wr_data_rom[13077]='h000004d1;
    rd_cycle[13078] = 1'b1;  wr_cycle[13078] = 1'b0;  addr_rom[13078]='h00000f48;  wr_data_rom[13078]='h00000000;
    rd_cycle[13079] = 1'b1;  wr_cycle[13079] = 1'b0;  addr_rom[13079]='h000021b4;  wr_data_rom[13079]='h00000000;
    rd_cycle[13080] = 1'b0;  wr_cycle[13080] = 1'b1;  addr_rom[13080]='h000028b4;  wr_data_rom[13080]='h000006de;
    rd_cycle[13081] = 1'b0;  wr_cycle[13081] = 1'b1;  addr_rom[13081]='h00000738;  wr_data_rom[13081]='h00000cf5;
    rd_cycle[13082] = 1'b1;  wr_cycle[13082] = 1'b0;  addr_rom[13082]='h00001440;  wr_data_rom[13082]='h00000000;
    rd_cycle[13083] = 1'b0;  wr_cycle[13083] = 1'b1;  addr_rom[13083]='h00003654;  wr_data_rom[13083]='h00000fbd;
    rd_cycle[13084] = 1'b0;  wr_cycle[13084] = 1'b1;  addr_rom[13084]='h00002cdc;  wr_data_rom[13084]='h0000153e;
    rd_cycle[13085] = 1'b0;  wr_cycle[13085] = 1'b1;  addr_rom[13085]='h00001290;  wr_data_rom[13085]='h00001f3c;
    rd_cycle[13086] = 1'b1;  wr_cycle[13086] = 1'b0;  addr_rom[13086]='h00002008;  wr_data_rom[13086]='h00000000;
    rd_cycle[13087] = 1'b0;  wr_cycle[13087] = 1'b1;  addr_rom[13087]='h00001208;  wr_data_rom[13087]='h00002305;
    rd_cycle[13088] = 1'b0;  wr_cycle[13088] = 1'b1;  addr_rom[13088]='h00000090;  wr_data_rom[13088]='h00000864;
    rd_cycle[13089] = 1'b1;  wr_cycle[13089] = 1'b0;  addr_rom[13089]='h00003cfc;  wr_data_rom[13089]='h00000000;
    rd_cycle[13090] = 1'b1;  wr_cycle[13090] = 1'b0;  addr_rom[13090]='h000015cc;  wr_data_rom[13090]='h00000000;
    rd_cycle[13091] = 1'b0;  wr_cycle[13091] = 1'b1;  addr_rom[13091]='h00002218;  wr_data_rom[13091]='h000035e0;
    rd_cycle[13092] = 1'b1;  wr_cycle[13092] = 1'b0;  addr_rom[13092]='h00000224;  wr_data_rom[13092]='h00000000;
    rd_cycle[13093] = 1'b0;  wr_cycle[13093] = 1'b1;  addr_rom[13093]='h000015d4;  wr_data_rom[13093]='h000019c8;
    rd_cycle[13094] = 1'b1;  wr_cycle[13094] = 1'b0;  addr_rom[13094]='h000018f4;  wr_data_rom[13094]='h00000000;
    rd_cycle[13095] = 1'b0;  wr_cycle[13095] = 1'b1;  addr_rom[13095]='h00001c54;  wr_data_rom[13095]='h00001b0d;
    rd_cycle[13096] = 1'b1;  wr_cycle[13096] = 1'b0;  addr_rom[13096]='h00000ce0;  wr_data_rom[13096]='h00000000;
    rd_cycle[13097] = 1'b0;  wr_cycle[13097] = 1'b1;  addr_rom[13097]='h0000254c;  wr_data_rom[13097]='h00001bbc;
    rd_cycle[13098] = 1'b1;  wr_cycle[13098] = 1'b0;  addr_rom[13098]='h0000222c;  wr_data_rom[13098]='h00000000;
    rd_cycle[13099] = 1'b0;  wr_cycle[13099] = 1'b1;  addr_rom[13099]='h00001230;  wr_data_rom[13099]='h00002e73;
    rd_cycle[13100] = 1'b0;  wr_cycle[13100] = 1'b1;  addr_rom[13100]='h00003694;  wr_data_rom[13100]='h00002b51;
    rd_cycle[13101] = 1'b0;  wr_cycle[13101] = 1'b1;  addr_rom[13101]='h000031e4;  wr_data_rom[13101]='h00003a25;
    rd_cycle[13102] = 1'b0;  wr_cycle[13102] = 1'b1;  addr_rom[13102]='h00001868;  wr_data_rom[13102]='h00002a71;
    rd_cycle[13103] = 1'b1;  wr_cycle[13103] = 1'b0;  addr_rom[13103]='h00003878;  wr_data_rom[13103]='h00000000;
    rd_cycle[13104] = 1'b0;  wr_cycle[13104] = 1'b1;  addr_rom[13104]='h000023e4;  wr_data_rom[13104]='h00003bcb;
    rd_cycle[13105] = 1'b0;  wr_cycle[13105] = 1'b1;  addr_rom[13105]='h0000290c;  wr_data_rom[13105]='h00001da9;
    rd_cycle[13106] = 1'b1;  wr_cycle[13106] = 1'b0;  addr_rom[13106]='h00003388;  wr_data_rom[13106]='h00000000;
    rd_cycle[13107] = 1'b1;  wr_cycle[13107] = 1'b0;  addr_rom[13107]='h0000368c;  wr_data_rom[13107]='h00000000;
    rd_cycle[13108] = 1'b0;  wr_cycle[13108] = 1'b1;  addr_rom[13108]='h00001d9c;  wr_data_rom[13108]='h00003c9f;
    rd_cycle[13109] = 1'b1;  wr_cycle[13109] = 1'b0;  addr_rom[13109]='h00002c70;  wr_data_rom[13109]='h00000000;
    rd_cycle[13110] = 1'b0;  wr_cycle[13110] = 1'b1;  addr_rom[13110]='h00002094;  wr_data_rom[13110]='h00003b2c;
    rd_cycle[13111] = 1'b1;  wr_cycle[13111] = 1'b0;  addr_rom[13111]='h00001214;  wr_data_rom[13111]='h00000000;
    rd_cycle[13112] = 1'b1;  wr_cycle[13112] = 1'b0;  addr_rom[13112]='h000007f8;  wr_data_rom[13112]='h00000000;
    rd_cycle[13113] = 1'b0;  wr_cycle[13113] = 1'b1;  addr_rom[13113]='h00000d34;  wr_data_rom[13113]='h0000234a;
    rd_cycle[13114] = 1'b0;  wr_cycle[13114] = 1'b1;  addr_rom[13114]='h000022a8;  wr_data_rom[13114]='h000000b0;
    rd_cycle[13115] = 1'b1;  wr_cycle[13115] = 1'b0;  addr_rom[13115]='h000028f8;  wr_data_rom[13115]='h00000000;
    rd_cycle[13116] = 1'b1;  wr_cycle[13116] = 1'b0;  addr_rom[13116]='h00002cd8;  wr_data_rom[13116]='h00000000;
    rd_cycle[13117] = 1'b1;  wr_cycle[13117] = 1'b0;  addr_rom[13117]='h00002aec;  wr_data_rom[13117]='h00000000;
    rd_cycle[13118] = 1'b0;  wr_cycle[13118] = 1'b1;  addr_rom[13118]='h000035fc;  wr_data_rom[13118]='h00002a67;
    rd_cycle[13119] = 1'b0;  wr_cycle[13119] = 1'b1;  addr_rom[13119]='h000022dc;  wr_data_rom[13119]='h0000309d;
    rd_cycle[13120] = 1'b0;  wr_cycle[13120] = 1'b1;  addr_rom[13120]='h00002d30;  wr_data_rom[13120]='h000020ee;
    rd_cycle[13121] = 1'b0;  wr_cycle[13121] = 1'b1;  addr_rom[13121]='h00003e04;  wr_data_rom[13121]='h00000676;
    rd_cycle[13122] = 1'b1;  wr_cycle[13122] = 1'b0;  addr_rom[13122]='h00000448;  wr_data_rom[13122]='h00000000;
    rd_cycle[13123] = 1'b0;  wr_cycle[13123] = 1'b1;  addr_rom[13123]='h00001be4;  wr_data_rom[13123]='h0000121a;
    rd_cycle[13124] = 1'b1;  wr_cycle[13124] = 1'b0;  addr_rom[13124]='h000036ec;  wr_data_rom[13124]='h00000000;
    rd_cycle[13125] = 1'b0;  wr_cycle[13125] = 1'b1;  addr_rom[13125]='h0000317c;  wr_data_rom[13125]='h00002e9f;
    rd_cycle[13126] = 1'b1;  wr_cycle[13126] = 1'b0;  addr_rom[13126]='h00003354;  wr_data_rom[13126]='h00000000;
    rd_cycle[13127] = 1'b0;  wr_cycle[13127] = 1'b1;  addr_rom[13127]='h00000a50;  wr_data_rom[13127]='h000001ed;
    rd_cycle[13128] = 1'b1;  wr_cycle[13128] = 1'b0;  addr_rom[13128]='h00003124;  wr_data_rom[13128]='h00000000;
    rd_cycle[13129] = 1'b0;  wr_cycle[13129] = 1'b1;  addr_rom[13129]='h0000053c;  wr_data_rom[13129]='h00000a7c;
    rd_cycle[13130] = 1'b0;  wr_cycle[13130] = 1'b1;  addr_rom[13130]='h00000ba0;  wr_data_rom[13130]='h00003989;
    rd_cycle[13131] = 1'b1;  wr_cycle[13131] = 1'b0;  addr_rom[13131]='h000012ac;  wr_data_rom[13131]='h00000000;
    rd_cycle[13132] = 1'b0;  wr_cycle[13132] = 1'b1;  addr_rom[13132]='h00003b94;  wr_data_rom[13132]='h0000093b;
    rd_cycle[13133] = 1'b0;  wr_cycle[13133] = 1'b1;  addr_rom[13133]='h00003d4c;  wr_data_rom[13133]='h000006d4;
    rd_cycle[13134] = 1'b1;  wr_cycle[13134] = 1'b0;  addr_rom[13134]='h00000d74;  wr_data_rom[13134]='h00000000;
    rd_cycle[13135] = 1'b1;  wr_cycle[13135] = 1'b0;  addr_rom[13135]='h00002d20;  wr_data_rom[13135]='h00000000;
    rd_cycle[13136] = 1'b0;  wr_cycle[13136] = 1'b1;  addr_rom[13136]='h00000710;  wr_data_rom[13136]='h00000fa8;
    rd_cycle[13137] = 1'b0;  wr_cycle[13137] = 1'b1;  addr_rom[13137]='h000013a4;  wr_data_rom[13137]='h00001941;
    rd_cycle[13138] = 1'b0;  wr_cycle[13138] = 1'b1;  addr_rom[13138]='h000023f8;  wr_data_rom[13138]='h00001fd7;
    rd_cycle[13139] = 1'b1;  wr_cycle[13139] = 1'b0;  addr_rom[13139]='h00000864;  wr_data_rom[13139]='h00000000;
    rd_cycle[13140] = 1'b1;  wr_cycle[13140] = 1'b0;  addr_rom[13140]='h00000774;  wr_data_rom[13140]='h00000000;
    rd_cycle[13141] = 1'b1;  wr_cycle[13141] = 1'b0;  addr_rom[13141]='h000017a4;  wr_data_rom[13141]='h00000000;
    rd_cycle[13142] = 1'b0;  wr_cycle[13142] = 1'b1;  addr_rom[13142]='h00002758;  wr_data_rom[13142]='h00000188;
    rd_cycle[13143] = 1'b1;  wr_cycle[13143] = 1'b0;  addr_rom[13143]='h00002d08;  wr_data_rom[13143]='h00000000;
    rd_cycle[13144] = 1'b1;  wr_cycle[13144] = 1'b0;  addr_rom[13144]='h00003ba4;  wr_data_rom[13144]='h00000000;
    rd_cycle[13145] = 1'b1;  wr_cycle[13145] = 1'b0;  addr_rom[13145]='h0000377c;  wr_data_rom[13145]='h00000000;
    rd_cycle[13146] = 1'b1;  wr_cycle[13146] = 1'b0;  addr_rom[13146]='h00001224;  wr_data_rom[13146]='h00000000;
    rd_cycle[13147] = 1'b1;  wr_cycle[13147] = 1'b0;  addr_rom[13147]='h00001d3c;  wr_data_rom[13147]='h00000000;
    rd_cycle[13148] = 1'b0;  wr_cycle[13148] = 1'b1;  addr_rom[13148]='h00000b00;  wr_data_rom[13148]='h00001091;
    rd_cycle[13149] = 1'b0;  wr_cycle[13149] = 1'b1;  addr_rom[13149]='h00002860;  wr_data_rom[13149]='h00003797;
    rd_cycle[13150] = 1'b0;  wr_cycle[13150] = 1'b1;  addr_rom[13150]='h000005fc;  wr_data_rom[13150]='h00003750;
    rd_cycle[13151] = 1'b0;  wr_cycle[13151] = 1'b1;  addr_rom[13151]='h000029b0;  wr_data_rom[13151]='h00001ea6;
    rd_cycle[13152] = 1'b1;  wr_cycle[13152] = 1'b0;  addr_rom[13152]='h00000320;  wr_data_rom[13152]='h00000000;
    rd_cycle[13153] = 1'b1;  wr_cycle[13153] = 1'b0;  addr_rom[13153]='h00000f10;  wr_data_rom[13153]='h00000000;
    rd_cycle[13154] = 1'b0;  wr_cycle[13154] = 1'b1;  addr_rom[13154]='h0000318c;  wr_data_rom[13154]='h000017ef;
    rd_cycle[13155] = 1'b1;  wr_cycle[13155] = 1'b0;  addr_rom[13155]='h00003250;  wr_data_rom[13155]='h00000000;
    rd_cycle[13156] = 1'b0;  wr_cycle[13156] = 1'b1;  addr_rom[13156]='h00002a98;  wr_data_rom[13156]='h00003638;
    rd_cycle[13157] = 1'b1;  wr_cycle[13157] = 1'b0;  addr_rom[13157]='h00000e00;  wr_data_rom[13157]='h00000000;
    rd_cycle[13158] = 1'b0;  wr_cycle[13158] = 1'b1;  addr_rom[13158]='h0000205c;  wr_data_rom[13158]='h00000488;
    rd_cycle[13159] = 1'b0;  wr_cycle[13159] = 1'b1;  addr_rom[13159]='h00003df0;  wr_data_rom[13159]='h000017ed;
    rd_cycle[13160] = 1'b0;  wr_cycle[13160] = 1'b1;  addr_rom[13160]='h00001140;  wr_data_rom[13160]='h000014f6;
    rd_cycle[13161] = 1'b1;  wr_cycle[13161] = 1'b0;  addr_rom[13161]='h0000144c;  wr_data_rom[13161]='h00000000;
    rd_cycle[13162] = 1'b0;  wr_cycle[13162] = 1'b1;  addr_rom[13162]='h00003e68;  wr_data_rom[13162]='h000039f2;
    rd_cycle[13163] = 1'b1;  wr_cycle[13163] = 1'b0;  addr_rom[13163]='h000014b4;  wr_data_rom[13163]='h00000000;
    rd_cycle[13164] = 1'b0;  wr_cycle[13164] = 1'b1;  addr_rom[13164]='h00003d4c;  wr_data_rom[13164]='h000022c0;
    rd_cycle[13165] = 1'b1;  wr_cycle[13165] = 1'b0;  addr_rom[13165]='h00002380;  wr_data_rom[13165]='h00000000;
    rd_cycle[13166] = 1'b0;  wr_cycle[13166] = 1'b1;  addr_rom[13166]='h00001980;  wr_data_rom[13166]='h0000049e;
    rd_cycle[13167] = 1'b1;  wr_cycle[13167] = 1'b0;  addr_rom[13167]='h000037e4;  wr_data_rom[13167]='h00000000;
    rd_cycle[13168] = 1'b1;  wr_cycle[13168] = 1'b0;  addr_rom[13168]='h00000e1c;  wr_data_rom[13168]='h00000000;
    rd_cycle[13169] = 1'b1;  wr_cycle[13169] = 1'b0;  addr_rom[13169]='h00003534;  wr_data_rom[13169]='h00000000;
    rd_cycle[13170] = 1'b0;  wr_cycle[13170] = 1'b1;  addr_rom[13170]='h00001cc8;  wr_data_rom[13170]='h0000366b;
    rd_cycle[13171] = 1'b1;  wr_cycle[13171] = 1'b0;  addr_rom[13171]='h00000090;  wr_data_rom[13171]='h00000000;
    rd_cycle[13172] = 1'b1;  wr_cycle[13172] = 1'b0;  addr_rom[13172]='h000021fc;  wr_data_rom[13172]='h00000000;
    rd_cycle[13173] = 1'b0;  wr_cycle[13173] = 1'b1;  addr_rom[13173]='h00001758;  wr_data_rom[13173]='h00003a21;
    rd_cycle[13174] = 1'b0;  wr_cycle[13174] = 1'b1;  addr_rom[13174]='h0000192c;  wr_data_rom[13174]='h000031b3;
    rd_cycle[13175] = 1'b0;  wr_cycle[13175] = 1'b1;  addr_rom[13175]='h00000bd4;  wr_data_rom[13175]='h0000270d;
    rd_cycle[13176] = 1'b1;  wr_cycle[13176] = 1'b0;  addr_rom[13176]='h000020bc;  wr_data_rom[13176]='h00000000;
    rd_cycle[13177] = 1'b1;  wr_cycle[13177] = 1'b0;  addr_rom[13177]='h00003558;  wr_data_rom[13177]='h00000000;
    rd_cycle[13178] = 1'b0;  wr_cycle[13178] = 1'b1;  addr_rom[13178]='h0000336c;  wr_data_rom[13178]='h000030b2;
    rd_cycle[13179] = 1'b0;  wr_cycle[13179] = 1'b1;  addr_rom[13179]='h00002ac8;  wr_data_rom[13179]='h0000245f;
    rd_cycle[13180] = 1'b1;  wr_cycle[13180] = 1'b0;  addr_rom[13180]='h000028e8;  wr_data_rom[13180]='h00000000;
    rd_cycle[13181] = 1'b0;  wr_cycle[13181] = 1'b1;  addr_rom[13181]='h00003160;  wr_data_rom[13181]='h000029ca;
    rd_cycle[13182] = 1'b0;  wr_cycle[13182] = 1'b1;  addr_rom[13182]='h00000c74;  wr_data_rom[13182]='h00001a13;
    rd_cycle[13183] = 1'b1;  wr_cycle[13183] = 1'b0;  addr_rom[13183]='h00003ef4;  wr_data_rom[13183]='h00000000;
    rd_cycle[13184] = 1'b1;  wr_cycle[13184] = 1'b0;  addr_rom[13184]='h00002e80;  wr_data_rom[13184]='h00000000;
    rd_cycle[13185] = 1'b1;  wr_cycle[13185] = 1'b0;  addr_rom[13185]='h00000c24;  wr_data_rom[13185]='h00000000;
    rd_cycle[13186] = 1'b1;  wr_cycle[13186] = 1'b0;  addr_rom[13186]='h000009dc;  wr_data_rom[13186]='h00000000;
    rd_cycle[13187] = 1'b1;  wr_cycle[13187] = 1'b0;  addr_rom[13187]='h00002220;  wr_data_rom[13187]='h00000000;
    rd_cycle[13188] = 1'b1;  wr_cycle[13188] = 1'b0;  addr_rom[13188]='h00000060;  wr_data_rom[13188]='h00000000;
    rd_cycle[13189] = 1'b0;  wr_cycle[13189] = 1'b1;  addr_rom[13189]='h000037d8;  wr_data_rom[13189]='h0000252b;
    rd_cycle[13190] = 1'b1;  wr_cycle[13190] = 1'b0;  addr_rom[13190]='h000017ac;  wr_data_rom[13190]='h00000000;
    rd_cycle[13191] = 1'b0;  wr_cycle[13191] = 1'b1;  addr_rom[13191]='h00000258;  wr_data_rom[13191]='h00002f83;
    rd_cycle[13192] = 1'b0;  wr_cycle[13192] = 1'b1;  addr_rom[13192]='h00002174;  wr_data_rom[13192]='h000004a6;
    rd_cycle[13193] = 1'b1;  wr_cycle[13193] = 1'b0;  addr_rom[13193]='h000012e8;  wr_data_rom[13193]='h00000000;
    rd_cycle[13194] = 1'b1;  wr_cycle[13194] = 1'b0;  addr_rom[13194]='h000026c4;  wr_data_rom[13194]='h00000000;
    rd_cycle[13195] = 1'b1;  wr_cycle[13195] = 1'b0;  addr_rom[13195]='h000014b4;  wr_data_rom[13195]='h00000000;
    rd_cycle[13196] = 1'b1;  wr_cycle[13196] = 1'b0;  addr_rom[13196]='h000027b4;  wr_data_rom[13196]='h00000000;
    rd_cycle[13197] = 1'b0;  wr_cycle[13197] = 1'b1;  addr_rom[13197]='h00000e04;  wr_data_rom[13197]='h000012e4;
    rd_cycle[13198] = 1'b0;  wr_cycle[13198] = 1'b1;  addr_rom[13198]='h00001094;  wr_data_rom[13198]='h000012fa;
    rd_cycle[13199] = 1'b0;  wr_cycle[13199] = 1'b1;  addr_rom[13199]='h00001ac0;  wr_data_rom[13199]='h000034f3;
    rd_cycle[13200] = 1'b0;  wr_cycle[13200] = 1'b1;  addr_rom[13200]='h00001ce4;  wr_data_rom[13200]='h00000f24;
    rd_cycle[13201] = 1'b0;  wr_cycle[13201] = 1'b1;  addr_rom[13201]='h00001484;  wr_data_rom[13201]='h000023a5;
    rd_cycle[13202] = 1'b0;  wr_cycle[13202] = 1'b1;  addr_rom[13202]='h00000768;  wr_data_rom[13202]='h00001de4;
    rd_cycle[13203] = 1'b1;  wr_cycle[13203] = 1'b0;  addr_rom[13203]='h0000092c;  wr_data_rom[13203]='h00000000;
    rd_cycle[13204] = 1'b0;  wr_cycle[13204] = 1'b1;  addr_rom[13204]='h00001e1c;  wr_data_rom[13204]='h00001b27;
    rd_cycle[13205] = 1'b0;  wr_cycle[13205] = 1'b1;  addr_rom[13205]='h00000bb0;  wr_data_rom[13205]='h00002b21;
    rd_cycle[13206] = 1'b1;  wr_cycle[13206] = 1'b0;  addr_rom[13206]='h0000317c;  wr_data_rom[13206]='h00000000;
    rd_cycle[13207] = 1'b0;  wr_cycle[13207] = 1'b1;  addr_rom[13207]='h000015d8;  wr_data_rom[13207]='h0000157e;
    rd_cycle[13208] = 1'b0;  wr_cycle[13208] = 1'b1;  addr_rom[13208]='h00000570;  wr_data_rom[13208]='h0000366e;
    rd_cycle[13209] = 1'b1;  wr_cycle[13209] = 1'b0;  addr_rom[13209]='h00003540;  wr_data_rom[13209]='h00000000;
    rd_cycle[13210] = 1'b1;  wr_cycle[13210] = 1'b0;  addr_rom[13210]='h00000894;  wr_data_rom[13210]='h00000000;
    rd_cycle[13211] = 1'b0;  wr_cycle[13211] = 1'b1;  addr_rom[13211]='h000013a4;  wr_data_rom[13211]='h00002a61;
    rd_cycle[13212] = 1'b0;  wr_cycle[13212] = 1'b1;  addr_rom[13212]='h00001d28;  wr_data_rom[13212]='h00001b85;
    rd_cycle[13213] = 1'b0;  wr_cycle[13213] = 1'b1;  addr_rom[13213]='h00001264;  wr_data_rom[13213]='h00003ba1;
    rd_cycle[13214] = 1'b1;  wr_cycle[13214] = 1'b0;  addr_rom[13214]='h00001a2c;  wr_data_rom[13214]='h00000000;
    rd_cycle[13215] = 1'b1;  wr_cycle[13215] = 1'b0;  addr_rom[13215]='h00000780;  wr_data_rom[13215]='h00000000;
    rd_cycle[13216] = 1'b0;  wr_cycle[13216] = 1'b1;  addr_rom[13216]='h00002eac;  wr_data_rom[13216]='h0000178b;
    rd_cycle[13217] = 1'b0;  wr_cycle[13217] = 1'b1;  addr_rom[13217]='h0000364c;  wr_data_rom[13217]='h0000121e;
    rd_cycle[13218] = 1'b0;  wr_cycle[13218] = 1'b1;  addr_rom[13218]='h00000b14;  wr_data_rom[13218]='h0000364c;
    rd_cycle[13219] = 1'b0;  wr_cycle[13219] = 1'b1;  addr_rom[13219]='h00002fa4;  wr_data_rom[13219]='h000025c4;
    rd_cycle[13220] = 1'b0;  wr_cycle[13220] = 1'b1;  addr_rom[13220]='h00000ef0;  wr_data_rom[13220]='h00002357;
    rd_cycle[13221] = 1'b0;  wr_cycle[13221] = 1'b1;  addr_rom[13221]='h000005a8;  wr_data_rom[13221]='h000001ce;
    rd_cycle[13222] = 1'b1;  wr_cycle[13222] = 1'b0;  addr_rom[13222]='h000011e4;  wr_data_rom[13222]='h00000000;
    rd_cycle[13223] = 1'b0;  wr_cycle[13223] = 1'b1;  addr_rom[13223]='h0000281c;  wr_data_rom[13223]='h000015c6;
    rd_cycle[13224] = 1'b1;  wr_cycle[13224] = 1'b0;  addr_rom[13224]='h00000350;  wr_data_rom[13224]='h00000000;
    rd_cycle[13225] = 1'b0;  wr_cycle[13225] = 1'b1;  addr_rom[13225]='h00002e6c;  wr_data_rom[13225]='h000011b2;
    rd_cycle[13226] = 1'b1;  wr_cycle[13226] = 1'b0;  addr_rom[13226]='h00001a88;  wr_data_rom[13226]='h00000000;
    rd_cycle[13227] = 1'b0;  wr_cycle[13227] = 1'b1;  addr_rom[13227]='h000034e8;  wr_data_rom[13227]='h00001c56;
    rd_cycle[13228] = 1'b0;  wr_cycle[13228] = 1'b1;  addr_rom[13228]='h00001148;  wr_data_rom[13228]='h0000074d;
    rd_cycle[13229] = 1'b0;  wr_cycle[13229] = 1'b1;  addr_rom[13229]='h00002a74;  wr_data_rom[13229]='h00001aeb;
    rd_cycle[13230] = 1'b1;  wr_cycle[13230] = 1'b0;  addr_rom[13230]='h00002918;  wr_data_rom[13230]='h00000000;
    rd_cycle[13231] = 1'b1;  wr_cycle[13231] = 1'b0;  addr_rom[13231]='h0000357c;  wr_data_rom[13231]='h00000000;
    rd_cycle[13232] = 1'b1;  wr_cycle[13232] = 1'b0;  addr_rom[13232]='h00001630;  wr_data_rom[13232]='h00000000;
    rd_cycle[13233] = 1'b0;  wr_cycle[13233] = 1'b1;  addr_rom[13233]='h00000fe8;  wr_data_rom[13233]='h00002ce5;
    rd_cycle[13234] = 1'b1;  wr_cycle[13234] = 1'b0;  addr_rom[13234]='h000018ac;  wr_data_rom[13234]='h00000000;
    rd_cycle[13235] = 1'b0;  wr_cycle[13235] = 1'b1;  addr_rom[13235]='h00002910;  wr_data_rom[13235]='h000035a6;
    rd_cycle[13236] = 1'b0;  wr_cycle[13236] = 1'b1;  addr_rom[13236]='h00001a58;  wr_data_rom[13236]='h00002a29;
    rd_cycle[13237] = 1'b0;  wr_cycle[13237] = 1'b1;  addr_rom[13237]='h00001174;  wr_data_rom[13237]='h0000123c;
    rd_cycle[13238] = 1'b1;  wr_cycle[13238] = 1'b0;  addr_rom[13238]='h00002b60;  wr_data_rom[13238]='h00000000;
    rd_cycle[13239] = 1'b0;  wr_cycle[13239] = 1'b1;  addr_rom[13239]='h00000810;  wr_data_rom[13239]='h0000163b;
    rd_cycle[13240] = 1'b0;  wr_cycle[13240] = 1'b1;  addr_rom[13240]='h00003128;  wr_data_rom[13240]='h00001efe;
    rd_cycle[13241] = 1'b0;  wr_cycle[13241] = 1'b1;  addr_rom[13241]='h00000ce8;  wr_data_rom[13241]='h00001410;
    rd_cycle[13242] = 1'b1;  wr_cycle[13242] = 1'b0;  addr_rom[13242]='h00000990;  wr_data_rom[13242]='h00000000;
    rd_cycle[13243] = 1'b1;  wr_cycle[13243] = 1'b0;  addr_rom[13243]='h00003228;  wr_data_rom[13243]='h00000000;
    rd_cycle[13244] = 1'b1;  wr_cycle[13244] = 1'b0;  addr_rom[13244]='h00002b1c;  wr_data_rom[13244]='h00000000;
    rd_cycle[13245] = 1'b1;  wr_cycle[13245] = 1'b0;  addr_rom[13245]='h00002fe8;  wr_data_rom[13245]='h00000000;
    rd_cycle[13246] = 1'b1;  wr_cycle[13246] = 1'b0;  addr_rom[13246]='h000000ac;  wr_data_rom[13246]='h00000000;
    rd_cycle[13247] = 1'b0;  wr_cycle[13247] = 1'b1;  addr_rom[13247]='h000032b4;  wr_data_rom[13247]='h00000f2d;
    rd_cycle[13248] = 1'b1;  wr_cycle[13248] = 1'b0;  addr_rom[13248]='h00003c28;  wr_data_rom[13248]='h00000000;
    rd_cycle[13249] = 1'b0;  wr_cycle[13249] = 1'b1;  addr_rom[13249]='h000028ec;  wr_data_rom[13249]='h000019e4;
    rd_cycle[13250] = 1'b1;  wr_cycle[13250] = 1'b0;  addr_rom[13250]='h000023ec;  wr_data_rom[13250]='h00000000;
    rd_cycle[13251] = 1'b1;  wr_cycle[13251] = 1'b0;  addr_rom[13251]='h00000958;  wr_data_rom[13251]='h00000000;
    rd_cycle[13252] = 1'b1;  wr_cycle[13252] = 1'b0;  addr_rom[13252]='h00003594;  wr_data_rom[13252]='h00000000;
    rd_cycle[13253] = 1'b1;  wr_cycle[13253] = 1'b0;  addr_rom[13253]='h000009e0;  wr_data_rom[13253]='h00000000;
    rd_cycle[13254] = 1'b1;  wr_cycle[13254] = 1'b0;  addr_rom[13254]='h000039a8;  wr_data_rom[13254]='h00000000;
    rd_cycle[13255] = 1'b0;  wr_cycle[13255] = 1'b1;  addr_rom[13255]='h00003660;  wr_data_rom[13255]='h00000274;
    rd_cycle[13256] = 1'b1;  wr_cycle[13256] = 1'b0;  addr_rom[13256]='h00001474;  wr_data_rom[13256]='h00000000;
    rd_cycle[13257] = 1'b1;  wr_cycle[13257] = 1'b0;  addr_rom[13257]='h000039c4;  wr_data_rom[13257]='h00000000;
    rd_cycle[13258] = 1'b0;  wr_cycle[13258] = 1'b1;  addr_rom[13258]='h0000145c;  wr_data_rom[13258]='h000029c9;
    rd_cycle[13259] = 1'b0;  wr_cycle[13259] = 1'b1;  addr_rom[13259]='h00002708;  wr_data_rom[13259]='h00000b02;
    rd_cycle[13260] = 1'b0;  wr_cycle[13260] = 1'b1;  addr_rom[13260]='h00002034;  wr_data_rom[13260]='h00003a9a;
    rd_cycle[13261] = 1'b1;  wr_cycle[13261] = 1'b0;  addr_rom[13261]='h000004b4;  wr_data_rom[13261]='h00000000;
    rd_cycle[13262] = 1'b1;  wr_cycle[13262] = 1'b0;  addr_rom[13262]='h00000668;  wr_data_rom[13262]='h00000000;
    rd_cycle[13263] = 1'b1;  wr_cycle[13263] = 1'b0;  addr_rom[13263]='h00001008;  wr_data_rom[13263]='h00000000;
    rd_cycle[13264] = 1'b1;  wr_cycle[13264] = 1'b0;  addr_rom[13264]='h00003ef4;  wr_data_rom[13264]='h00000000;
    rd_cycle[13265] = 1'b1;  wr_cycle[13265] = 1'b0;  addr_rom[13265]='h000034cc;  wr_data_rom[13265]='h00000000;
    rd_cycle[13266] = 1'b0;  wr_cycle[13266] = 1'b1;  addr_rom[13266]='h0000284c;  wr_data_rom[13266]='h00001792;
    rd_cycle[13267] = 1'b1;  wr_cycle[13267] = 1'b0;  addr_rom[13267]='h000009c8;  wr_data_rom[13267]='h00000000;
    rd_cycle[13268] = 1'b0;  wr_cycle[13268] = 1'b1;  addr_rom[13268]='h00001eb0;  wr_data_rom[13268]='h00000b86;
    rd_cycle[13269] = 1'b1;  wr_cycle[13269] = 1'b0;  addr_rom[13269]='h00000870;  wr_data_rom[13269]='h00000000;
    rd_cycle[13270] = 1'b0;  wr_cycle[13270] = 1'b1;  addr_rom[13270]='h00000f34;  wr_data_rom[13270]='h00003f6e;
    rd_cycle[13271] = 1'b1;  wr_cycle[13271] = 1'b0;  addr_rom[13271]='h00002c80;  wr_data_rom[13271]='h00000000;
    rd_cycle[13272] = 1'b1;  wr_cycle[13272] = 1'b0;  addr_rom[13272]='h000020d8;  wr_data_rom[13272]='h00000000;
    rd_cycle[13273] = 1'b0;  wr_cycle[13273] = 1'b1;  addr_rom[13273]='h0000138c;  wr_data_rom[13273]='h00001b8f;
    rd_cycle[13274] = 1'b0;  wr_cycle[13274] = 1'b1;  addr_rom[13274]='h000026e0;  wr_data_rom[13274]='h00002d32;
    rd_cycle[13275] = 1'b0;  wr_cycle[13275] = 1'b1;  addr_rom[13275]='h00002520;  wr_data_rom[13275]='h00003b9e;
    rd_cycle[13276] = 1'b0;  wr_cycle[13276] = 1'b1;  addr_rom[13276]='h00001a70;  wr_data_rom[13276]='h0000089d;
    rd_cycle[13277] = 1'b1;  wr_cycle[13277] = 1'b0;  addr_rom[13277]='h000002d8;  wr_data_rom[13277]='h00000000;
    rd_cycle[13278] = 1'b0;  wr_cycle[13278] = 1'b1;  addr_rom[13278]='h00002234;  wr_data_rom[13278]='h00001f5e;
    rd_cycle[13279] = 1'b1;  wr_cycle[13279] = 1'b0;  addr_rom[13279]='h00003174;  wr_data_rom[13279]='h00000000;
    rd_cycle[13280] = 1'b0;  wr_cycle[13280] = 1'b1;  addr_rom[13280]='h00000880;  wr_data_rom[13280]='h000022fa;
    rd_cycle[13281] = 1'b0;  wr_cycle[13281] = 1'b1;  addr_rom[13281]='h00000498;  wr_data_rom[13281]='h00000cbe;
    rd_cycle[13282] = 1'b1;  wr_cycle[13282] = 1'b0;  addr_rom[13282]='h00003398;  wr_data_rom[13282]='h00000000;
    rd_cycle[13283] = 1'b0;  wr_cycle[13283] = 1'b1;  addr_rom[13283]='h00002ad4;  wr_data_rom[13283]='h000006b8;
    rd_cycle[13284] = 1'b0;  wr_cycle[13284] = 1'b1;  addr_rom[13284]='h00001d20;  wr_data_rom[13284]='h00001abd;
    rd_cycle[13285] = 1'b1;  wr_cycle[13285] = 1'b0;  addr_rom[13285]='h00003000;  wr_data_rom[13285]='h00000000;
    rd_cycle[13286] = 1'b1;  wr_cycle[13286] = 1'b0;  addr_rom[13286]='h00000e4c;  wr_data_rom[13286]='h00000000;
    rd_cycle[13287] = 1'b0;  wr_cycle[13287] = 1'b1;  addr_rom[13287]='h00001b2c;  wr_data_rom[13287]='h0000064e;
    rd_cycle[13288] = 1'b0;  wr_cycle[13288] = 1'b1;  addr_rom[13288]='h00000e18;  wr_data_rom[13288]='h00000af3;
    rd_cycle[13289] = 1'b0;  wr_cycle[13289] = 1'b1;  addr_rom[13289]='h00001974;  wr_data_rom[13289]='h00003186;
    rd_cycle[13290] = 1'b0;  wr_cycle[13290] = 1'b1;  addr_rom[13290]='h000027e4;  wr_data_rom[13290]='h00002d8f;
    rd_cycle[13291] = 1'b0;  wr_cycle[13291] = 1'b1;  addr_rom[13291]='h000037dc;  wr_data_rom[13291]='h00001762;
    rd_cycle[13292] = 1'b1;  wr_cycle[13292] = 1'b0;  addr_rom[13292]='h000017c0;  wr_data_rom[13292]='h00000000;
    rd_cycle[13293] = 1'b0;  wr_cycle[13293] = 1'b1;  addr_rom[13293]='h00002b48;  wr_data_rom[13293]='h000002c6;
    rd_cycle[13294] = 1'b1;  wr_cycle[13294] = 1'b0;  addr_rom[13294]='h0000395c;  wr_data_rom[13294]='h00000000;
    rd_cycle[13295] = 1'b0;  wr_cycle[13295] = 1'b1;  addr_rom[13295]='h000034a8;  wr_data_rom[13295]='h00001bab;
    rd_cycle[13296] = 1'b0;  wr_cycle[13296] = 1'b1;  addr_rom[13296]='h00003eec;  wr_data_rom[13296]='h000037e0;
    rd_cycle[13297] = 1'b1;  wr_cycle[13297] = 1'b0;  addr_rom[13297]='h000020bc;  wr_data_rom[13297]='h00000000;
    rd_cycle[13298] = 1'b1;  wr_cycle[13298] = 1'b0;  addr_rom[13298]='h000003dc;  wr_data_rom[13298]='h00000000;
    rd_cycle[13299] = 1'b0;  wr_cycle[13299] = 1'b1;  addr_rom[13299]='h000031b0;  wr_data_rom[13299]='h00002864;
    rd_cycle[13300] = 1'b1;  wr_cycle[13300] = 1'b0;  addr_rom[13300]='h000002f8;  wr_data_rom[13300]='h00000000;
    rd_cycle[13301] = 1'b1;  wr_cycle[13301] = 1'b0;  addr_rom[13301]='h000016b0;  wr_data_rom[13301]='h00000000;
    rd_cycle[13302] = 1'b0;  wr_cycle[13302] = 1'b1;  addr_rom[13302]='h00002b50;  wr_data_rom[13302]='h00001cf0;
    rd_cycle[13303] = 1'b0;  wr_cycle[13303] = 1'b1;  addr_rom[13303]='h000012c8;  wr_data_rom[13303]='h0000164a;
    rd_cycle[13304] = 1'b0;  wr_cycle[13304] = 1'b1;  addr_rom[13304]='h000008c8;  wr_data_rom[13304]='h00003333;
    rd_cycle[13305] = 1'b1;  wr_cycle[13305] = 1'b0;  addr_rom[13305]='h00000a5c;  wr_data_rom[13305]='h00000000;
    rd_cycle[13306] = 1'b1;  wr_cycle[13306] = 1'b0;  addr_rom[13306]='h00001780;  wr_data_rom[13306]='h00000000;
    rd_cycle[13307] = 1'b1;  wr_cycle[13307] = 1'b0;  addr_rom[13307]='h00003134;  wr_data_rom[13307]='h00000000;
    rd_cycle[13308] = 1'b0;  wr_cycle[13308] = 1'b1;  addr_rom[13308]='h00003914;  wr_data_rom[13308]='h00000434;
    rd_cycle[13309] = 1'b0;  wr_cycle[13309] = 1'b1;  addr_rom[13309]='h00003538;  wr_data_rom[13309]='h000028d2;
    rd_cycle[13310] = 1'b1;  wr_cycle[13310] = 1'b0;  addr_rom[13310]='h00001ba8;  wr_data_rom[13310]='h00000000;
    rd_cycle[13311] = 1'b1;  wr_cycle[13311] = 1'b0;  addr_rom[13311]='h0000009c;  wr_data_rom[13311]='h00000000;
    rd_cycle[13312] = 1'b1;  wr_cycle[13312] = 1'b0;  addr_rom[13312]='h00000dd8;  wr_data_rom[13312]='h00000000;
    rd_cycle[13313] = 1'b1;  wr_cycle[13313] = 1'b0;  addr_rom[13313]='h00002270;  wr_data_rom[13313]='h00000000;
    rd_cycle[13314] = 1'b1;  wr_cycle[13314] = 1'b0;  addr_rom[13314]='h000007a4;  wr_data_rom[13314]='h00000000;
    rd_cycle[13315] = 1'b0;  wr_cycle[13315] = 1'b1;  addr_rom[13315]='h00000ea4;  wr_data_rom[13315]='h00001783;
    rd_cycle[13316] = 1'b0;  wr_cycle[13316] = 1'b1;  addr_rom[13316]='h000005d4;  wr_data_rom[13316]='h00003acf;
    rd_cycle[13317] = 1'b1;  wr_cycle[13317] = 1'b0;  addr_rom[13317]='h0000382c;  wr_data_rom[13317]='h00000000;
    rd_cycle[13318] = 1'b0;  wr_cycle[13318] = 1'b1;  addr_rom[13318]='h00000024;  wr_data_rom[13318]='h000035da;
    rd_cycle[13319] = 1'b1;  wr_cycle[13319] = 1'b0;  addr_rom[13319]='h0000081c;  wr_data_rom[13319]='h00000000;
    rd_cycle[13320] = 1'b0;  wr_cycle[13320] = 1'b1;  addr_rom[13320]='h00002730;  wr_data_rom[13320]='h00003610;
    rd_cycle[13321] = 1'b0;  wr_cycle[13321] = 1'b1;  addr_rom[13321]='h00002930;  wr_data_rom[13321]='h00001a8a;
    rd_cycle[13322] = 1'b0;  wr_cycle[13322] = 1'b1;  addr_rom[13322]='h0000349c;  wr_data_rom[13322]='h00001c74;
    rd_cycle[13323] = 1'b0;  wr_cycle[13323] = 1'b1;  addr_rom[13323]='h00002948;  wr_data_rom[13323]='h00000d7c;
    rd_cycle[13324] = 1'b1;  wr_cycle[13324] = 1'b0;  addr_rom[13324]='h00000fc0;  wr_data_rom[13324]='h00000000;
    rd_cycle[13325] = 1'b1;  wr_cycle[13325] = 1'b0;  addr_rom[13325]='h00002f18;  wr_data_rom[13325]='h00000000;
    rd_cycle[13326] = 1'b0;  wr_cycle[13326] = 1'b1;  addr_rom[13326]='h00003e34;  wr_data_rom[13326]='h000003c5;
    rd_cycle[13327] = 1'b1;  wr_cycle[13327] = 1'b0;  addr_rom[13327]='h00001d28;  wr_data_rom[13327]='h00000000;
    rd_cycle[13328] = 1'b1;  wr_cycle[13328] = 1'b0;  addr_rom[13328]='h00001900;  wr_data_rom[13328]='h00000000;
    rd_cycle[13329] = 1'b1;  wr_cycle[13329] = 1'b0;  addr_rom[13329]='h00003274;  wr_data_rom[13329]='h00000000;
    rd_cycle[13330] = 1'b0;  wr_cycle[13330] = 1'b1;  addr_rom[13330]='h00002d9c;  wr_data_rom[13330]='h00001a74;
    rd_cycle[13331] = 1'b0;  wr_cycle[13331] = 1'b1;  addr_rom[13331]='h00001d90;  wr_data_rom[13331]='h000012b0;
    rd_cycle[13332] = 1'b1;  wr_cycle[13332] = 1'b0;  addr_rom[13332]='h000007b0;  wr_data_rom[13332]='h00000000;
    rd_cycle[13333] = 1'b0;  wr_cycle[13333] = 1'b1;  addr_rom[13333]='h00000fec;  wr_data_rom[13333]='h00003f78;
    rd_cycle[13334] = 1'b1;  wr_cycle[13334] = 1'b0;  addr_rom[13334]='h000004a8;  wr_data_rom[13334]='h00000000;
    rd_cycle[13335] = 1'b0;  wr_cycle[13335] = 1'b1;  addr_rom[13335]='h0000337c;  wr_data_rom[13335]='h000021d6;
    rd_cycle[13336] = 1'b0;  wr_cycle[13336] = 1'b1;  addr_rom[13336]='h00001abc;  wr_data_rom[13336]='h00002bd8;
    rd_cycle[13337] = 1'b1;  wr_cycle[13337] = 1'b0;  addr_rom[13337]='h00000928;  wr_data_rom[13337]='h00000000;
    rd_cycle[13338] = 1'b0;  wr_cycle[13338] = 1'b1;  addr_rom[13338]='h00000370;  wr_data_rom[13338]='h00000855;
    rd_cycle[13339] = 1'b1;  wr_cycle[13339] = 1'b0;  addr_rom[13339]='h00000df4;  wr_data_rom[13339]='h00000000;
    rd_cycle[13340] = 1'b1;  wr_cycle[13340] = 1'b0;  addr_rom[13340]='h000037cc;  wr_data_rom[13340]='h00000000;
    rd_cycle[13341] = 1'b1;  wr_cycle[13341] = 1'b0;  addr_rom[13341]='h00002210;  wr_data_rom[13341]='h00000000;
    rd_cycle[13342] = 1'b1;  wr_cycle[13342] = 1'b0;  addr_rom[13342]='h00003c5c;  wr_data_rom[13342]='h00000000;
    rd_cycle[13343] = 1'b1;  wr_cycle[13343] = 1'b0;  addr_rom[13343]='h00001a70;  wr_data_rom[13343]='h00000000;
    rd_cycle[13344] = 1'b0;  wr_cycle[13344] = 1'b1;  addr_rom[13344]='h00002b30;  wr_data_rom[13344]='h00001565;
    rd_cycle[13345] = 1'b0;  wr_cycle[13345] = 1'b1;  addr_rom[13345]='h00001e24;  wr_data_rom[13345]='h00003369;
    rd_cycle[13346] = 1'b1;  wr_cycle[13346] = 1'b0;  addr_rom[13346]='h0000048c;  wr_data_rom[13346]='h00000000;
    rd_cycle[13347] = 1'b1;  wr_cycle[13347] = 1'b0;  addr_rom[13347]='h000011b4;  wr_data_rom[13347]='h00000000;
    rd_cycle[13348] = 1'b1;  wr_cycle[13348] = 1'b0;  addr_rom[13348]='h000002e8;  wr_data_rom[13348]='h00000000;
    rd_cycle[13349] = 1'b0;  wr_cycle[13349] = 1'b1;  addr_rom[13349]='h000023a8;  wr_data_rom[13349]='h000015e9;
    rd_cycle[13350] = 1'b0;  wr_cycle[13350] = 1'b1;  addr_rom[13350]='h000010e0;  wr_data_rom[13350]='h0000100a;
    rd_cycle[13351] = 1'b0;  wr_cycle[13351] = 1'b1;  addr_rom[13351]='h000025f8;  wr_data_rom[13351]='h00002fed;
    rd_cycle[13352] = 1'b0;  wr_cycle[13352] = 1'b1;  addr_rom[13352]='h000028a8;  wr_data_rom[13352]='h000029bb;
    rd_cycle[13353] = 1'b1;  wr_cycle[13353] = 1'b0;  addr_rom[13353]='h00000544;  wr_data_rom[13353]='h00000000;
    rd_cycle[13354] = 1'b0;  wr_cycle[13354] = 1'b1;  addr_rom[13354]='h00001350;  wr_data_rom[13354]='h00000c90;
    rd_cycle[13355] = 1'b0;  wr_cycle[13355] = 1'b1;  addr_rom[13355]='h00003d10;  wr_data_rom[13355]='h00002805;
    rd_cycle[13356] = 1'b1;  wr_cycle[13356] = 1'b0;  addr_rom[13356]='h00001a88;  wr_data_rom[13356]='h00000000;
    rd_cycle[13357] = 1'b0;  wr_cycle[13357] = 1'b1;  addr_rom[13357]='h00000854;  wr_data_rom[13357]='h00001ee7;
    rd_cycle[13358] = 1'b1;  wr_cycle[13358] = 1'b0;  addr_rom[13358]='h000034dc;  wr_data_rom[13358]='h00000000;
    rd_cycle[13359] = 1'b0;  wr_cycle[13359] = 1'b1;  addr_rom[13359]='h00000c44;  wr_data_rom[13359]='h00001bd4;
    rd_cycle[13360] = 1'b1;  wr_cycle[13360] = 1'b0;  addr_rom[13360]='h00001548;  wr_data_rom[13360]='h00000000;
    rd_cycle[13361] = 1'b1;  wr_cycle[13361] = 1'b0;  addr_rom[13361]='h00000c7c;  wr_data_rom[13361]='h00000000;
    rd_cycle[13362] = 1'b1;  wr_cycle[13362] = 1'b0;  addr_rom[13362]='h00001a3c;  wr_data_rom[13362]='h00000000;
    rd_cycle[13363] = 1'b0;  wr_cycle[13363] = 1'b1;  addr_rom[13363]='h00002d50;  wr_data_rom[13363]='h00000894;
    rd_cycle[13364] = 1'b0;  wr_cycle[13364] = 1'b1;  addr_rom[13364]='h00003c64;  wr_data_rom[13364]='h00000ff4;
    rd_cycle[13365] = 1'b0;  wr_cycle[13365] = 1'b1;  addr_rom[13365]='h00000820;  wr_data_rom[13365]='h0000133e;
    rd_cycle[13366] = 1'b1;  wr_cycle[13366] = 1'b0;  addr_rom[13366]='h00000650;  wr_data_rom[13366]='h00000000;
    rd_cycle[13367] = 1'b1;  wr_cycle[13367] = 1'b0;  addr_rom[13367]='h0000374c;  wr_data_rom[13367]='h00000000;
    rd_cycle[13368] = 1'b0;  wr_cycle[13368] = 1'b1;  addr_rom[13368]='h00002b1c;  wr_data_rom[13368]='h00002b71;
    rd_cycle[13369] = 1'b0;  wr_cycle[13369] = 1'b1;  addr_rom[13369]='h00002b7c;  wr_data_rom[13369]='h00002401;
    rd_cycle[13370] = 1'b1;  wr_cycle[13370] = 1'b0;  addr_rom[13370]='h0000263c;  wr_data_rom[13370]='h00000000;
    rd_cycle[13371] = 1'b0;  wr_cycle[13371] = 1'b1;  addr_rom[13371]='h00000818;  wr_data_rom[13371]='h000033a2;
    rd_cycle[13372] = 1'b1;  wr_cycle[13372] = 1'b0;  addr_rom[13372]='h00001de8;  wr_data_rom[13372]='h00000000;
    rd_cycle[13373] = 1'b1;  wr_cycle[13373] = 1'b0;  addr_rom[13373]='h00003a6c;  wr_data_rom[13373]='h00000000;
    rd_cycle[13374] = 1'b0;  wr_cycle[13374] = 1'b1;  addr_rom[13374]='h00001124;  wr_data_rom[13374]='h00000cef;
    rd_cycle[13375] = 1'b1;  wr_cycle[13375] = 1'b0;  addr_rom[13375]='h00000f58;  wr_data_rom[13375]='h00000000;
    rd_cycle[13376] = 1'b1;  wr_cycle[13376] = 1'b0;  addr_rom[13376]='h000035e8;  wr_data_rom[13376]='h00000000;
    rd_cycle[13377] = 1'b0;  wr_cycle[13377] = 1'b1;  addr_rom[13377]='h00001788;  wr_data_rom[13377]='h000003d0;
    rd_cycle[13378] = 1'b0;  wr_cycle[13378] = 1'b1;  addr_rom[13378]='h00000ce0;  wr_data_rom[13378]='h000026c4;
    rd_cycle[13379] = 1'b0;  wr_cycle[13379] = 1'b1;  addr_rom[13379]='h00000954;  wr_data_rom[13379]='h000024b0;
    rd_cycle[13380] = 1'b0;  wr_cycle[13380] = 1'b1;  addr_rom[13380]='h000031e8;  wr_data_rom[13380]='h00002efe;
    rd_cycle[13381] = 1'b1;  wr_cycle[13381] = 1'b0;  addr_rom[13381]='h00002c78;  wr_data_rom[13381]='h00000000;
    rd_cycle[13382] = 1'b1;  wr_cycle[13382] = 1'b0;  addr_rom[13382]='h0000229c;  wr_data_rom[13382]='h00000000;
    rd_cycle[13383] = 1'b1;  wr_cycle[13383] = 1'b0;  addr_rom[13383]='h00003134;  wr_data_rom[13383]='h00000000;
    rd_cycle[13384] = 1'b0;  wr_cycle[13384] = 1'b1;  addr_rom[13384]='h00002008;  wr_data_rom[13384]='h00002d00;
    rd_cycle[13385] = 1'b0;  wr_cycle[13385] = 1'b1;  addr_rom[13385]='h00001ea8;  wr_data_rom[13385]='h000019ea;
    rd_cycle[13386] = 1'b0;  wr_cycle[13386] = 1'b1;  addr_rom[13386]='h0000305c;  wr_data_rom[13386]='h00002247;
    rd_cycle[13387] = 1'b0;  wr_cycle[13387] = 1'b1;  addr_rom[13387]='h00003d5c;  wr_data_rom[13387]='h000011b4;
    rd_cycle[13388] = 1'b0;  wr_cycle[13388] = 1'b1;  addr_rom[13388]='h00002c88;  wr_data_rom[13388]='h00003d56;
    rd_cycle[13389] = 1'b1;  wr_cycle[13389] = 1'b0;  addr_rom[13389]='h0000080c;  wr_data_rom[13389]='h00000000;
    rd_cycle[13390] = 1'b1;  wr_cycle[13390] = 1'b0;  addr_rom[13390]='h000011c8;  wr_data_rom[13390]='h00000000;
    rd_cycle[13391] = 1'b1;  wr_cycle[13391] = 1'b0;  addr_rom[13391]='h00001e48;  wr_data_rom[13391]='h00000000;
    rd_cycle[13392] = 1'b0;  wr_cycle[13392] = 1'b1;  addr_rom[13392]='h000029bc;  wr_data_rom[13392]='h000015e1;
    rd_cycle[13393] = 1'b0;  wr_cycle[13393] = 1'b1;  addr_rom[13393]='h00001b10;  wr_data_rom[13393]='h00000f17;
    rd_cycle[13394] = 1'b0;  wr_cycle[13394] = 1'b1;  addr_rom[13394]='h00001dfc;  wr_data_rom[13394]='h00001523;
    rd_cycle[13395] = 1'b0;  wr_cycle[13395] = 1'b1;  addr_rom[13395]='h00003ad4;  wr_data_rom[13395]='h00000963;
    rd_cycle[13396] = 1'b1;  wr_cycle[13396] = 1'b0;  addr_rom[13396]='h00001424;  wr_data_rom[13396]='h00000000;
    rd_cycle[13397] = 1'b1;  wr_cycle[13397] = 1'b0;  addr_rom[13397]='h0000289c;  wr_data_rom[13397]='h00000000;
    rd_cycle[13398] = 1'b1;  wr_cycle[13398] = 1'b0;  addr_rom[13398]='h00002f2c;  wr_data_rom[13398]='h00000000;
    rd_cycle[13399] = 1'b0;  wr_cycle[13399] = 1'b1;  addr_rom[13399]='h000018a8;  wr_data_rom[13399]='h00000632;
    rd_cycle[13400] = 1'b0;  wr_cycle[13400] = 1'b1;  addr_rom[13400]='h000032a4;  wr_data_rom[13400]='h000027a9;
    rd_cycle[13401] = 1'b0;  wr_cycle[13401] = 1'b1;  addr_rom[13401]='h00001534;  wr_data_rom[13401]='h00002c07;
    rd_cycle[13402] = 1'b1;  wr_cycle[13402] = 1'b0;  addr_rom[13402]='h00000da4;  wr_data_rom[13402]='h00000000;
    rd_cycle[13403] = 1'b0;  wr_cycle[13403] = 1'b1;  addr_rom[13403]='h00003dfc;  wr_data_rom[13403]='h00000a3e;
    rd_cycle[13404] = 1'b1;  wr_cycle[13404] = 1'b0;  addr_rom[13404]='h00002c48;  wr_data_rom[13404]='h00000000;
    rd_cycle[13405] = 1'b0;  wr_cycle[13405] = 1'b1;  addr_rom[13405]='h00001974;  wr_data_rom[13405]='h00001a2f;
    rd_cycle[13406] = 1'b0;  wr_cycle[13406] = 1'b1;  addr_rom[13406]='h00002748;  wr_data_rom[13406]='h000012ea;
    rd_cycle[13407] = 1'b0;  wr_cycle[13407] = 1'b1;  addr_rom[13407]='h0000068c;  wr_data_rom[13407]='h00001041;
    rd_cycle[13408] = 1'b0;  wr_cycle[13408] = 1'b1;  addr_rom[13408]='h00003fdc;  wr_data_rom[13408]='h00000ee7;
    rd_cycle[13409] = 1'b1;  wr_cycle[13409] = 1'b0;  addr_rom[13409]='h00003db4;  wr_data_rom[13409]='h00000000;
    rd_cycle[13410] = 1'b1;  wr_cycle[13410] = 1'b0;  addr_rom[13410]='h00003b98;  wr_data_rom[13410]='h00000000;
    rd_cycle[13411] = 1'b0;  wr_cycle[13411] = 1'b1;  addr_rom[13411]='h000034ec;  wr_data_rom[13411]='h000026c5;
    rd_cycle[13412] = 1'b1;  wr_cycle[13412] = 1'b0;  addr_rom[13412]='h00002e70;  wr_data_rom[13412]='h00000000;
    rd_cycle[13413] = 1'b1;  wr_cycle[13413] = 1'b0;  addr_rom[13413]='h000018f0;  wr_data_rom[13413]='h00000000;
    rd_cycle[13414] = 1'b0;  wr_cycle[13414] = 1'b1;  addr_rom[13414]='h000007cc;  wr_data_rom[13414]='h00002705;
    rd_cycle[13415] = 1'b1;  wr_cycle[13415] = 1'b0;  addr_rom[13415]='h000001f0;  wr_data_rom[13415]='h00000000;
    rd_cycle[13416] = 1'b0;  wr_cycle[13416] = 1'b1;  addr_rom[13416]='h00001584;  wr_data_rom[13416]='h00002240;
    rd_cycle[13417] = 1'b1;  wr_cycle[13417] = 1'b0;  addr_rom[13417]='h000038d8;  wr_data_rom[13417]='h00000000;
    rd_cycle[13418] = 1'b0;  wr_cycle[13418] = 1'b1;  addr_rom[13418]='h0000269c;  wr_data_rom[13418]='h00003a58;
    rd_cycle[13419] = 1'b0;  wr_cycle[13419] = 1'b1;  addr_rom[13419]='h00002a40;  wr_data_rom[13419]='h00000a75;
    rd_cycle[13420] = 1'b1;  wr_cycle[13420] = 1'b0;  addr_rom[13420]='h00001b00;  wr_data_rom[13420]='h00000000;
    rd_cycle[13421] = 1'b1;  wr_cycle[13421] = 1'b0;  addr_rom[13421]='h00002f28;  wr_data_rom[13421]='h00000000;
    rd_cycle[13422] = 1'b0;  wr_cycle[13422] = 1'b1;  addr_rom[13422]='h00003bcc;  wr_data_rom[13422]='h00003b5f;
    rd_cycle[13423] = 1'b0;  wr_cycle[13423] = 1'b1;  addr_rom[13423]='h000038c8;  wr_data_rom[13423]='h00000a41;
    rd_cycle[13424] = 1'b0;  wr_cycle[13424] = 1'b1;  addr_rom[13424]='h000003b0;  wr_data_rom[13424]='h00001689;
    rd_cycle[13425] = 1'b1;  wr_cycle[13425] = 1'b0;  addr_rom[13425]='h00003b30;  wr_data_rom[13425]='h00000000;
    rd_cycle[13426] = 1'b0;  wr_cycle[13426] = 1'b1;  addr_rom[13426]='h00002030;  wr_data_rom[13426]='h00001e2b;
    rd_cycle[13427] = 1'b0;  wr_cycle[13427] = 1'b1;  addr_rom[13427]='h00000108;  wr_data_rom[13427]='h00001680;
    rd_cycle[13428] = 1'b1;  wr_cycle[13428] = 1'b0;  addr_rom[13428]='h000028b4;  wr_data_rom[13428]='h00000000;
    rd_cycle[13429] = 1'b0;  wr_cycle[13429] = 1'b1;  addr_rom[13429]='h00003420;  wr_data_rom[13429]='h00000919;
    rd_cycle[13430] = 1'b0;  wr_cycle[13430] = 1'b1;  addr_rom[13430]='h00001b60;  wr_data_rom[13430]='h00002f99;
    rd_cycle[13431] = 1'b0;  wr_cycle[13431] = 1'b1;  addr_rom[13431]='h00002584;  wr_data_rom[13431]='h0000397a;
    rd_cycle[13432] = 1'b0;  wr_cycle[13432] = 1'b1;  addr_rom[13432]='h00003264;  wr_data_rom[13432]='h000025cd;
    rd_cycle[13433] = 1'b0;  wr_cycle[13433] = 1'b1;  addr_rom[13433]='h0000289c;  wr_data_rom[13433]='h0000356c;
    rd_cycle[13434] = 1'b1;  wr_cycle[13434] = 1'b0;  addr_rom[13434]='h00002d78;  wr_data_rom[13434]='h00000000;
    rd_cycle[13435] = 1'b1;  wr_cycle[13435] = 1'b0;  addr_rom[13435]='h00001360;  wr_data_rom[13435]='h00000000;
    rd_cycle[13436] = 1'b1;  wr_cycle[13436] = 1'b0;  addr_rom[13436]='h00003870;  wr_data_rom[13436]='h00000000;
    rd_cycle[13437] = 1'b1;  wr_cycle[13437] = 1'b0;  addr_rom[13437]='h00001790;  wr_data_rom[13437]='h00000000;
    rd_cycle[13438] = 1'b1;  wr_cycle[13438] = 1'b0;  addr_rom[13438]='h0000229c;  wr_data_rom[13438]='h00000000;
    rd_cycle[13439] = 1'b0;  wr_cycle[13439] = 1'b1;  addr_rom[13439]='h00003358;  wr_data_rom[13439]='h00002b04;
    rd_cycle[13440] = 1'b1;  wr_cycle[13440] = 1'b0;  addr_rom[13440]='h000009f0;  wr_data_rom[13440]='h00000000;
    rd_cycle[13441] = 1'b0;  wr_cycle[13441] = 1'b1;  addr_rom[13441]='h00001480;  wr_data_rom[13441]='h00001eeb;
    rd_cycle[13442] = 1'b0;  wr_cycle[13442] = 1'b1;  addr_rom[13442]='h00000d80;  wr_data_rom[13442]='h000000f1;
    rd_cycle[13443] = 1'b1;  wr_cycle[13443] = 1'b0;  addr_rom[13443]='h00001f60;  wr_data_rom[13443]='h00000000;
    rd_cycle[13444] = 1'b1;  wr_cycle[13444] = 1'b0;  addr_rom[13444]='h000024c8;  wr_data_rom[13444]='h00000000;
    rd_cycle[13445] = 1'b1;  wr_cycle[13445] = 1'b0;  addr_rom[13445]='h00000ff0;  wr_data_rom[13445]='h00000000;
    rd_cycle[13446] = 1'b0;  wr_cycle[13446] = 1'b1;  addr_rom[13446]='h00001464;  wr_data_rom[13446]='h0000368c;
    rd_cycle[13447] = 1'b1;  wr_cycle[13447] = 1'b0;  addr_rom[13447]='h0000360c;  wr_data_rom[13447]='h00000000;
    rd_cycle[13448] = 1'b1;  wr_cycle[13448] = 1'b0;  addr_rom[13448]='h00003a14;  wr_data_rom[13448]='h00000000;
    rd_cycle[13449] = 1'b0;  wr_cycle[13449] = 1'b1;  addr_rom[13449]='h00002818;  wr_data_rom[13449]='h000019a3;
    rd_cycle[13450] = 1'b1;  wr_cycle[13450] = 1'b0;  addr_rom[13450]='h00001e34;  wr_data_rom[13450]='h00000000;
    rd_cycle[13451] = 1'b1;  wr_cycle[13451] = 1'b0;  addr_rom[13451]='h00002d00;  wr_data_rom[13451]='h00000000;
    rd_cycle[13452] = 1'b1;  wr_cycle[13452] = 1'b0;  addr_rom[13452]='h00002b50;  wr_data_rom[13452]='h00000000;
    rd_cycle[13453] = 1'b0;  wr_cycle[13453] = 1'b1;  addr_rom[13453]='h000037ec;  wr_data_rom[13453]='h00002c45;
    rd_cycle[13454] = 1'b0;  wr_cycle[13454] = 1'b1;  addr_rom[13454]='h00001af8;  wr_data_rom[13454]='h00003b51;
    rd_cycle[13455] = 1'b0;  wr_cycle[13455] = 1'b1;  addr_rom[13455]='h000031f0;  wr_data_rom[13455]='h00000e0d;
    rd_cycle[13456] = 1'b0;  wr_cycle[13456] = 1'b1;  addr_rom[13456]='h00002950;  wr_data_rom[13456]='h00002ef6;
    rd_cycle[13457] = 1'b1;  wr_cycle[13457] = 1'b0;  addr_rom[13457]='h00001340;  wr_data_rom[13457]='h00000000;
    rd_cycle[13458] = 1'b0;  wr_cycle[13458] = 1'b1;  addr_rom[13458]='h00002e1c;  wr_data_rom[13458]='h0000222d;
    rd_cycle[13459] = 1'b1;  wr_cycle[13459] = 1'b0;  addr_rom[13459]='h000011ac;  wr_data_rom[13459]='h00000000;
    rd_cycle[13460] = 1'b1;  wr_cycle[13460] = 1'b0;  addr_rom[13460]='h00000eac;  wr_data_rom[13460]='h00000000;
    rd_cycle[13461] = 1'b0;  wr_cycle[13461] = 1'b1;  addr_rom[13461]='h0000302c;  wr_data_rom[13461]='h00003465;
    rd_cycle[13462] = 1'b0;  wr_cycle[13462] = 1'b1;  addr_rom[13462]='h000031a8;  wr_data_rom[13462]='h000033d9;
    rd_cycle[13463] = 1'b1;  wr_cycle[13463] = 1'b0;  addr_rom[13463]='h00003aa8;  wr_data_rom[13463]='h00000000;
    rd_cycle[13464] = 1'b0;  wr_cycle[13464] = 1'b1;  addr_rom[13464]='h000024ec;  wr_data_rom[13464]='h000027b0;
    rd_cycle[13465] = 1'b0;  wr_cycle[13465] = 1'b1;  addr_rom[13465]='h00002a30;  wr_data_rom[13465]='h000015d3;
    rd_cycle[13466] = 1'b1;  wr_cycle[13466] = 1'b0;  addr_rom[13466]='h00003090;  wr_data_rom[13466]='h00000000;
    rd_cycle[13467] = 1'b1;  wr_cycle[13467] = 1'b0;  addr_rom[13467]='h00002a70;  wr_data_rom[13467]='h00000000;
    rd_cycle[13468] = 1'b0;  wr_cycle[13468] = 1'b1;  addr_rom[13468]='h000000c8;  wr_data_rom[13468]='h000013f3;
    rd_cycle[13469] = 1'b1;  wr_cycle[13469] = 1'b0;  addr_rom[13469]='h0000373c;  wr_data_rom[13469]='h00000000;
    rd_cycle[13470] = 1'b1;  wr_cycle[13470] = 1'b0;  addr_rom[13470]='h00002ee0;  wr_data_rom[13470]='h00000000;
    rd_cycle[13471] = 1'b1;  wr_cycle[13471] = 1'b0;  addr_rom[13471]='h00003bac;  wr_data_rom[13471]='h00000000;
    rd_cycle[13472] = 1'b1;  wr_cycle[13472] = 1'b0;  addr_rom[13472]='h00002250;  wr_data_rom[13472]='h00000000;
    rd_cycle[13473] = 1'b0;  wr_cycle[13473] = 1'b1;  addr_rom[13473]='h000015bc;  wr_data_rom[13473]='h00003228;
    rd_cycle[13474] = 1'b0;  wr_cycle[13474] = 1'b1;  addr_rom[13474]='h00002b84;  wr_data_rom[13474]='h00002eab;
    rd_cycle[13475] = 1'b1;  wr_cycle[13475] = 1'b0;  addr_rom[13475]='h00003bc8;  wr_data_rom[13475]='h00000000;
    rd_cycle[13476] = 1'b1;  wr_cycle[13476] = 1'b0;  addr_rom[13476]='h00000508;  wr_data_rom[13476]='h00000000;
    rd_cycle[13477] = 1'b1;  wr_cycle[13477] = 1'b0;  addr_rom[13477]='h00001e10;  wr_data_rom[13477]='h00000000;
    rd_cycle[13478] = 1'b0;  wr_cycle[13478] = 1'b1;  addr_rom[13478]='h00001ab0;  wr_data_rom[13478]='h00002bb4;
    rd_cycle[13479] = 1'b0;  wr_cycle[13479] = 1'b1;  addr_rom[13479]='h00000abc;  wr_data_rom[13479]='h00003e4b;
    rd_cycle[13480] = 1'b1;  wr_cycle[13480] = 1'b0;  addr_rom[13480]='h00001050;  wr_data_rom[13480]='h00000000;
    rd_cycle[13481] = 1'b1;  wr_cycle[13481] = 1'b0;  addr_rom[13481]='h00003a14;  wr_data_rom[13481]='h00000000;
    rd_cycle[13482] = 1'b1;  wr_cycle[13482] = 1'b0;  addr_rom[13482]='h00002f74;  wr_data_rom[13482]='h00000000;
    rd_cycle[13483] = 1'b1;  wr_cycle[13483] = 1'b0;  addr_rom[13483]='h000022a8;  wr_data_rom[13483]='h00000000;
    rd_cycle[13484] = 1'b0;  wr_cycle[13484] = 1'b1;  addr_rom[13484]='h000002e0;  wr_data_rom[13484]='h00002a1f;
    rd_cycle[13485] = 1'b1;  wr_cycle[13485] = 1'b0;  addr_rom[13485]='h00001ec4;  wr_data_rom[13485]='h00000000;
    rd_cycle[13486] = 1'b1;  wr_cycle[13486] = 1'b0;  addr_rom[13486]='h00001c7c;  wr_data_rom[13486]='h00000000;
    rd_cycle[13487] = 1'b1;  wr_cycle[13487] = 1'b0;  addr_rom[13487]='h000031cc;  wr_data_rom[13487]='h00000000;
    rd_cycle[13488] = 1'b1;  wr_cycle[13488] = 1'b0;  addr_rom[13488]='h00003e34;  wr_data_rom[13488]='h00000000;
    rd_cycle[13489] = 1'b1;  wr_cycle[13489] = 1'b0;  addr_rom[13489]='h00003f88;  wr_data_rom[13489]='h00000000;
    rd_cycle[13490] = 1'b0;  wr_cycle[13490] = 1'b1;  addr_rom[13490]='h00001350;  wr_data_rom[13490]='h00000740;
    rd_cycle[13491] = 1'b1;  wr_cycle[13491] = 1'b0;  addr_rom[13491]='h00001e9c;  wr_data_rom[13491]='h00000000;
    rd_cycle[13492] = 1'b1;  wr_cycle[13492] = 1'b0;  addr_rom[13492]='h00001ec0;  wr_data_rom[13492]='h00000000;
    rd_cycle[13493] = 1'b1;  wr_cycle[13493] = 1'b0;  addr_rom[13493]='h00001630;  wr_data_rom[13493]='h00000000;
    rd_cycle[13494] = 1'b0;  wr_cycle[13494] = 1'b1;  addr_rom[13494]='h0000110c;  wr_data_rom[13494]='h00001e53;
    rd_cycle[13495] = 1'b1;  wr_cycle[13495] = 1'b0;  addr_rom[13495]='h000015ac;  wr_data_rom[13495]='h00000000;
    rd_cycle[13496] = 1'b0;  wr_cycle[13496] = 1'b1;  addr_rom[13496]='h00002b4c;  wr_data_rom[13496]='h00001d75;
    rd_cycle[13497] = 1'b0;  wr_cycle[13497] = 1'b1;  addr_rom[13497]='h00000b8c;  wr_data_rom[13497]='h00002213;
    rd_cycle[13498] = 1'b1;  wr_cycle[13498] = 1'b0;  addr_rom[13498]='h000038f0;  wr_data_rom[13498]='h00000000;
    rd_cycle[13499] = 1'b0;  wr_cycle[13499] = 1'b1;  addr_rom[13499]='h000022b8;  wr_data_rom[13499]='h00002943;
    rd_cycle[13500] = 1'b1;  wr_cycle[13500] = 1'b0;  addr_rom[13500]='h000014bc;  wr_data_rom[13500]='h00000000;
    rd_cycle[13501] = 1'b1;  wr_cycle[13501] = 1'b0;  addr_rom[13501]='h00003f50;  wr_data_rom[13501]='h00000000;
    rd_cycle[13502] = 1'b0;  wr_cycle[13502] = 1'b1;  addr_rom[13502]='h00003254;  wr_data_rom[13502]='h00001091;
    rd_cycle[13503] = 1'b0;  wr_cycle[13503] = 1'b1;  addr_rom[13503]='h00000e18;  wr_data_rom[13503]='h00001f2e;
    rd_cycle[13504] = 1'b1;  wr_cycle[13504] = 1'b0;  addr_rom[13504]='h00001840;  wr_data_rom[13504]='h00000000;
    rd_cycle[13505] = 1'b0;  wr_cycle[13505] = 1'b1;  addr_rom[13505]='h000039c4;  wr_data_rom[13505]='h00003a21;
    rd_cycle[13506] = 1'b0;  wr_cycle[13506] = 1'b1;  addr_rom[13506]='h000010f8;  wr_data_rom[13506]='h0000362c;
    rd_cycle[13507] = 1'b1;  wr_cycle[13507] = 1'b0;  addr_rom[13507]='h00003ef0;  wr_data_rom[13507]='h00000000;
    rd_cycle[13508] = 1'b0;  wr_cycle[13508] = 1'b1;  addr_rom[13508]='h00000844;  wr_data_rom[13508]='h00001202;
    rd_cycle[13509] = 1'b0;  wr_cycle[13509] = 1'b1;  addr_rom[13509]='h00001b24;  wr_data_rom[13509]='h000003ac;
    rd_cycle[13510] = 1'b1;  wr_cycle[13510] = 1'b0;  addr_rom[13510]='h00000564;  wr_data_rom[13510]='h00000000;
    rd_cycle[13511] = 1'b1;  wr_cycle[13511] = 1'b0;  addr_rom[13511]='h0000301c;  wr_data_rom[13511]='h00000000;
    rd_cycle[13512] = 1'b1;  wr_cycle[13512] = 1'b0;  addr_rom[13512]='h00001ad4;  wr_data_rom[13512]='h00000000;
    rd_cycle[13513] = 1'b0;  wr_cycle[13513] = 1'b1;  addr_rom[13513]='h00003a74;  wr_data_rom[13513]='h00000e28;
    rd_cycle[13514] = 1'b0;  wr_cycle[13514] = 1'b1;  addr_rom[13514]='h00001dd4;  wr_data_rom[13514]='h00003028;
    rd_cycle[13515] = 1'b1;  wr_cycle[13515] = 1'b0;  addr_rom[13515]='h000036b8;  wr_data_rom[13515]='h00000000;
    rd_cycle[13516] = 1'b0;  wr_cycle[13516] = 1'b1;  addr_rom[13516]='h00001a80;  wr_data_rom[13516]='h000033ef;
    rd_cycle[13517] = 1'b0;  wr_cycle[13517] = 1'b1;  addr_rom[13517]='h000007b0;  wr_data_rom[13517]='h000031b1;
    rd_cycle[13518] = 1'b1;  wr_cycle[13518] = 1'b0;  addr_rom[13518]='h00002540;  wr_data_rom[13518]='h00000000;
    rd_cycle[13519] = 1'b0;  wr_cycle[13519] = 1'b1;  addr_rom[13519]='h0000014c;  wr_data_rom[13519]='h00003e3f;
    rd_cycle[13520] = 1'b0;  wr_cycle[13520] = 1'b1;  addr_rom[13520]='h00001968;  wr_data_rom[13520]='h0000169c;
    rd_cycle[13521] = 1'b1;  wr_cycle[13521] = 1'b0;  addr_rom[13521]='h00003608;  wr_data_rom[13521]='h00000000;
    rd_cycle[13522] = 1'b1;  wr_cycle[13522] = 1'b0;  addr_rom[13522]='h0000095c;  wr_data_rom[13522]='h00000000;
    rd_cycle[13523] = 1'b1;  wr_cycle[13523] = 1'b0;  addr_rom[13523]='h0000179c;  wr_data_rom[13523]='h00000000;
    rd_cycle[13524] = 1'b1;  wr_cycle[13524] = 1'b0;  addr_rom[13524]='h000011f4;  wr_data_rom[13524]='h00000000;
    rd_cycle[13525] = 1'b1;  wr_cycle[13525] = 1'b0;  addr_rom[13525]='h00003230;  wr_data_rom[13525]='h00000000;
    rd_cycle[13526] = 1'b0;  wr_cycle[13526] = 1'b1;  addr_rom[13526]='h00001454;  wr_data_rom[13526]='h000007fa;
    rd_cycle[13527] = 1'b1;  wr_cycle[13527] = 1'b0;  addr_rom[13527]='h00001dc8;  wr_data_rom[13527]='h00000000;
    rd_cycle[13528] = 1'b1;  wr_cycle[13528] = 1'b0;  addr_rom[13528]='h00002954;  wr_data_rom[13528]='h00000000;
    rd_cycle[13529] = 1'b0;  wr_cycle[13529] = 1'b1;  addr_rom[13529]='h000006fc;  wr_data_rom[13529]='h00000487;
    rd_cycle[13530] = 1'b0;  wr_cycle[13530] = 1'b1;  addr_rom[13530]='h00003518;  wr_data_rom[13530]='h00000b6a;
    rd_cycle[13531] = 1'b1;  wr_cycle[13531] = 1'b0;  addr_rom[13531]='h000038b8;  wr_data_rom[13531]='h00000000;
    rd_cycle[13532] = 1'b0;  wr_cycle[13532] = 1'b1;  addr_rom[13532]='h00002d4c;  wr_data_rom[13532]='h00002b7d;
    rd_cycle[13533] = 1'b1;  wr_cycle[13533] = 1'b0;  addr_rom[13533]='h000032c8;  wr_data_rom[13533]='h00000000;
    rd_cycle[13534] = 1'b0;  wr_cycle[13534] = 1'b1;  addr_rom[13534]='h00002dac;  wr_data_rom[13534]='h000024c3;
    rd_cycle[13535] = 1'b1;  wr_cycle[13535] = 1'b0;  addr_rom[13535]='h000010d8;  wr_data_rom[13535]='h00000000;
    rd_cycle[13536] = 1'b1;  wr_cycle[13536] = 1'b0;  addr_rom[13536]='h00003c4c;  wr_data_rom[13536]='h00000000;
    rd_cycle[13537] = 1'b0;  wr_cycle[13537] = 1'b1;  addr_rom[13537]='h000010f4;  wr_data_rom[13537]='h000027b3;
    rd_cycle[13538] = 1'b0;  wr_cycle[13538] = 1'b1;  addr_rom[13538]='h00002ca0;  wr_data_rom[13538]='h00002ee1;
    rd_cycle[13539] = 1'b0;  wr_cycle[13539] = 1'b1;  addr_rom[13539]='h000024f0;  wr_data_rom[13539]='h0000110d;
    rd_cycle[13540] = 1'b0;  wr_cycle[13540] = 1'b1;  addr_rom[13540]='h00002c0c;  wr_data_rom[13540]='h00002040;
    rd_cycle[13541] = 1'b1;  wr_cycle[13541] = 1'b0;  addr_rom[13541]='h000018d8;  wr_data_rom[13541]='h00000000;
    rd_cycle[13542] = 1'b1;  wr_cycle[13542] = 1'b0;  addr_rom[13542]='h00001174;  wr_data_rom[13542]='h00000000;
    rd_cycle[13543] = 1'b1;  wr_cycle[13543] = 1'b0;  addr_rom[13543]='h000018dc;  wr_data_rom[13543]='h00000000;
    rd_cycle[13544] = 1'b0;  wr_cycle[13544] = 1'b1;  addr_rom[13544]='h000036e0;  wr_data_rom[13544]='h0000357a;
    rd_cycle[13545] = 1'b1;  wr_cycle[13545] = 1'b0;  addr_rom[13545]='h00003008;  wr_data_rom[13545]='h00000000;
    rd_cycle[13546] = 1'b0;  wr_cycle[13546] = 1'b1;  addr_rom[13546]='h0000174c;  wr_data_rom[13546]='h0000100a;
    rd_cycle[13547] = 1'b0;  wr_cycle[13547] = 1'b1;  addr_rom[13547]='h00000d1c;  wr_data_rom[13547]='h00002e6c;
    rd_cycle[13548] = 1'b1;  wr_cycle[13548] = 1'b0;  addr_rom[13548]='h00000c8c;  wr_data_rom[13548]='h00000000;
    rd_cycle[13549] = 1'b0;  wr_cycle[13549] = 1'b1;  addr_rom[13549]='h00002744;  wr_data_rom[13549]='h00002933;
    rd_cycle[13550] = 1'b0;  wr_cycle[13550] = 1'b1;  addr_rom[13550]='h000026c4;  wr_data_rom[13550]='h00001832;
    rd_cycle[13551] = 1'b1;  wr_cycle[13551] = 1'b0;  addr_rom[13551]='h00001280;  wr_data_rom[13551]='h00000000;
    rd_cycle[13552] = 1'b0;  wr_cycle[13552] = 1'b1;  addr_rom[13552]='h000016e8;  wr_data_rom[13552]='h00000aba;
    rd_cycle[13553] = 1'b0;  wr_cycle[13553] = 1'b1;  addr_rom[13553]='h00001b24;  wr_data_rom[13553]='h000032dd;
    rd_cycle[13554] = 1'b0;  wr_cycle[13554] = 1'b1;  addr_rom[13554]='h00001b04;  wr_data_rom[13554]='h00001a02;
    rd_cycle[13555] = 1'b0;  wr_cycle[13555] = 1'b1;  addr_rom[13555]='h000001d8;  wr_data_rom[13555]='h00003966;
    rd_cycle[13556] = 1'b1;  wr_cycle[13556] = 1'b0;  addr_rom[13556]='h000035ac;  wr_data_rom[13556]='h00000000;
    rd_cycle[13557] = 1'b0;  wr_cycle[13557] = 1'b1;  addr_rom[13557]='h00003e14;  wr_data_rom[13557]='h0000375e;
    rd_cycle[13558] = 1'b1;  wr_cycle[13558] = 1'b0;  addr_rom[13558]='h000027b4;  wr_data_rom[13558]='h00000000;
    rd_cycle[13559] = 1'b1;  wr_cycle[13559] = 1'b0;  addr_rom[13559]='h000023c8;  wr_data_rom[13559]='h00000000;
    rd_cycle[13560] = 1'b1;  wr_cycle[13560] = 1'b0;  addr_rom[13560]='h000036fc;  wr_data_rom[13560]='h00000000;
    rd_cycle[13561] = 1'b1;  wr_cycle[13561] = 1'b0;  addr_rom[13561]='h00002e90;  wr_data_rom[13561]='h00000000;
    rd_cycle[13562] = 1'b0;  wr_cycle[13562] = 1'b1;  addr_rom[13562]='h0000281c;  wr_data_rom[13562]='h000008b0;
    rd_cycle[13563] = 1'b0;  wr_cycle[13563] = 1'b1;  addr_rom[13563]='h00003d14;  wr_data_rom[13563]='h00002623;
    rd_cycle[13564] = 1'b0;  wr_cycle[13564] = 1'b1;  addr_rom[13564]='h000004f0;  wr_data_rom[13564]='h00001fc8;
    rd_cycle[13565] = 1'b0;  wr_cycle[13565] = 1'b1;  addr_rom[13565]='h000005a8;  wr_data_rom[13565]='h000024b7;
    rd_cycle[13566] = 1'b0;  wr_cycle[13566] = 1'b1;  addr_rom[13566]='h00002fe8;  wr_data_rom[13566]='h00000fa5;
    rd_cycle[13567] = 1'b1;  wr_cycle[13567] = 1'b0;  addr_rom[13567]='h00002074;  wr_data_rom[13567]='h00000000;
    rd_cycle[13568] = 1'b0;  wr_cycle[13568] = 1'b1;  addr_rom[13568]='h00000ed0;  wr_data_rom[13568]='h00001441;
    rd_cycle[13569] = 1'b0;  wr_cycle[13569] = 1'b1;  addr_rom[13569]='h00002724;  wr_data_rom[13569]='h00001a73;
    rd_cycle[13570] = 1'b1;  wr_cycle[13570] = 1'b0;  addr_rom[13570]='h00000594;  wr_data_rom[13570]='h00000000;
    rd_cycle[13571] = 1'b1;  wr_cycle[13571] = 1'b0;  addr_rom[13571]='h0000389c;  wr_data_rom[13571]='h00000000;
    rd_cycle[13572] = 1'b1;  wr_cycle[13572] = 1'b0;  addr_rom[13572]='h00003180;  wr_data_rom[13572]='h00000000;
    rd_cycle[13573] = 1'b0;  wr_cycle[13573] = 1'b1;  addr_rom[13573]='h000019c4;  wr_data_rom[13573]='h000010dd;
    rd_cycle[13574] = 1'b0;  wr_cycle[13574] = 1'b1;  addr_rom[13574]='h00000ae0;  wr_data_rom[13574]='h00001501;
    rd_cycle[13575] = 1'b1;  wr_cycle[13575] = 1'b0;  addr_rom[13575]='h00003738;  wr_data_rom[13575]='h00000000;
    rd_cycle[13576] = 1'b0;  wr_cycle[13576] = 1'b1;  addr_rom[13576]='h00002d44;  wr_data_rom[13576]='h00001f44;
    rd_cycle[13577] = 1'b1;  wr_cycle[13577] = 1'b0;  addr_rom[13577]='h00001354;  wr_data_rom[13577]='h00000000;
    rd_cycle[13578] = 1'b0;  wr_cycle[13578] = 1'b1;  addr_rom[13578]='h00002cbc;  wr_data_rom[13578]='h000010d3;
    rd_cycle[13579] = 1'b0;  wr_cycle[13579] = 1'b1;  addr_rom[13579]='h00001824;  wr_data_rom[13579]='h000027e2;
    rd_cycle[13580] = 1'b1;  wr_cycle[13580] = 1'b0;  addr_rom[13580]='h00003b94;  wr_data_rom[13580]='h00000000;
    rd_cycle[13581] = 1'b1;  wr_cycle[13581] = 1'b0;  addr_rom[13581]='h000023fc;  wr_data_rom[13581]='h00000000;
    rd_cycle[13582] = 1'b1;  wr_cycle[13582] = 1'b0;  addr_rom[13582]='h0000245c;  wr_data_rom[13582]='h00000000;
    rd_cycle[13583] = 1'b0;  wr_cycle[13583] = 1'b1;  addr_rom[13583]='h00001500;  wr_data_rom[13583]='h00002ba3;
    rd_cycle[13584] = 1'b1;  wr_cycle[13584] = 1'b0;  addr_rom[13584]='h00001098;  wr_data_rom[13584]='h00000000;
    rd_cycle[13585] = 1'b1;  wr_cycle[13585] = 1'b0;  addr_rom[13585]='h00002f44;  wr_data_rom[13585]='h00000000;
    rd_cycle[13586] = 1'b1;  wr_cycle[13586] = 1'b0;  addr_rom[13586]='h000012ec;  wr_data_rom[13586]='h00000000;
    rd_cycle[13587] = 1'b1;  wr_cycle[13587] = 1'b0;  addr_rom[13587]='h00001c14;  wr_data_rom[13587]='h00000000;
    rd_cycle[13588] = 1'b1;  wr_cycle[13588] = 1'b0;  addr_rom[13588]='h000002b0;  wr_data_rom[13588]='h00000000;
    rd_cycle[13589] = 1'b1;  wr_cycle[13589] = 1'b0;  addr_rom[13589]='h000013e4;  wr_data_rom[13589]='h00000000;
    rd_cycle[13590] = 1'b1;  wr_cycle[13590] = 1'b0;  addr_rom[13590]='h000013a0;  wr_data_rom[13590]='h00000000;
    rd_cycle[13591] = 1'b1;  wr_cycle[13591] = 1'b0;  addr_rom[13591]='h000029c8;  wr_data_rom[13591]='h00000000;
    rd_cycle[13592] = 1'b0;  wr_cycle[13592] = 1'b1;  addr_rom[13592]='h00001c7c;  wr_data_rom[13592]='h00000b78;
    rd_cycle[13593] = 1'b0;  wr_cycle[13593] = 1'b1;  addr_rom[13593]='h00002324;  wr_data_rom[13593]='h00003642;
    rd_cycle[13594] = 1'b1;  wr_cycle[13594] = 1'b0;  addr_rom[13594]='h0000287c;  wr_data_rom[13594]='h00000000;
    rd_cycle[13595] = 1'b1;  wr_cycle[13595] = 1'b0;  addr_rom[13595]='h000035c4;  wr_data_rom[13595]='h00000000;
    rd_cycle[13596] = 1'b1;  wr_cycle[13596] = 1'b0;  addr_rom[13596]='h000009f4;  wr_data_rom[13596]='h00000000;
    rd_cycle[13597] = 1'b1;  wr_cycle[13597] = 1'b0;  addr_rom[13597]='h0000325c;  wr_data_rom[13597]='h00000000;
    rd_cycle[13598] = 1'b1;  wr_cycle[13598] = 1'b0;  addr_rom[13598]='h00002bfc;  wr_data_rom[13598]='h00000000;
    rd_cycle[13599] = 1'b0;  wr_cycle[13599] = 1'b1;  addr_rom[13599]='h00001ad0;  wr_data_rom[13599]='h00003ec4;
    rd_cycle[13600] = 1'b1;  wr_cycle[13600] = 1'b0;  addr_rom[13600]='h00000a34;  wr_data_rom[13600]='h00000000;
    rd_cycle[13601] = 1'b1;  wr_cycle[13601] = 1'b0;  addr_rom[13601]='h000006e4;  wr_data_rom[13601]='h00000000;
    rd_cycle[13602] = 1'b1;  wr_cycle[13602] = 1'b0;  addr_rom[13602]='h0000065c;  wr_data_rom[13602]='h00000000;
    rd_cycle[13603] = 1'b0;  wr_cycle[13603] = 1'b1;  addr_rom[13603]='h00001d3c;  wr_data_rom[13603]='h0000282c;
    rd_cycle[13604] = 1'b1;  wr_cycle[13604] = 1'b0;  addr_rom[13604]='h00002ca8;  wr_data_rom[13604]='h00000000;
    rd_cycle[13605] = 1'b1;  wr_cycle[13605] = 1'b0;  addr_rom[13605]='h00003650;  wr_data_rom[13605]='h00000000;
    rd_cycle[13606] = 1'b1;  wr_cycle[13606] = 1'b0;  addr_rom[13606]='h00001420;  wr_data_rom[13606]='h00000000;
    rd_cycle[13607] = 1'b0;  wr_cycle[13607] = 1'b1;  addr_rom[13607]='h00000de8;  wr_data_rom[13607]='h00003f5e;
    rd_cycle[13608] = 1'b0;  wr_cycle[13608] = 1'b1;  addr_rom[13608]='h00000d10;  wr_data_rom[13608]='h00003fb3;
    rd_cycle[13609] = 1'b1;  wr_cycle[13609] = 1'b0;  addr_rom[13609]='h00002638;  wr_data_rom[13609]='h00000000;
    rd_cycle[13610] = 1'b1;  wr_cycle[13610] = 1'b0;  addr_rom[13610]='h00000014;  wr_data_rom[13610]='h00000000;
    rd_cycle[13611] = 1'b1;  wr_cycle[13611] = 1'b0;  addr_rom[13611]='h00002ee8;  wr_data_rom[13611]='h00000000;
    rd_cycle[13612] = 1'b1;  wr_cycle[13612] = 1'b0;  addr_rom[13612]='h00003348;  wr_data_rom[13612]='h00000000;
    rd_cycle[13613] = 1'b0;  wr_cycle[13613] = 1'b1;  addr_rom[13613]='h00000b1c;  wr_data_rom[13613]='h00001598;
    rd_cycle[13614] = 1'b1;  wr_cycle[13614] = 1'b0;  addr_rom[13614]='h00001618;  wr_data_rom[13614]='h00000000;
    rd_cycle[13615] = 1'b0;  wr_cycle[13615] = 1'b1;  addr_rom[13615]='h00000b4c;  wr_data_rom[13615]='h000039c6;
    rd_cycle[13616] = 1'b1;  wr_cycle[13616] = 1'b0;  addr_rom[13616]='h00002974;  wr_data_rom[13616]='h00000000;
    rd_cycle[13617] = 1'b0;  wr_cycle[13617] = 1'b1;  addr_rom[13617]='h000030cc;  wr_data_rom[13617]='h0000103d;
    rd_cycle[13618] = 1'b1;  wr_cycle[13618] = 1'b0;  addr_rom[13618]='h000008dc;  wr_data_rom[13618]='h00000000;
    rd_cycle[13619] = 1'b1;  wr_cycle[13619] = 1'b0;  addr_rom[13619]='h000000cc;  wr_data_rom[13619]='h00000000;
    rd_cycle[13620] = 1'b0;  wr_cycle[13620] = 1'b1;  addr_rom[13620]='h00000f28;  wr_data_rom[13620]='h00000be4;
    rd_cycle[13621] = 1'b1;  wr_cycle[13621] = 1'b0;  addr_rom[13621]='h000039a8;  wr_data_rom[13621]='h00000000;
    rd_cycle[13622] = 1'b1;  wr_cycle[13622] = 1'b0;  addr_rom[13622]='h00001fbc;  wr_data_rom[13622]='h00000000;
    rd_cycle[13623] = 1'b0;  wr_cycle[13623] = 1'b1;  addr_rom[13623]='h0000254c;  wr_data_rom[13623]='h00000478;
    rd_cycle[13624] = 1'b1;  wr_cycle[13624] = 1'b0;  addr_rom[13624]='h0000333c;  wr_data_rom[13624]='h00000000;
    rd_cycle[13625] = 1'b1;  wr_cycle[13625] = 1'b0;  addr_rom[13625]='h000031c4;  wr_data_rom[13625]='h00000000;
    rd_cycle[13626] = 1'b1;  wr_cycle[13626] = 1'b0;  addr_rom[13626]='h000006a4;  wr_data_rom[13626]='h00000000;
    rd_cycle[13627] = 1'b0;  wr_cycle[13627] = 1'b1;  addr_rom[13627]='h00003f18;  wr_data_rom[13627]='h0000070e;
    rd_cycle[13628] = 1'b1;  wr_cycle[13628] = 1'b0;  addr_rom[13628]='h0000037c;  wr_data_rom[13628]='h00000000;
    rd_cycle[13629] = 1'b1;  wr_cycle[13629] = 1'b0;  addr_rom[13629]='h00002ed8;  wr_data_rom[13629]='h00000000;
    rd_cycle[13630] = 1'b1;  wr_cycle[13630] = 1'b0;  addr_rom[13630]='h00000cd4;  wr_data_rom[13630]='h00000000;
    rd_cycle[13631] = 1'b0;  wr_cycle[13631] = 1'b1;  addr_rom[13631]='h000034c0;  wr_data_rom[13631]='h00001dab;
    rd_cycle[13632] = 1'b0;  wr_cycle[13632] = 1'b1;  addr_rom[13632]='h000003dc;  wr_data_rom[13632]='h00000b69;
    rd_cycle[13633] = 1'b0;  wr_cycle[13633] = 1'b1;  addr_rom[13633]='h00002b98;  wr_data_rom[13633]='h000001e0;
    rd_cycle[13634] = 1'b0;  wr_cycle[13634] = 1'b1;  addr_rom[13634]='h00002714;  wr_data_rom[13634]='h000019cb;
    rd_cycle[13635] = 1'b0;  wr_cycle[13635] = 1'b1;  addr_rom[13635]='h00001088;  wr_data_rom[13635]='h00003ec6;
    rd_cycle[13636] = 1'b0;  wr_cycle[13636] = 1'b1;  addr_rom[13636]='h000033cc;  wr_data_rom[13636]='h000024c5;
    rd_cycle[13637] = 1'b1;  wr_cycle[13637] = 1'b0;  addr_rom[13637]='h00000c24;  wr_data_rom[13637]='h00000000;
    rd_cycle[13638] = 1'b1;  wr_cycle[13638] = 1'b0;  addr_rom[13638]='h00003b6c;  wr_data_rom[13638]='h00000000;
    rd_cycle[13639] = 1'b1;  wr_cycle[13639] = 1'b0;  addr_rom[13639]='h00002c1c;  wr_data_rom[13639]='h00000000;
    rd_cycle[13640] = 1'b0;  wr_cycle[13640] = 1'b1;  addr_rom[13640]='h00003bd0;  wr_data_rom[13640]='h00002107;
    rd_cycle[13641] = 1'b1;  wr_cycle[13641] = 1'b0;  addr_rom[13641]='h00003f88;  wr_data_rom[13641]='h00000000;
    rd_cycle[13642] = 1'b0;  wr_cycle[13642] = 1'b1;  addr_rom[13642]='h000004e8;  wr_data_rom[13642]='h00003f74;
    rd_cycle[13643] = 1'b1;  wr_cycle[13643] = 1'b0;  addr_rom[13643]='h00000280;  wr_data_rom[13643]='h00000000;
    rd_cycle[13644] = 1'b0;  wr_cycle[13644] = 1'b1;  addr_rom[13644]='h00001054;  wr_data_rom[13644]='h00003af5;
    rd_cycle[13645] = 1'b1;  wr_cycle[13645] = 1'b0;  addr_rom[13645]='h00002fd4;  wr_data_rom[13645]='h00000000;
    rd_cycle[13646] = 1'b1;  wr_cycle[13646] = 1'b0;  addr_rom[13646]='h00001604;  wr_data_rom[13646]='h00000000;
    rd_cycle[13647] = 1'b0;  wr_cycle[13647] = 1'b1;  addr_rom[13647]='h0000216c;  wr_data_rom[13647]='h000017b9;
    rd_cycle[13648] = 1'b1;  wr_cycle[13648] = 1'b0;  addr_rom[13648]='h0000256c;  wr_data_rom[13648]='h00000000;
    rd_cycle[13649] = 1'b0;  wr_cycle[13649] = 1'b1;  addr_rom[13649]='h000018dc;  wr_data_rom[13649]='h00003cad;
    rd_cycle[13650] = 1'b0;  wr_cycle[13650] = 1'b1;  addr_rom[13650]='h000031d8;  wr_data_rom[13650]='h000027c7;
    rd_cycle[13651] = 1'b1;  wr_cycle[13651] = 1'b0;  addr_rom[13651]='h00000fc4;  wr_data_rom[13651]='h00000000;
    rd_cycle[13652] = 1'b1;  wr_cycle[13652] = 1'b0;  addr_rom[13652]='h00000688;  wr_data_rom[13652]='h00000000;
    rd_cycle[13653] = 1'b1;  wr_cycle[13653] = 1'b0;  addr_rom[13653]='h00003b24;  wr_data_rom[13653]='h00000000;
    rd_cycle[13654] = 1'b0;  wr_cycle[13654] = 1'b1;  addr_rom[13654]='h00002a58;  wr_data_rom[13654]='h0000013b;
    rd_cycle[13655] = 1'b0;  wr_cycle[13655] = 1'b1;  addr_rom[13655]='h00003990;  wr_data_rom[13655]='h00003528;
    rd_cycle[13656] = 1'b1;  wr_cycle[13656] = 1'b0;  addr_rom[13656]='h00002a54;  wr_data_rom[13656]='h00000000;
    rd_cycle[13657] = 1'b1;  wr_cycle[13657] = 1'b0;  addr_rom[13657]='h00003c70;  wr_data_rom[13657]='h00000000;
    rd_cycle[13658] = 1'b0;  wr_cycle[13658] = 1'b1;  addr_rom[13658]='h000024dc;  wr_data_rom[13658]='h000026a5;
    rd_cycle[13659] = 1'b1;  wr_cycle[13659] = 1'b0;  addr_rom[13659]='h000010b4;  wr_data_rom[13659]='h00000000;
    rd_cycle[13660] = 1'b0;  wr_cycle[13660] = 1'b1;  addr_rom[13660]='h000039cc;  wr_data_rom[13660]='h00000653;
    rd_cycle[13661] = 1'b1;  wr_cycle[13661] = 1'b0;  addr_rom[13661]='h000008cc;  wr_data_rom[13661]='h00000000;
    rd_cycle[13662] = 1'b0;  wr_cycle[13662] = 1'b1;  addr_rom[13662]='h000010b0;  wr_data_rom[13662]='h00000e69;
    rd_cycle[13663] = 1'b1;  wr_cycle[13663] = 1'b0;  addr_rom[13663]='h00000fd0;  wr_data_rom[13663]='h00000000;
    rd_cycle[13664] = 1'b0;  wr_cycle[13664] = 1'b1;  addr_rom[13664]='h000030ac;  wr_data_rom[13664]='h000017c7;
    rd_cycle[13665] = 1'b0;  wr_cycle[13665] = 1'b1;  addr_rom[13665]='h00000cb0;  wr_data_rom[13665]='h0000385f;
    rd_cycle[13666] = 1'b1;  wr_cycle[13666] = 1'b0;  addr_rom[13666]='h00001d94;  wr_data_rom[13666]='h00000000;
    rd_cycle[13667] = 1'b1;  wr_cycle[13667] = 1'b0;  addr_rom[13667]='h00003428;  wr_data_rom[13667]='h00000000;
    rd_cycle[13668] = 1'b1;  wr_cycle[13668] = 1'b0;  addr_rom[13668]='h00002350;  wr_data_rom[13668]='h00000000;
    rd_cycle[13669] = 1'b0;  wr_cycle[13669] = 1'b1;  addr_rom[13669]='h00000820;  wr_data_rom[13669]='h000021ae;
    rd_cycle[13670] = 1'b0;  wr_cycle[13670] = 1'b1;  addr_rom[13670]='h000005f4;  wr_data_rom[13670]='h00001985;
    rd_cycle[13671] = 1'b0;  wr_cycle[13671] = 1'b1;  addr_rom[13671]='h000005b0;  wr_data_rom[13671]='h00000c63;
    rd_cycle[13672] = 1'b1;  wr_cycle[13672] = 1'b0;  addr_rom[13672]='h0000312c;  wr_data_rom[13672]='h00000000;
    rd_cycle[13673] = 1'b0;  wr_cycle[13673] = 1'b1;  addr_rom[13673]='h0000321c;  wr_data_rom[13673]='h000005e9;
    rd_cycle[13674] = 1'b1;  wr_cycle[13674] = 1'b0;  addr_rom[13674]='h0000303c;  wr_data_rom[13674]='h00000000;
    rd_cycle[13675] = 1'b1;  wr_cycle[13675] = 1'b0;  addr_rom[13675]='h000018d0;  wr_data_rom[13675]='h00000000;
    rd_cycle[13676] = 1'b1;  wr_cycle[13676] = 1'b0;  addr_rom[13676]='h00002630;  wr_data_rom[13676]='h00000000;
    rd_cycle[13677] = 1'b0;  wr_cycle[13677] = 1'b1;  addr_rom[13677]='h000028d0;  wr_data_rom[13677]='h00002194;
    rd_cycle[13678] = 1'b1;  wr_cycle[13678] = 1'b0;  addr_rom[13678]='h0000293c;  wr_data_rom[13678]='h00000000;
    rd_cycle[13679] = 1'b1;  wr_cycle[13679] = 1'b0;  addr_rom[13679]='h00001fa8;  wr_data_rom[13679]='h00000000;
    rd_cycle[13680] = 1'b0;  wr_cycle[13680] = 1'b1;  addr_rom[13680]='h00002d38;  wr_data_rom[13680]='h00003790;
    rd_cycle[13681] = 1'b0;  wr_cycle[13681] = 1'b1;  addr_rom[13681]='h000030f0;  wr_data_rom[13681]='h000006cc;
    rd_cycle[13682] = 1'b1;  wr_cycle[13682] = 1'b0;  addr_rom[13682]='h00002224;  wr_data_rom[13682]='h00000000;
    rd_cycle[13683] = 1'b1;  wr_cycle[13683] = 1'b0;  addr_rom[13683]='h0000366c;  wr_data_rom[13683]='h00000000;
    rd_cycle[13684] = 1'b1;  wr_cycle[13684] = 1'b0;  addr_rom[13684]='h000026ec;  wr_data_rom[13684]='h00000000;
    rd_cycle[13685] = 1'b0;  wr_cycle[13685] = 1'b1;  addr_rom[13685]='h000017f4;  wr_data_rom[13685]='h0000227c;
    rd_cycle[13686] = 1'b1;  wr_cycle[13686] = 1'b0;  addr_rom[13686]='h000010d4;  wr_data_rom[13686]='h00000000;
    rd_cycle[13687] = 1'b0;  wr_cycle[13687] = 1'b1;  addr_rom[13687]='h00003138;  wr_data_rom[13687]='h000013d7;
    rd_cycle[13688] = 1'b0;  wr_cycle[13688] = 1'b1;  addr_rom[13688]='h00001cd4;  wr_data_rom[13688]='h00000a5a;
    rd_cycle[13689] = 1'b1;  wr_cycle[13689] = 1'b0;  addr_rom[13689]='h000017a4;  wr_data_rom[13689]='h00000000;
    rd_cycle[13690] = 1'b0;  wr_cycle[13690] = 1'b1;  addr_rom[13690]='h00001ee8;  wr_data_rom[13690]='h000002d5;
    rd_cycle[13691] = 1'b1;  wr_cycle[13691] = 1'b0;  addr_rom[13691]='h00000a78;  wr_data_rom[13691]='h00000000;
    rd_cycle[13692] = 1'b1;  wr_cycle[13692] = 1'b0;  addr_rom[13692]='h00000f44;  wr_data_rom[13692]='h00000000;
    rd_cycle[13693] = 1'b0;  wr_cycle[13693] = 1'b1;  addr_rom[13693]='h00003038;  wr_data_rom[13693]='h000010e8;
    rd_cycle[13694] = 1'b0;  wr_cycle[13694] = 1'b1;  addr_rom[13694]='h00001c7c;  wr_data_rom[13694]='h00000441;
    rd_cycle[13695] = 1'b1;  wr_cycle[13695] = 1'b0;  addr_rom[13695]='h000009e0;  wr_data_rom[13695]='h00000000;
    rd_cycle[13696] = 1'b1;  wr_cycle[13696] = 1'b0;  addr_rom[13696]='h00003d5c;  wr_data_rom[13696]='h00000000;
    rd_cycle[13697] = 1'b1;  wr_cycle[13697] = 1'b0;  addr_rom[13697]='h00001a00;  wr_data_rom[13697]='h00000000;
    rd_cycle[13698] = 1'b0;  wr_cycle[13698] = 1'b1;  addr_rom[13698]='h000017d0;  wr_data_rom[13698]='h00001fd4;
    rd_cycle[13699] = 1'b0;  wr_cycle[13699] = 1'b1;  addr_rom[13699]='h00002c6c;  wr_data_rom[13699]='h00003a6f;
    rd_cycle[13700] = 1'b1;  wr_cycle[13700] = 1'b0;  addr_rom[13700]='h00001e58;  wr_data_rom[13700]='h00000000;
    rd_cycle[13701] = 1'b1;  wr_cycle[13701] = 1'b0;  addr_rom[13701]='h00002c08;  wr_data_rom[13701]='h00000000;
    rd_cycle[13702] = 1'b1;  wr_cycle[13702] = 1'b0;  addr_rom[13702]='h00002b38;  wr_data_rom[13702]='h00000000;
    rd_cycle[13703] = 1'b1;  wr_cycle[13703] = 1'b0;  addr_rom[13703]='h00003ed0;  wr_data_rom[13703]='h00000000;
    rd_cycle[13704] = 1'b1;  wr_cycle[13704] = 1'b0;  addr_rom[13704]='h00003658;  wr_data_rom[13704]='h00000000;
    rd_cycle[13705] = 1'b1;  wr_cycle[13705] = 1'b0;  addr_rom[13705]='h00001da4;  wr_data_rom[13705]='h00000000;
    rd_cycle[13706] = 1'b1;  wr_cycle[13706] = 1'b0;  addr_rom[13706]='h00003714;  wr_data_rom[13706]='h00000000;
    rd_cycle[13707] = 1'b1;  wr_cycle[13707] = 1'b0;  addr_rom[13707]='h00001d4c;  wr_data_rom[13707]='h00000000;
    rd_cycle[13708] = 1'b1;  wr_cycle[13708] = 1'b0;  addr_rom[13708]='h00003ed8;  wr_data_rom[13708]='h00000000;
    rd_cycle[13709] = 1'b0;  wr_cycle[13709] = 1'b1;  addr_rom[13709]='h0000186c;  wr_data_rom[13709]='h00001a6a;
    rd_cycle[13710] = 1'b0;  wr_cycle[13710] = 1'b1;  addr_rom[13710]='h00001b28;  wr_data_rom[13710]='h00002110;
    rd_cycle[13711] = 1'b1;  wr_cycle[13711] = 1'b0;  addr_rom[13711]='h00001c1c;  wr_data_rom[13711]='h00000000;
    rd_cycle[13712] = 1'b1;  wr_cycle[13712] = 1'b0;  addr_rom[13712]='h00002aac;  wr_data_rom[13712]='h00000000;
    rd_cycle[13713] = 1'b1;  wr_cycle[13713] = 1'b0;  addr_rom[13713]='h00002b10;  wr_data_rom[13713]='h00000000;
    rd_cycle[13714] = 1'b0;  wr_cycle[13714] = 1'b1;  addr_rom[13714]='h00000b88;  wr_data_rom[13714]='h00002a5e;
    rd_cycle[13715] = 1'b0;  wr_cycle[13715] = 1'b1;  addr_rom[13715]='h00000b5c;  wr_data_rom[13715]='h000003dc;
    rd_cycle[13716] = 1'b1;  wr_cycle[13716] = 1'b0;  addr_rom[13716]='h000033d4;  wr_data_rom[13716]='h00000000;
    rd_cycle[13717] = 1'b1;  wr_cycle[13717] = 1'b0;  addr_rom[13717]='h0000207c;  wr_data_rom[13717]='h00000000;
    rd_cycle[13718] = 1'b0;  wr_cycle[13718] = 1'b1;  addr_rom[13718]='h00001c60;  wr_data_rom[13718]='h00003ca1;
    rd_cycle[13719] = 1'b0;  wr_cycle[13719] = 1'b1;  addr_rom[13719]='h000002f0;  wr_data_rom[13719]='h00000102;
    rd_cycle[13720] = 1'b1;  wr_cycle[13720] = 1'b0;  addr_rom[13720]='h000020d4;  wr_data_rom[13720]='h00000000;
    rd_cycle[13721] = 1'b0;  wr_cycle[13721] = 1'b1;  addr_rom[13721]='h00003684;  wr_data_rom[13721]='h00002b54;
    rd_cycle[13722] = 1'b1;  wr_cycle[13722] = 1'b0;  addr_rom[13722]='h00000368;  wr_data_rom[13722]='h00000000;
    rd_cycle[13723] = 1'b0;  wr_cycle[13723] = 1'b1;  addr_rom[13723]='h0000082c;  wr_data_rom[13723]='h00001992;
    rd_cycle[13724] = 1'b0;  wr_cycle[13724] = 1'b1;  addr_rom[13724]='h0000369c;  wr_data_rom[13724]='h00001200;
    rd_cycle[13725] = 1'b0;  wr_cycle[13725] = 1'b1;  addr_rom[13725]='h000026ac;  wr_data_rom[13725]='h00002ddc;
    rd_cycle[13726] = 1'b1;  wr_cycle[13726] = 1'b0;  addr_rom[13726]='h00000e0c;  wr_data_rom[13726]='h00000000;
    rd_cycle[13727] = 1'b0;  wr_cycle[13727] = 1'b1;  addr_rom[13727]='h000018dc;  wr_data_rom[13727]='h00000195;
    rd_cycle[13728] = 1'b1;  wr_cycle[13728] = 1'b0;  addr_rom[13728]='h00001c18;  wr_data_rom[13728]='h00000000;
    rd_cycle[13729] = 1'b0;  wr_cycle[13729] = 1'b1;  addr_rom[13729]='h000005bc;  wr_data_rom[13729]='h0000082a;
    rd_cycle[13730] = 1'b1;  wr_cycle[13730] = 1'b0;  addr_rom[13730]='h0000072c;  wr_data_rom[13730]='h00000000;
    rd_cycle[13731] = 1'b0;  wr_cycle[13731] = 1'b1;  addr_rom[13731]='h000009ec;  wr_data_rom[13731]='h000002d9;
    rd_cycle[13732] = 1'b1;  wr_cycle[13732] = 1'b0;  addr_rom[13732]='h00000570;  wr_data_rom[13732]='h00000000;
    rd_cycle[13733] = 1'b0;  wr_cycle[13733] = 1'b1;  addr_rom[13733]='h00001b24;  wr_data_rom[13733]='h0000192f;
    rd_cycle[13734] = 1'b1;  wr_cycle[13734] = 1'b0;  addr_rom[13734]='h00002128;  wr_data_rom[13734]='h00000000;
    rd_cycle[13735] = 1'b1;  wr_cycle[13735] = 1'b0;  addr_rom[13735]='h000012cc;  wr_data_rom[13735]='h00000000;
    rd_cycle[13736] = 1'b0;  wr_cycle[13736] = 1'b1;  addr_rom[13736]='h00001b1c;  wr_data_rom[13736]='h00000a5e;
    rd_cycle[13737] = 1'b0;  wr_cycle[13737] = 1'b1;  addr_rom[13737]='h00000e10;  wr_data_rom[13737]='h00000659;
    rd_cycle[13738] = 1'b1;  wr_cycle[13738] = 1'b0;  addr_rom[13738]='h00002bbc;  wr_data_rom[13738]='h00000000;
    rd_cycle[13739] = 1'b0;  wr_cycle[13739] = 1'b1;  addr_rom[13739]='h00002cac;  wr_data_rom[13739]='h00002db7;
    rd_cycle[13740] = 1'b1;  wr_cycle[13740] = 1'b0;  addr_rom[13740]='h00003eec;  wr_data_rom[13740]='h00000000;
    rd_cycle[13741] = 1'b1;  wr_cycle[13741] = 1'b0;  addr_rom[13741]='h00000f14;  wr_data_rom[13741]='h00000000;
    rd_cycle[13742] = 1'b0;  wr_cycle[13742] = 1'b1;  addr_rom[13742]='h00002d28;  wr_data_rom[13742]='h000033cc;
    rd_cycle[13743] = 1'b1;  wr_cycle[13743] = 1'b0;  addr_rom[13743]='h00000074;  wr_data_rom[13743]='h00000000;
    rd_cycle[13744] = 1'b1;  wr_cycle[13744] = 1'b0;  addr_rom[13744]='h00003f4c;  wr_data_rom[13744]='h00000000;
    rd_cycle[13745] = 1'b0;  wr_cycle[13745] = 1'b1;  addr_rom[13745]='h00002680;  wr_data_rom[13745]='h00001ebd;
    rd_cycle[13746] = 1'b0;  wr_cycle[13746] = 1'b1;  addr_rom[13746]='h00001b98;  wr_data_rom[13746]='h0000211f;
    rd_cycle[13747] = 1'b1;  wr_cycle[13747] = 1'b0;  addr_rom[13747]='h00000710;  wr_data_rom[13747]='h00000000;
    rd_cycle[13748] = 1'b1;  wr_cycle[13748] = 1'b0;  addr_rom[13748]='h00003c10;  wr_data_rom[13748]='h00000000;
    rd_cycle[13749] = 1'b0;  wr_cycle[13749] = 1'b1;  addr_rom[13749]='h00001cec;  wr_data_rom[13749]='h00001c4c;
    rd_cycle[13750] = 1'b0;  wr_cycle[13750] = 1'b1;  addr_rom[13750]='h000010a0;  wr_data_rom[13750]='h00002096;
    rd_cycle[13751] = 1'b1;  wr_cycle[13751] = 1'b0;  addr_rom[13751]='h000024d4;  wr_data_rom[13751]='h00000000;
    rd_cycle[13752] = 1'b1;  wr_cycle[13752] = 1'b0;  addr_rom[13752]='h000033d4;  wr_data_rom[13752]='h00000000;
    rd_cycle[13753] = 1'b0;  wr_cycle[13753] = 1'b1;  addr_rom[13753]='h000009fc;  wr_data_rom[13753]='h000001fe;
    rd_cycle[13754] = 1'b1;  wr_cycle[13754] = 1'b0;  addr_rom[13754]='h00003e5c;  wr_data_rom[13754]='h00000000;
    rd_cycle[13755] = 1'b0;  wr_cycle[13755] = 1'b1;  addr_rom[13755]='h00003eb0;  wr_data_rom[13755]='h00002c60;
    rd_cycle[13756] = 1'b1;  wr_cycle[13756] = 1'b0;  addr_rom[13756]='h00000ed4;  wr_data_rom[13756]='h00000000;
    rd_cycle[13757] = 1'b1;  wr_cycle[13757] = 1'b0;  addr_rom[13757]='h00000924;  wr_data_rom[13757]='h00000000;
    rd_cycle[13758] = 1'b0;  wr_cycle[13758] = 1'b1;  addr_rom[13758]='h000035e8;  wr_data_rom[13758]='h00002e6f;
    rd_cycle[13759] = 1'b1;  wr_cycle[13759] = 1'b0;  addr_rom[13759]='h00002e6c;  wr_data_rom[13759]='h00000000;
    rd_cycle[13760] = 1'b0;  wr_cycle[13760] = 1'b1;  addr_rom[13760]='h00002080;  wr_data_rom[13760]='h000037c8;
    rd_cycle[13761] = 1'b1;  wr_cycle[13761] = 1'b0;  addr_rom[13761]='h000033b0;  wr_data_rom[13761]='h00000000;
    rd_cycle[13762] = 1'b0;  wr_cycle[13762] = 1'b1;  addr_rom[13762]='h00003c80;  wr_data_rom[13762]='h000038c0;
    rd_cycle[13763] = 1'b1;  wr_cycle[13763] = 1'b0;  addr_rom[13763]='h00000628;  wr_data_rom[13763]='h00000000;
    rd_cycle[13764] = 1'b1;  wr_cycle[13764] = 1'b0;  addr_rom[13764]='h00003dc0;  wr_data_rom[13764]='h00000000;
    rd_cycle[13765] = 1'b1;  wr_cycle[13765] = 1'b0;  addr_rom[13765]='h000015fc;  wr_data_rom[13765]='h00000000;
    rd_cycle[13766] = 1'b1;  wr_cycle[13766] = 1'b0;  addr_rom[13766]='h00001c10;  wr_data_rom[13766]='h00000000;
    rd_cycle[13767] = 1'b1;  wr_cycle[13767] = 1'b0;  addr_rom[13767]='h000030f8;  wr_data_rom[13767]='h00000000;
    rd_cycle[13768] = 1'b0;  wr_cycle[13768] = 1'b1;  addr_rom[13768]='h0000106c;  wr_data_rom[13768]='h00002920;
    rd_cycle[13769] = 1'b0;  wr_cycle[13769] = 1'b1;  addr_rom[13769]='h00000bb4;  wr_data_rom[13769]='h00003b85;
    rd_cycle[13770] = 1'b1;  wr_cycle[13770] = 1'b0;  addr_rom[13770]='h000033dc;  wr_data_rom[13770]='h00000000;
    rd_cycle[13771] = 1'b1;  wr_cycle[13771] = 1'b0;  addr_rom[13771]='h0000105c;  wr_data_rom[13771]='h00000000;
    rd_cycle[13772] = 1'b0;  wr_cycle[13772] = 1'b1;  addr_rom[13772]='h00000e50;  wr_data_rom[13772]='h0000196d;
    rd_cycle[13773] = 1'b0;  wr_cycle[13773] = 1'b1;  addr_rom[13773]='h00000e98;  wr_data_rom[13773]='h0000301d;
    rd_cycle[13774] = 1'b0;  wr_cycle[13774] = 1'b1;  addr_rom[13774]='h0000241c;  wr_data_rom[13774]='h0000099f;
    rd_cycle[13775] = 1'b1;  wr_cycle[13775] = 1'b0;  addr_rom[13775]='h000013ac;  wr_data_rom[13775]='h00000000;
    rd_cycle[13776] = 1'b0;  wr_cycle[13776] = 1'b1;  addr_rom[13776]='h000032cc;  wr_data_rom[13776]='h00000f19;
    rd_cycle[13777] = 1'b0;  wr_cycle[13777] = 1'b1;  addr_rom[13777]='h00002b18;  wr_data_rom[13777]='h00000bda;
    rd_cycle[13778] = 1'b0;  wr_cycle[13778] = 1'b1;  addr_rom[13778]='h00002578;  wr_data_rom[13778]='h00000a9b;
    rd_cycle[13779] = 1'b0;  wr_cycle[13779] = 1'b1;  addr_rom[13779]='h00002e0c;  wr_data_rom[13779]='h00000377;
    rd_cycle[13780] = 1'b0;  wr_cycle[13780] = 1'b1;  addr_rom[13780]='h00002ed4;  wr_data_rom[13780]='h00001573;
    rd_cycle[13781] = 1'b1;  wr_cycle[13781] = 1'b0;  addr_rom[13781]='h00000344;  wr_data_rom[13781]='h00000000;
    rd_cycle[13782] = 1'b0;  wr_cycle[13782] = 1'b1;  addr_rom[13782]='h0000058c;  wr_data_rom[13782]='h00002000;
    rd_cycle[13783] = 1'b0;  wr_cycle[13783] = 1'b1;  addr_rom[13783]='h0000007c;  wr_data_rom[13783]='h000020a1;
    rd_cycle[13784] = 1'b1;  wr_cycle[13784] = 1'b0;  addr_rom[13784]='h00002de8;  wr_data_rom[13784]='h00000000;
    rd_cycle[13785] = 1'b1;  wr_cycle[13785] = 1'b0;  addr_rom[13785]='h00001e94;  wr_data_rom[13785]='h00000000;
    rd_cycle[13786] = 1'b0;  wr_cycle[13786] = 1'b1;  addr_rom[13786]='h00003588;  wr_data_rom[13786]='h00001e3a;
    rd_cycle[13787] = 1'b0;  wr_cycle[13787] = 1'b1;  addr_rom[13787]='h00001154;  wr_data_rom[13787]='h00002ced;
    rd_cycle[13788] = 1'b1;  wr_cycle[13788] = 1'b0;  addr_rom[13788]='h000010f8;  wr_data_rom[13788]='h00000000;
    rd_cycle[13789] = 1'b1;  wr_cycle[13789] = 1'b0;  addr_rom[13789]='h000025a4;  wr_data_rom[13789]='h00000000;
    rd_cycle[13790] = 1'b1;  wr_cycle[13790] = 1'b0;  addr_rom[13790]='h000015a8;  wr_data_rom[13790]='h00000000;
    rd_cycle[13791] = 1'b1;  wr_cycle[13791] = 1'b0;  addr_rom[13791]='h00000398;  wr_data_rom[13791]='h00000000;
    rd_cycle[13792] = 1'b1;  wr_cycle[13792] = 1'b0;  addr_rom[13792]='h0000093c;  wr_data_rom[13792]='h00000000;
    rd_cycle[13793] = 1'b0;  wr_cycle[13793] = 1'b1;  addr_rom[13793]='h00002f00;  wr_data_rom[13793]='h0000004e;
    rd_cycle[13794] = 1'b1;  wr_cycle[13794] = 1'b0;  addr_rom[13794]='h00001ec8;  wr_data_rom[13794]='h00000000;
    rd_cycle[13795] = 1'b1;  wr_cycle[13795] = 1'b0;  addr_rom[13795]='h00003cd8;  wr_data_rom[13795]='h00000000;
    rd_cycle[13796] = 1'b1;  wr_cycle[13796] = 1'b0;  addr_rom[13796]='h00000c54;  wr_data_rom[13796]='h00000000;
    rd_cycle[13797] = 1'b1;  wr_cycle[13797] = 1'b0;  addr_rom[13797]='h00000438;  wr_data_rom[13797]='h00000000;
    rd_cycle[13798] = 1'b0;  wr_cycle[13798] = 1'b1;  addr_rom[13798]='h0000217c;  wr_data_rom[13798]='h00001e01;
    rd_cycle[13799] = 1'b1;  wr_cycle[13799] = 1'b0;  addr_rom[13799]='h00001b64;  wr_data_rom[13799]='h00000000;
    rd_cycle[13800] = 1'b0;  wr_cycle[13800] = 1'b1;  addr_rom[13800]='h00002a50;  wr_data_rom[13800]='h00003b9a;
    rd_cycle[13801] = 1'b1;  wr_cycle[13801] = 1'b0;  addr_rom[13801]='h00002d50;  wr_data_rom[13801]='h00000000;
    rd_cycle[13802] = 1'b1;  wr_cycle[13802] = 1'b0;  addr_rom[13802]='h00000018;  wr_data_rom[13802]='h00000000;
    rd_cycle[13803] = 1'b1;  wr_cycle[13803] = 1'b0;  addr_rom[13803]='h00003df4;  wr_data_rom[13803]='h00000000;
    rd_cycle[13804] = 1'b1;  wr_cycle[13804] = 1'b0;  addr_rom[13804]='h00003d5c;  wr_data_rom[13804]='h00000000;
    rd_cycle[13805] = 1'b0;  wr_cycle[13805] = 1'b1;  addr_rom[13805]='h00002b68;  wr_data_rom[13805]='h00001238;
    rd_cycle[13806] = 1'b0;  wr_cycle[13806] = 1'b1;  addr_rom[13806]='h00001ca0;  wr_data_rom[13806]='h00002684;
    rd_cycle[13807] = 1'b1;  wr_cycle[13807] = 1'b0;  addr_rom[13807]='h00002898;  wr_data_rom[13807]='h00000000;
    rd_cycle[13808] = 1'b0;  wr_cycle[13808] = 1'b1;  addr_rom[13808]='h00002ad4;  wr_data_rom[13808]='h00002974;
    rd_cycle[13809] = 1'b1;  wr_cycle[13809] = 1'b0;  addr_rom[13809]='h00003b00;  wr_data_rom[13809]='h00000000;
    rd_cycle[13810] = 1'b1;  wr_cycle[13810] = 1'b0;  addr_rom[13810]='h00003358;  wr_data_rom[13810]='h00000000;
    rd_cycle[13811] = 1'b1;  wr_cycle[13811] = 1'b0;  addr_rom[13811]='h0000190c;  wr_data_rom[13811]='h00000000;
    rd_cycle[13812] = 1'b0;  wr_cycle[13812] = 1'b1;  addr_rom[13812]='h00003f74;  wr_data_rom[13812]='h000000fc;
    rd_cycle[13813] = 1'b1;  wr_cycle[13813] = 1'b0;  addr_rom[13813]='h00003514;  wr_data_rom[13813]='h00000000;
    rd_cycle[13814] = 1'b1;  wr_cycle[13814] = 1'b0;  addr_rom[13814]='h00000078;  wr_data_rom[13814]='h00000000;
    rd_cycle[13815] = 1'b1;  wr_cycle[13815] = 1'b0;  addr_rom[13815]='h00001268;  wr_data_rom[13815]='h00000000;
    rd_cycle[13816] = 1'b0;  wr_cycle[13816] = 1'b1;  addr_rom[13816]='h00003c34;  wr_data_rom[13816]='h00000061;
    rd_cycle[13817] = 1'b1;  wr_cycle[13817] = 1'b0;  addr_rom[13817]='h000002bc;  wr_data_rom[13817]='h00000000;
    rd_cycle[13818] = 1'b1;  wr_cycle[13818] = 1'b0;  addr_rom[13818]='h000004d8;  wr_data_rom[13818]='h00000000;
    rd_cycle[13819] = 1'b1;  wr_cycle[13819] = 1'b0;  addr_rom[13819]='h00001c20;  wr_data_rom[13819]='h00000000;
    rd_cycle[13820] = 1'b0;  wr_cycle[13820] = 1'b1;  addr_rom[13820]='h000033a4;  wr_data_rom[13820]='h000034f9;
    rd_cycle[13821] = 1'b0;  wr_cycle[13821] = 1'b1;  addr_rom[13821]='h0000028c;  wr_data_rom[13821]='h0000013d;
    rd_cycle[13822] = 1'b1;  wr_cycle[13822] = 1'b0;  addr_rom[13822]='h00002b30;  wr_data_rom[13822]='h00000000;
    rd_cycle[13823] = 1'b0;  wr_cycle[13823] = 1'b1;  addr_rom[13823]='h000023c4;  wr_data_rom[13823]='h0000241a;
    rd_cycle[13824] = 1'b0;  wr_cycle[13824] = 1'b1;  addr_rom[13824]='h00000610;  wr_data_rom[13824]='h00000fb2;
    rd_cycle[13825] = 1'b0;  wr_cycle[13825] = 1'b1;  addr_rom[13825]='h00003108;  wr_data_rom[13825]='h00000daf;
    rd_cycle[13826] = 1'b0;  wr_cycle[13826] = 1'b1;  addr_rom[13826]='h0000079c;  wr_data_rom[13826]='h00003b4c;
    rd_cycle[13827] = 1'b0;  wr_cycle[13827] = 1'b1;  addr_rom[13827]='h00000354;  wr_data_rom[13827]='h00000933;
    rd_cycle[13828] = 1'b0;  wr_cycle[13828] = 1'b1;  addr_rom[13828]='h00002650;  wr_data_rom[13828]='h00001863;
    rd_cycle[13829] = 1'b0;  wr_cycle[13829] = 1'b1;  addr_rom[13829]='h000030a0;  wr_data_rom[13829]='h000009d0;
    rd_cycle[13830] = 1'b0;  wr_cycle[13830] = 1'b1;  addr_rom[13830]='h00003550;  wr_data_rom[13830]='h00002fe8;
    rd_cycle[13831] = 1'b0;  wr_cycle[13831] = 1'b1;  addr_rom[13831]='h0000387c;  wr_data_rom[13831]='h00000b7c;
    rd_cycle[13832] = 1'b1;  wr_cycle[13832] = 1'b0;  addr_rom[13832]='h00002f44;  wr_data_rom[13832]='h00000000;
    rd_cycle[13833] = 1'b0;  wr_cycle[13833] = 1'b1;  addr_rom[13833]='h00001df4;  wr_data_rom[13833]='h00003329;
    rd_cycle[13834] = 1'b1;  wr_cycle[13834] = 1'b0;  addr_rom[13834]='h00001dec;  wr_data_rom[13834]='h00000000;
    rd_cycle[13835] = 1'b0;  wr_cycle[13835] = 1'b1;  addr_rom[13835]='h00001218;  wr_data_rom[13835]='h00001d0e;
    rd_cycle[13836] = 1'b0;  wr_cycle[13836] = 1'b1;  addr_rom[13836]='h00000210;  wr_data_rom[13836]='h00003b74;
    rd_cycle[13837] = 1'b1;  wr_cycle[13837] = 1'b0;  addr_rom[13837]='h0000237c;  wr_data_rom[13837]='h00000000;
    rd_cycle[13838] = 1'b1;  wr_cycle[13838] = 1'b0;  addr_rom[13838]='h00001ca4;  wr_data_rom[13838]='h00000000;
    rd_cycle[13839] = 1'b1;  wr_cycle[13839] = 1'b0;  addr_rom[13839]='h0000232c;  wr_data_rom[13839]='h00000000;
    rd_cycle[13840] = 1'b0;  wr_cycle[13840] = 1'b1;  addr_rom[13840]='h0000013c;  wr_data_rom[13840]='h00001f3e;
    rd_cycle[13841] = 1'b1;  wr_cycle[13841] = 1'b0;  addr_rom[13841]='h00003078;  wr_data_rom[13841]='h00000000;
    rd_cycle[13842] = 1'b0;  wr_cycle[13842] = 1'b1;  addr_rom[13842]='h00000a88;  wr_data_rom[13842]='h00000d98;
    rd_cycle[13843] = 1'b1;  wr_cycle[13843] = 1'b0;  addr_rom[13843]='h000033f0;  wr_data_rom[13843]='h00000000;
    rd_cycle[13844] = 1'b1;  wr_cycle[13844] = 1'b0;  addr_rom[13844]='h0000160c;  wr_data_rom[13844]='h00000000;
    rd_cycle[13845] = 1'b1;  wr_cycle[13845] = 1'b0;  addr_rom[13845]='h00002dd4;  wr_data_rom[13845]='h00000000;
    rd_cycle[13846] = 1'b0;  wr_cycle[13846] = 1'b1;  addr_rom[13846]='h00001320;  wr_data_rom[13846]='h000034ee;
    rd_cycle[13847] = 1'b1;  wr_cycle[13847] = 1'b0;  addr_rom[13847]='h00003ad4;  wr_data_rom[13847]='h00000000;
    rd_cycle[13848] = 1'b0;  wr_cycle[13848] = 1'b1;  addr_rom[13848]='h00003148;  wr_data_rom[13848]='h00003e2a;
    rd_cycle[13849] = 1'b0;  wr_cycle[13849] = 1'b1;  addr_rom[13849]='h000015bc;  wr_data_rom[13849]='h00003354;
    rd_cycle[13850] = 1'b1;  wr_cycle[13850] = 1'b0;  addr_rom[13850]='h000000e0;  wr_data_rom[13850]='h00000000;
    rd_cycle[13851] = 1'b1;  wr_cycle[13851] = 1'b0;  addr_rom[13851]='h000025a4;  wr_data_rom[13851]='h00000000;
    rd_cycle[13852] = 1'b0;  wr_cycle[13852] = 1'b1;  addr_rom[13852]='h00000ab4;  wr_data_rom[13852]='h00002561;
    rd_cycle[13853] = 1'b0;  wr_cycle[13853] = 1'b1;  addr_rom[13853]='h00000f28;  wr_data_rom[13853]='h000029b4;
    rd_cycle[13854] = 1'b0;  wr_cycle[13854] = 1'b1;  addr_rom[13854]='h00002e24;  wr_data_rom[13854]='h0000255a;
    rd_cycle[13855] = 1'b1;  wr_cycle[13855] = 1'b0;  addr_rom[13855]='h00002be0;  wr_data_rom[13855]='h00000000;
    rd_cycle[13856] = 1'b1;  wr_cycle[13856] = 1'b0;  addr_rom[13856]='h000028d8;  wr_data_rom[13856]='h00000000;
    rd_cycle[13857] = 1'b0;  wr_cycle[13857] = 1'b1;  addr_rom[13857]='h00001930;  wr_data_rom[13857]='h000004d8;
    rd_cycle[13858] = 1'b0;  wr_cycle[13858] = 1'b1;  addr_rom[13858]='h00002120;  wr_data_rom[13858]='h0000014f;
    rd_cycle[13859] = 1'b1;  wr_cycle[13859] = 1'b0;  addr_rom[13859]='h000000a4;  wr_data_rom[13859]='h00000000;
    rd_cycle[13860] = 1'b1;  wr_cycle[13860] = 1'b0;  addr_rom[13860]='h0000389c;  wr_data_rom[13860]='h00000000;
    rd_cycle[13861] = 1'b1;  wr_cycle[13861] = 1'b0;  addr_rom[13861]='h0000107c;  wr_data_rom[13861]='h00000000;
    rd_cycle[13862] = 1'b1;  wr_cycle[13862] = 1'b0;  addr_rom[13862]='h00001a04;  wr_data_rom[13862]='h00000000;
    rd_cycle[13863] = 1'b1;  wr_cycle[13863] = 1'b0;  addr_rom[13863]='h000026f0;  wr_data_rom[13863]='h00000000;
    rd_cycle[13864] = 1'b1;  wr_cycle[13864] = 1'b0;  addr_rom[13864]='h00001c78;  wr_data_rom[13864]='h00000000;
    rd_cycle[13865] = 1'b1;  wr_cycle[13865] = 1'b0;  addr_rom[13865]='h00001940;  wr_data_rom[13865]='h00000000;
    rd_cycle[13866] = 1'b0;  wr_cycle[13866] = 1'b1;  addr_rom[13866]='h00002d48;  wr_data_rom[13866]='h00003484;
    rd_cycle[13867] = 1'b0;  wr_cycle[13867] = 1'b1;  addr_rom[13867]='h000015c4;  wr_data_rom[13867]='h00001efe;
    rd_cycle[13868] = 1'b0;  wr_cycle[13868] = 1'b1;  addr_rom[13868]='h00001518;  wr_data_rom[13868]='h00003744;
    rd_cycle[13869] = 1'b0;  wr_cycle[13869] = 1'b1;  addr_rom[13869]='h000005f4;  wr_data_rom[13869]='h00001026;
    rd_cycle[13870] = 1'b0;  wr_cycle[13870] = 1'b1;  addr_rom[13870]='h00001784;  wr_data_rom[13870]='h00001d85;
    rd_cycle[13871] = 1'b0;  wr_cycle[13871] = 1'b1;  addr_rom[13871]='h00001464;  wr_data_rom[13871]='h0000144d;
    rd_cycle[13872] = 1'b1;  wr_cycle[13872] = 1'b0;  addr_rom[13872]='h00002498;  wr_data_rom[13872]='h00000000;
    rd_cycle[13873] = 1'b0;  wr_cycle[13873] = 1'b1;  addr_rom[13873]='h00002a50;  wr_data_rom[13873]='h00002ea0;
    rd_cycle[13874] = 1'b1;  wr_cycle[13874] = 1'b0;  addr_rom[13874]='h00001b30;  wr_data_rom[13874]='h00000000;
    rd_cycle[13875] = 1'b1;  wr_cycle[13875] = 1'b0;  addr_rom[13875]='h00002da4;  wr_data_rom[13875]='h00000000;
    rd_cycle[13876] = 1'b1;  wr_cycle[13876] = 1'b0;  addr_rom[13876]='h00001260;  wr_data_rom[13876]='h00000000;
    rd_cycle[13877] = 1'b0;  wr_cycle[13877] = 1'b1;  addr_rom[13877]='h000005bc;  wr_data_rom[13877]='h00000917;
    rd_cycle[13878] = 1'b1;  wr_cycle[13878] = 1'b0;  addr_rom[13878]='h000011b0;  wr_data_rom[13878]='h00000000;
    rd_cycle[13879] = 1'b1;  wr_cycle[13879] = 1'b0;  addr_rom[13879]='h00000698;  wr_data_rom[13879]='h00000000;
    rd_cycle[13880] = 1'b0;  wr_cycle[13880] = 1'b1;  addr_rom[13880]='h00001384;  wr_data_rom[13880]='h00000b8b;
    rd_cycle[13881] = 1'b1;  wr_cycle[13881] = 1'b0;  addr_rom[13881]='h00003e3c;  wr_data_rom[13881]='h00000000;
    rd_cycle[13882] = 1'b1;  wr_cycle[13882] = 1'b0;  addr_rom[13882]='h00003948;  wr_data_rom[13882]='h00000000;
    rd_cycle[13883] = 1'b1;  wr_cycle[13883] = 1'b0;  addr_rom[13883]='h00001b98;  wr_data_rom[13883]='h00000000;
    rd_cycle[13884] = 1'b1;  wr_cycle[13884] = 1'b0;  addr_rom[13884]='h00002d9c;  wr_data_rom[13884]='h00000000;
    rd_cycle[13885] = 1'b1;  wr_cycle[13885] = 1'b0;  addr_rom[13885]='h00003008;  wr_data_rom[13885]='h00000000;
    rd_cycle[13886] = 1'b1;  wr_cycle[13886] = 1'b0;  addr_rom[13886]='h0000056c;  wr_data_rom[13886]='h00000000;
    rd_cycle[13887] = 1'b1;  wr_cycle[13887] = 1'b0;  addr_rom[13887]='h0000038c;  wr_data_rom[13887]='h00000000;
    rd_cycle[13888] = 1'b1;  wr_cycle[13888] = 1'b0;  addr_rom[13888]='h00001980;  wr_data_rom[13888]='h00000000;
    rd_cycle[13889] = 1'b1;  wr_cycle[13889] = 1'b0;  addr_rom[13889]='h00003584;  wr_data_rom[13889]='h00000000;
    rd_cycle[13890] = 1'b1;  wr_cycle[13890] = 1'b0;  addr_rom[13890]='h00002f28;  wr_data_rom[13890]='h00000000;
    rd_cycle[13891] = 1'b0;  wr_cycle[13891] = 1'b1;  addr_rom[13891]='h00000ddc;  wr_data_rom[13891]='h000010c3;
    rd_cycle[13892] = 1'b0;  wr_cycle[13892] = 1'b1;  addr_rom[13892]='h00000ec0;  wr_data_rom[13892]='h000021eb;
    rd_cycle[13893] = 1'b1;  wr_cycle[13893] = 1'b0;  addr_rom[13893]='h00000788;  wr_data_rom[13893]='h00000000;
    rd_cycle[13894] = 1'b1;  wr_cycle[13894] = 1'b0;  addr_rom[13894]='h0000335c;  wr_data_rom[13894]='h00000000;
    rd_cycle[13895] = 1'b1;  wr_cycle[13895] = 1'b0;  addr_rom[13895]='h00001a1c;  wr_data_rom[13895]='h00000000;
    rd_cycle[13896] = 1'b0;  wr_cycle[13896] = 1'b1;  addr_rom[13896]='h000016b4;  wr_data_rom[13896]='h00001bca;
    rd_cycle[13897] = 1'b1;  wr_cycle[13897] = 1'b0;  addr_rom[13897]='h0000250c;  wr_data_rom[13897]='h00000000;
    rd_cycle[13898] = 1'b0;  wr_cycle[13898] = 1'b1;  addr_rom[13898]='h000021ac;  wr_data_rom[13898]='h00003595;
    rd_cycle[13899] = 1'b0;  wr_cycle[13899] = 1'b1;  addr_rom[13899]='h00003284;  wr_data_rom[13899]='h000035d6;
    rd_cycle[13900] = 1'b0;  wr_cycle[13900] = 1'b1;  addr_rom[13900]='h00003484;  wr_data_rom[13900]='h00000245;
    rd_cycle[13901] = 1'b0;  wr_cycle[13901] = 1'b1;  addr_rom[13901]='h00001c48;  wr_data_rom[13901]='h00003a13;
    rd_cycle[13902] = 1'b0;  wr_cycle[13902] = 1'b1;  addr_rom[13902]='h00003e80;  wr_data_rom[13902]='h00003eba;
    rd_cycle[13903] = 1'b0;  wr_cycle[13903] = 1'b1;  addr_rom[13903]='h00001cb4;  wr_data_rom[13903]='h0000213b;
    rd_cycle[13904] = 1'b1;  wr_cycle[13904] = 1'b0;  addr_rom[13904]='h00001bb0;  wr_data_rom[13904]='h00000000;
    rd_cycle[13905] = 1'b0;  wr_cycle[13905] = 1'b1;  addr_rom[13905]='h00000d50;  wr_data_rom[13905]='h000003e3;
    rd_cycle[13906] = 1'b1;  wr_cycle[13906] = 1'b0;  addr_rom[13906]='h00003e94;  wr_data_rom[13906]='h00000000;
    rd_cycle[13907] = 1'b1;  wr_cycle[13907] = 1'b0;  addr_rom[13907]='h00003e98;  wr_data_rom[13907]='h00000000;
    rd_cycle[13908] = 1'b0;  wr_cycle[13908] = 1'b1;  addr_rom[13908]='h00000228;  wr_data_rom[13908]='h00001875;
    rd_cycle[13909] = 1'b1;  wr_cycle[13909] = 1'b0;  addr_rom[13909]='h000034e4;  wr_data_rom[13909]='h00000000;
    rd_cycle[13910] = 1'b0;  wr_cycle[13910] = 1'b1;  addr_rom[13910]='h000010b8;  wr_data_rom[13910]='h0000006d;
    rd_cycle[13911] = 1'b1;  wr_cycle[13911] = 1'b0;  addr_rom[13911]='h00001fbc;  wr_data_rom[13911]='h00000000;
    rd_cycle[13912] = 1'b0;  wr_cycle[13912] = 1'b1;  addr_rom[13912]='h00001d04;  wr_data_rom[13912]='h0000163b;
    rd_cycle[13913] = 1'b1;  wr_cycle[13913] = 1'b0;  addr_rom[13913]='h000004b8;  wr_data_rom[13913]='h00000000;
    rd_cycle[13914] = 1'b1;  wr_cycle[13914] = 1'b0;  addr_rom[13914]='h00003274;  wr_data_rom[13914]='h00000000;
    rd_cycle[13915] = 1'b0;  wr_cycle[13915] = 1'b1;  addr_rom[13915]='h000010a0;  wr_data_rom[13915]='h0000381f;
    rd_cycle[13916] = 1'b1;  wr_cycle[13916] = 1'b0;  addr_rom[13916]='h00002658;  wr_data_rom[13916]='h00000000;
    rd_cycle[13917] = 1'b0;  wr_cycle[13917] = 1'b1;  addr_rom[13917]='h000034a4;  wr_data_rom[13917]='h000017f2;
    rd_cycle[13918] = 1'b0;  wr_cycle[13918] = 1'b1;  addr_rom[13918]='h000026bc;  wr_data_rom[13918]='h00000a01;
    rd_cycle[13919] = 1'b1;  wr_cycle[13919] = 1'b0;  addr_rom[13919]='h00001ef8;  wr_data_rom[13919]='h00000000;
    rd_cycle[13920] = 1'b1;  wr_cycle[13920] = 1'b0;  addr_rom[13920]='h000031c8;  wr_data_rom[13920]='h00000000;
    rd_cycle[13921] = 1'b1;  wr_cycle[13921] = 1'b0;  addr_rom[13921]='h000032a8;  wr_data_rom[13921]='h00000000;
    rd_cycle[13922] = 1'b0;  wr_cycle[13922] = 1'b1;  addr_rom[13922]='h0000228c;  wr_data_rom[13922]='h00000d24;
    rd_cycle[13923] = 1'b0;  wr_cycle[13923] = 1'b1;  addr_rom[13923]='h00001168;  wr_data_rom[13923]='h000002d1;
    rd_cycle[13924] = 1'b1;  wr_cycle[13924] = 1'b0;  addr_rom[13924]='h0000396c;  wr_data_rom[13924]='h00000000;
    rd_cycle[13925] = 1'b1;  wr_cycle[13925] = 1'b0;  addr_rom[13925]='h00000d98;  wr_data_rom[13925]='h00000000;
    rd_cycle[13926] = 1'b1;  wr_cycle[13926] = 1'b0;  addr_rom[13926]='h000004c8;  wr_data_rom[13926]='h00000000;
    rd_cycle[13927] = 1'b0;  wr_cycle[13927] = 1'b1;  addr_rom[13927]='h00001978;  wr_data_rom[13927]='h000036ef;
    rd_cycle[13928] = 1'b1;  wr_cycle[13928] = 1'b0;  addr_rom[13928]='h000007c0;  wr_data_rom[13928]='h00000000;
    rd_cycle[13929] = 1'b1;  wr_cycle[13929] = 1'b0;  addr_rom[13929]='h00003310;  wr_data_rom[13929]='h00000000;
    rd_cycle[13930] = 1'b1;  wr_cycle[13930] = 1'b0;  addr_rom[13930]='h00002770;  wr_data_rom[13930]='h00000000;
    rd_cycle[13931] = 1'b1;  wr_cycle[13931] = 1'b0;  addr_rom[13931]='h000027c0;  wr_data_rom[13931]='h00000000;
    rd_cycle[13932] = 1'b1;  wr_cycle[13932] = 1'b0;  addr_rom[13932]='h0000343c;  wr_data_rom[13932]='h00000000;
    rd_cycle[13933] = 1'b0;  wr_cycle[13933] = 1'b1;  addr_rom[13933]='h00001a2c;  wr_data_rom[13933]='h00002a86;
    rd_cycle[13934] = 1'b1;  wr_cycle[13934] = 1'b0;  addr_rom[13934]='h000022f4;  wr_data_rom[13934]='h00000000;
    rd_cycle[13935] = 1'b0;  wr_cycle[13935] = 1'b1;  addr_rom[13935]='h00003eac;  wr_data_rom[13935]='h000020e2;
    rd_cycle[13936] = 1'b0;  wr_cycle[13936] = 1'b1;  addr_rom[13936]='h00000e08;  wr_data_rom[13936]='h00001f9f;
    rd_cycle[13937] = 1'b1;  wr_cycle[13937] = 1'b0;  addr_rom[13937]='h0000328c;  wr_data_rom[13937]='h00000000;
    rd_cycle[13938] = 1'b1;  wr_cycle[13938] = 1'b0;  addr_rom[13938]='h00000274;  wr_data_rom[13938]='h00000000;
    rd_cycle[13939] = 1'b1;  wr_cycle[13939] = 1'b0;  addr_rom[13939]='h00001ce0;  wr_data_rom[13939]='h00000000;
    rd_cycle[13940] = 1'b0;  wr_cycle[13940] = 1'b1;  addr_rom[13940]='h000032d0;  wr_data_rom[13940]='h00002a8a;
    rd_cycle[13941] = 1'b1;  wr_cycle[13941] = 1'b0;  addr_rom[13941]='h000033ec;  wr_data_rom[13941]='h00000000;
    rd_cycle[13942] = 1'b1;  wr_cycle[13942] = 1'b0;  addr_rom[13942]='h00001874;  wr_data_rom[13942]='h00000000;
    rd_cycle[13943] = 1'b1;  wr_cycle[13943] = 1'b0;  addr_rom[13943]='h000008a8;  wr_data_rom[13943]='h00000000;
    rd_cycle[13944] = 1'b1;  wr_cycle[13944] = 1'b0;  addr_rom[13944]='h00003d10;  wr_data_rom[13944]='h00000000;
    rd_cycle[13945] = 1'b1;  wr_cycle[13945] = 1'b0;  addr_rom[13945]='h0000043c;  wr_data_rom[13945]='h00000000;
    rd_cycle[13946] = 1'b0;  wr_cycle[13946] = 1'b1;  addr_rom[13946]='h000017f0;  wr_data_rom[13946]='h00002da5;
    rd_cycle[13947] = 1'b1;  wr_cycle[13947] = 1'b0;  addr_rom[13947]='h00002500;  wr_data_rom[13947]='h00000000;
    rd_cycle[13948] = 1'b0;  wr_cycle[13948] = 1'b1;  addr_rom[13948]='h00001e88;  wr_data_rom[13948]='h0000094a;
    rd_cycle[13949] = 1'b1;  wr_cycle[13949] = 1'b0;  addr_rom[13949]='h00002714;  wr_data_rom[13949]='h00000000;
    rd_cycle[13950] = 1'b1;  wr_cycle[13950] = 1'b0;  addr_rom[13950]='h000020c4;  wr_data_rom[13950]='h00000000;
    rd_cycle[13951] = 1'b1;  wr_cycle[13951] = 1'b0;  addr_rom[13951]='h00000ca0;  wr_data_rom[13951]='h00000000;
    rd_cycle[13952] = 1'b0;  wr_cycle[13952] = 1'b1;  addr_rom[13952]='h00000b34;  wr_data_rom[13952]='h000011fe;
    rd_cycle[13953] = 1'b0;  wr_cycle[13953] = 1'b1;  addr_rom[13953]='h00001d7c;  wr_data_rom[13953]='h00003cc8;
    rd_cycle[13954] = 1'b1;  wr_cycle[13954] = 1'b0;  addr_rom[13954]='h00000ca4;  wr_data_rom[13954]='h00000000;
    rd_cycle[13955] = 1'b0;  wr_cycle[13955] = 1'b1;  addr_rom[13955]='h00000d28;  wr_data_rom[13955]='h0000344b;
    rd_cycle[13956] = 1'b0;  wr_cycle[13956] = 1'b1;  addr_rom[13956]='h00000ef8;  wr_data_rom[13956]='h0000093a;
    rd_cycle[13957] = 1'b1;  wr_cycle[13957] = 1'b0;  addr_rom[13957]='h00000210;  wr_data_rom[13957]='h00000000;
    rd_cycle[13958] = 1'b1;  wr_cycle[13958] = 1'b0;  addr_rom[13958]='h000023d4;  wr_data_rom[13958]='h00000000;
    rd_cycle[13959] = 1'b1;  wr_cycle[13959] = 1'b0;  addr_rom[13959]='h0000374c;  wr_data_rom[13959]='h00000000;
    rd_cycle[13960] = 1'b0;  wr_cycle[13960] = 1'b1;  addr_rom[13960]='h00001398;  wr_data_rom[13960]='h000019b9;
    rd_cycle[13961] = 1'b1;  wr_cycle[13961] = 1'b0;  addr_rom[13961]='h00000df8;  wr_data_rom[13961]='h00000000;
    rd_cycle[13962] = 1'b1;  wr_cycle[13962] = 1'b0;  addr_rom[13962]='h00002824;  wr_data_rom[13962]='h00000000;
    rd_cycle[13963] = 1'b0;  wr_cycle[13963] = 1'b1;  addr_rom[13963]='h000011a0;  wr_data_rom[13963]='h000035a6;
    rd_cycle[13964] = 1'b1;  wr_cycle[13964] = 1'b0;  addr_rom[13964]='h00003970;  wr_data_rom[13964]='h00000000;
    rd_cycle[13965] = 1'b0;  wr_cycle[13965] = 1'b1;  addr_rom[13965]='h000028b8;  wr_data_rom[13965]='h0000349d;
    rd_cycle[13966] = 1'b0;  wr_cycle[13966] = 1'b1;  addr_rom[13966]='h000005d8;  wr_data_rom[13966]='h00000203;
    rd_cycle[13967] = 1'b1;  wr_cycle[13967] = 1'b0;  addr_rom[13967]='h00003144;  wr_data_rom[13967]='h00000000;
    rd_cycle[13968] = 1'b0;  wr_cycle[13968] = 1'b1;  addr_rom[13968]='h00000e74;  wr_data_rom[13968]='h0000354b;
    rd_cycle[13969] = 1'b0;  wr_cycle[13969] = 1'b1;  addr_rom[13969]='h000035ec;  wr_data_rom[13969]='h0000075c;
    rd_cycle[13970] = 1'b1;  wr_cycle[13970] = 1'b0;  addr_rom[13970]='h0000183c;  wr_data_rom[13970]='h00000000;
    rd_cycle[13971] = 1'b1;  wr_cycle[13971] = 1'b0;  addr_rom[13971]='h00003928;  wr_data_rom[13971]='h00000000;
    rd_cycle[13972] = 1'b1;  wr_cycle[13972] = 1'b0;  addr_rom[13972]='h0000357c;  wr_data_rom[13972]='h00000000;
    rd_cycle[13973] = 1'b1;  wr_cycle[13973] = 1'b0;  addr_rom[13973]='h00001fe8;  wr_data_rom[13973]='h00000000;
    rd_cycle[13974] = 1'b0;  wr_cycle[13974] = 1'b1;  addr_rom[13974]='h00001f3c;  wr_data_rom[13974]='h000011eb;
    rd_cycle[13975] = 1'b1;  wr_cycle[13975] = 1'b0;  addr_rom[13975]='h000037cc;  wr_data_rom[13975]='h00000000;
    rd_cycle[13976] = 1'b1;  wr_cycle[13976] = 1'b0;  addr_rom[13976]='h00001478;  wr_data_rom[13976]='h00000000;
    rd_cycle[13977] = 1'b0;  wr_cycle[13977] = 1'b1;  addr_rom[13977]='h00003ec0;  wr_data_rom[13977]='h000037ab;
    rd_cycle[13978] = 1'b0;  wr_cycle[13978] = 1'b1;  addr_rom[13978]='h000012c8;  wr_data_rom[13978]='h00003d36;
    rd_cycle[13979] = 1'b1;  wr_cycle[13979] = 1'b0;  addr_rom[13979]='h0000315c;  wr_data_rom[13979]='h00000000;
    rd_cycle[13980] = 1'b1;  wr_cycle[13980] = 1'b0;  addr_rom[13980]='h00000644;  wr_data_rom[13980]='h00000000;
    rd_cycle[13981] = 1'b0;  wr_cycle[13981] = 1'b1;  addr_rom[13981]='h000003c4;  wr_data_rom[13981]='h0000396b;
    rd_cycle[13982] = 1'b0;  wr_cycle[13982] = 1'b1;  addr_rom[13982]='h00003520;  wr_data_rom[13982]='h000034cc;
    rd_cycle[13983] = 1'b0;  wr_cycle[13983] = 1'b1;  addr_rom[13983]='h00002fd4;  wr_data_rom[13983]='h0000070a;
    rd_cycle[13984] = 1'b1;  wr_cycle[13984] = 1'b0;  addr_rom[13984]='h00000e9c;  wr_data_rom[13984]='h00000000;
    rd_cycle[13985] = 1'b1;  wr_cycle[13985] = 1'b0;  addr_rom[13985]='h000012f0;  wr_data_rom[13985]='h00000000;
    rd_cycle[13986] = 1'b1;  wr_cycle[13986] = 1'b0;  addr_rom[13986]='h00003848;  wr_data_rom[13986]='h00000000;
    rd_cycle[13987] = 1'b1;  wr_cycle[13987] = 1'b0;  addr_rom[13987]='h00000c1c;  wr_data_rom[13987]='h00000000;
    rd_cycle[13988] = 1'b0;  wr_cycle[13988] = 1'b1;  addr_rom[13988]='h000011b0;  wr_data_rom[13988]='h00000a7f;
    rd_cycle[13989] = 1'b0;  wr_cycle[13989] = 1'b1;  addr_rom[13989]='h00002a00;  wr_data_rom[13989]='h000012ef;
    rd_cycle[13990] = 1'b1;  wr_cycle[13990] = 1'b0;  addr_rom[13990]='h00003cdc;  wr_data_rom[13990]='h00000000;
    rd_cycle[13991] = 1'b1;  wr_cycle[13991] = 1'b0;  addr_rom[13991]='h00000178;  wr_data_rom[13991]='h00000000;
    rd_cycle[13992] = 1'b0;  wr_cycle[13992] = 1'b1;  addr_rom[13992]='h00003b3c;  wr_data_rom[13992]='h00002a18;
    rd_cycle[13993] = 1'b0;  wr_cycle[13993] = 1'b1;  addr_rom[13993]='h000039a8;  wr_data_rom[13993]='h000002d3;
    rd_cycle[13994] = 1'b0;  wr_cycle[13994] = 1'b1;  addr_rom[13994]='h00003238;  wr_data_rom[13994]='h00002be9;
    rd_cycle[13995] = 1'b1;  wr_cycle[13995] = 1'b0;  addr_rom[13995]='h00001490;  wr_data_rom[13995]='h00000000;
    rd_cycle[13996] = 1'b1;  wr_cycle[13996] = 1'b0;  addr_rom[13996]='h000005ec;  wr_data_rom[13996]='h00000000;
    rd_cycle[13997] = 1'b1;  wr_cycle[13997] = 1'b0;  addr_rom[13997]='h00003590;  wr_data_rom[13997]='h00000000;
    rd_cycle[13998] = 1'b1;  wr_cycle[13998] = 1'b0;  addr_rom[13998]='h00002ebc;  wr_data_rom[13998]='h00000000;
    rd_cycle[13999] = 1'b1;  wr_cycle[13999] = 1'b0;  addr_rom[13999]='h00002c24;  wr_data_rom[13999]='h00000000;
    rd_cycle[14000] = 1'b1;  wr_cycle[14000] = 1'b0;  addr_rom[14000]='h00001adc;  wr_data_rom[14000]='h00000000;
    rd_cycle[14001] = 1'b0;  wr_cycle[14001] = 1'b1;  addr_rom[14001]='h0000269c;  wr_data_rom[14001]='h000024cb;
    rd_cycle[14002] = 1'b0;  wr_cycle[14002] = 1'b1;  addr_rom[14002]='h00002178;  wr_data_rom[14002]='h00003a91;
    rd_cycle[14003] = 1'b0;  wr_cycle[14003] = 1'b1;  addr_rom[14003]='h00001fbc;  wr_data_rom[14003]='h000013d8;
    rd_cycle[14004] = 1'b0;  wr_cycle[14004] = 1'b1;  addr_rom[14004]='h000017c4;  wr_data_rom[14004]='h000007ce;
    rd_cycle[14005] = 1'b1;  wr_cycle[14005] = 1'b0;  addr_rom[14005]='h00000a6c;  wr_data_rom[14005]='h00000000;
    rd_cycle[14006] = 1'b1;  wr_cycle[14006] = 1'b0;  addr_rom[14006]='h000020ac;  wr_data_rom[14006]='h00000000;
    rd_cycle[14007] = 1'b1;  wr_cycle[14007] = 1'b0;  addr_rom[14007]='h0000103c;  wr_data_rom[14007]='h00000000;
    rd_cycle[14008] = 1'b1;  wr_cycle[14008] = 1'b0;  addr_rom[14008]='h00003e3c;  wr_data_rom[14008]='h00000000;
    rd_cycle[14009] = 1'b0;  wr_cycle[14009] = 1'b1;  addr_rom[14009]='h000018b4;  wr_data_rom[14009]='h00000e0f;
    rd_cycle[14010] = 1'b1;  wr_cycle[14010] = 1'b0;  addr_rom[14010]='h00003d4c;  wr_data_rom[14010]='h00000000;
    rd_cycle[14011] = 1'b1;  wr_cycle[14011] = 1'b0;  addr_rom[14011]='h000036f4;  wr_data_rom[14011]='h00000000;
    rd_cycle[14012] = 1'b1;  wr_cycle[14012] = 1'b0;  addr_rom[14012]='h00001adc;  wr_data_rom[14012]='h00000000;
    rd_cycle[14013] = 1'b0;  wr_cycle[14013] = 1'b1;  addr_rom[14013]='h000009cc;  wr_data_rom[14013]='h0000218e;
    rd_cycle[14014] = 1'b0;  wr_cycle[14014] = 1'b1;  addr_rom[14014]='h00003678;  wr_data_rom[14014]='h0000203a;
    rd_cycle[14015] = 1'b0;  wr_cycle[14015] = 1'b1;  addr_rom[14015]='h000032a0;  wr_data_rom[14015]='h000027fa;
    rd_cycle[14016] = 1'b1;  wr_cycle[14016] = 1'b0;  addr_rom[14016]='h00001054;  wr_data_rom[14016]='h00000000;
    rd_cycle[14017] = 1'b1;  wr_cycle[14017] = 1'b0;  addr_rom[14017]='h00003c40;  wr_data_rom[14017]='h00000000;
    rd_cycle[14018] = 1'b1;  wr_cycle[14018] = 1'b0;  addr_rom[14018]='h000000f0;  wr_data_rom[14018]='h00000000;
    rd_cycle[14019] = 1'b1;  wr_cycle[14019] = 1'b0;  addr_rom[14019]='h00000914;  wr_data_rom[14019]='h00000000;
    rd_cycle[14020] = 1'b1;  wr_cycle[14020] = 1'b0;  addr_rom[14020]='h00000764;  wr_data_rom[14020]='h00000000;
    rd_cycle[14021] = 1'b0;  wr_cycle[14021] = 1'b1;  addr_rom[14021]='h00002de0;  wr_data_rom[14021]='h00001860;
    rd_cycle[14022] = 1'b0;  wr_cycle[14022] = 1'b1;  addr_rom[14022]='h000031a4;  wr_data_rom[14022]='h000023d2;
    rd_cycle[14023] = 1'b0;  wr_cycle[14023] = 1'b1;  addr_rom[14023]='h0000076c;  wr_data_rom[14023]='h000038bb;
    rd_cycle[14024] = 1'b1;  wr_cycle[14024] = 1'b0;  addr_rom[14024]='h00000ed8;  wr_data_rom[14024]='h00000000;
    rd_cycle[14025] = 1'b0;  wr_cycle[14025] = 1'b1;  addr_rom[14025]='h00002050;  wr_data_rom[14025]='h00002a0f;
    rd_cycle[14026] = 1'b0;  wr_cycle[14026] = 1'b1;  addr_rom[14026]='h0000049c;  wr_data_rom[14026]='h000009d6;
    rd_cycle[14027] = 1'b0;  wr_cycle[14027] = 1'b1;  addr_rom[14027]='h00003ba4;  wr_data_rom[14027]='h0000065a;
    rd_cycle[14028] = 1'b0;  wr_cycle[14028] = 1'b1;  addr_rom[14028]='h00001860;  wr_data_rom[14028]='h00002be3;
    rd_cycle[14029] = 1'b1;  wr_cycle[14029] = 1'b0;  addr_rom[14029]='h000025f0;  wr_data_rom[14029]='h00000000;
    rd_cycle[14030] = 1'b0;  wr_cycle[14030] = 1'b1;  addr_rom[14030]='h00000ba0;  wr_data_rom[14030]='h0000146c;
    rd_cycle[14031] = 1'b1;  wr_cycle[14031] = 1'b0;  addr_rom[14031]='h000039fc;  wr_data_rom[14031]='h00000000;
    rd_cycle[14032] = 1'b1;  wr_cycle[14032] = 1'b0;  addr_rom[14032]='h00001a60;  wr_data_rom[14032]='h00000000;
    rd_cycle[14033] = 1'b0;  wr_cycle[14033] = 1'b1;  addr_rom[14033]='h00003720;  wr_data_rom[14033]='h000036fb;
    rd_cycle[14034] = 1'b0;  wr_cycle[14034] = 1'b1;  addr_rom[14034]='h00002e14;  wr_data_rom[14034]='h000001bb;
    rd_cycle[14035] = 1'b1;  wr_cycle[14035] = 1'b0;  addr_rom[14035]='h00002100;  wr_data_rom[14035]='h00000000;
    rd_cycle[14036] = 1'b0;  wr_cycle[14036] = 1'b1;  addr_rom[14036]='h0000299c;  wr_data_rom[14036]='h000008d5;
    rd_cycle[14037] = 1'b1;  wr_cycle[14037] = 1'b0;  addr_rom[14037]='h000035a8;  wr_data_rom[14037]='h00000000;
    rd_cycle[14038] = 1'b0;  wr_cycle[14038] = 1'b1;  addr_rom[14038]='h00003290;  wr_data_rom[14038]='h000024a4;
    rd_cycle[14039] = 1'b1;  wr_cycle[14039] = 1'b0;  addr_rom[14039]='h0000006c;  wr_data_rom[14039]='h00000000;
    rd_cycle[14040] = 1'b1;  wr_cycle[14040] = 1'b0;  addr_rom[14040]='h00002b54;  wr_data_rom[14040]='h00000000;
    rd_cycle[14041] = 1'b0;  wr_cycle[14041] = 1'b1;  addr_rom[14041]='h000006b4;  wr_data_rom[14041]='h00000028;
    rd_cycle[14042] = 1'b1;  wr_cycle[14042] = 1'b0;  addr_rom[14042]='h00001938;  wr_data_rom[14042]='h00000000;
    rd_cycle[14043] = 1'b0;  wr_cycle[14043] = 1'b1;  addr_rom[14043]='h000008e0;  wr_data_rom[14043]='h00003a45;
    rd_cycle[14044] = 1'b1;  wr_cycle[14044] = 1'b0;  addr_rom[14044]='h000027d0;  wr_data_rom[14044]='h00000000;
    rd_cycle[14045] = 1'b1;  wr_cycle[14045] = 1'b0;  addr_rom[14045]='h000028a0;  wr_data_rom[14045]='h00000000;
    rd_cycle[14046] = 1'b1;  wr_cycle[14046] = 1'b0;  addr_rom[14046]='h00002544;  wr_data_rom[14046]='h00000000;
    rd_cycle[14047] = 1'b0;  wr_cycle[14047] = 1'b1;  addr_rom[14047]='h00001648;  wr_data_rom[14047]='h000023e8;
    rd_cycle[14048] = 1'b1;  wr_cycle[14048] = 1'b0;  addr_rom[14048]='h0000292c;  wr_data_rom[14048]='h00000000;
    rd_cycle[14049] = 1'b1;  wr_cycle[14049] = 1'b0;  addr_rom[14049]='h000025bc;  wr_data_rom[14049]='h00000000;
    rd_cycle[14050] = 1'b0;  wr_cycle[14050] = 1'b1;  addr_rom[14050]='h00000854;  wr_data_rom[14050]='h00002b99;
    rd_cycle[14051] = 1'b1;  wr_cycle[14051] = 1'b0;  addr_rom[14051]='h000032ac;  wr_data_rom[14051]='h00000000;
    rd_cycle[14052] = 1'b0;  wr_cycle[14052] = 1'b1;  addr_rom[14052]='h00000a78;  wr_data_rom[14052]='h00001895;
    rd_cycle[14053] = 1'b1;  wr_cycle[14053] = 1'b0;  addr_rom[14053]='h0000071c;  wr_data_rom[14053]='h00000000;
    rd_cycle[14054] = 1'b1;  wr_cycle[14054] = 1'b0;  addr_rom[14054]='h00001a10;  wr_data_rom[14054]='h00000000;
    rd_cycle[14055] = 1'b1;  wr_cycle[14055] = 1'b0;  addr_rom[14055]='h000009e0;  wr_data_rom[14055]='h00000000;
    rd_cycle[14056] = 1'b1;  wr_cycle[14056] = 1'b0;  addr_rom[14056]='h000022fc;  wr_data_rom[14056]='h00000000;
    rd_cycle[14057] = 1'b1;  wr_cycle[14057] = 1'b0;  addr_rom[14057]='h00003374;  wr_data_rom[14057]='h00000000;
    rd_cycle[14058] = 1'b1;  wr_cycle[14058] = 1'b0;  addr_rom[14058]='h00001088;  wr_data_rom[14058]='h00000000;
    rd_cycle[14059] = 1'b0;  wr_cycle[14059] = 1'b1;  addr_rom[14059]='h00003a18;  wr_data_rom[14059]='h00003270;
    rd_cycle[14060] = 1'b1;  wr_cycle[14060] = 1'b0;  addr_rom[14060]='h00001910;  wr_data_rom[14060]='h00000000;
    rd_cycle[14061] = 1'b1;  wr_cycle[14061] = 1'b0;  addr_rom[14061]='h00000d50;  wr_data_rom[14061]='h00000000;
    rd_cycle[14062] = 1'b1;  wr_cycle[14062] = 1'b0;  addr_rom[14062]='h00000408;  wr_data_rom[14062]='h00000000;
    rd_cycle[14063] = 1'b0;  wr_cycle[14063] = 1'b1;  addr_rom[14063]='h00000cf8;  wr_data_rom[14063]='h00000b0c;
    rd_cycle[14064] = 1'b1;  wr_cycle[14064] = 1'b0;  addr_rom[14064]='h00002be4;  wr_data_rom[14064]='h00000000;
    rd_cycle[14065] = 1'b1;  wr_cycle[14065] = 1'b0;  addr_rom[14065]='h00000cc0;  wr_data_rom[14065]='h00000000;
    rd_cycle[14066] = 1'b1;  wr_cycle[14066] = 1'b0;  addr_rom[14066]='h00000488;  wr_data_rom[14066]='h00000000;
    rd_cycle[14067] = 1'b0;  wr_cycle[14067] = 1'b1;  addr_rom[14067]='h00003678;  wr_data_rom[14067]='h00000a3b;
    rd_cycle[14068] = 1'b1;  wr_cycle[14068] = 1'b0;  addr_rom[14068]='h00002ad8;  wr_data_rom[14068]='h00000000;
    rd_cycle[14069] = 1'b0;  wr_cycle[14069] = 1'b1;  addr_rom[14069]='h0000138c;  wr_data_rom[14069]='h00003451;
    rd_cycle[14070] = 1'b0;  wr_cycle[14070] = 1'b1;  addr_rom[14070]='h00003194;  wr_data_rom[14070]='h000035ef;
    rd_cycle[14071] = 1'b0;  wr_cycle[14071] = 1'b1;  addr_rom[14071]='h00001474;  wr_data_rom[14071]='h0000117f;
    rd_cycle[14072] = 1'b0;  wr_cycle[14072] = 1'b1;  addr_rom[14072]='h00001ce0;  wr_data_rom[14072]='h00000f8c;
    rd_cycle[14073] = 1'b1;  wr_cycle[14073] = 1'b0;  addr_rom[14073]='h00001e38;  wr_data_rom[14073]='h00000000;
    rd_cycle[14074] = 1'b0;  wr_cycle[14074] = 1'b1;  addr_rom[14074]='h00003f08;  wr_data_rom[14074]='h00001762;
    rd_cycle[14075] = 1'b0;  wr_cycle[14075] = 1'b1;  addr_rom[14075]='h00001d54;  wr_data_rom[14075]='h000010d3;
    rd_cycle[14076] = 1'b0;  wr_cycle[14076] = 1'b1;  addr_rom[14076]='h00003f20;  wr_data_rom[14076]='h000038eb;
    rd_cycle[14077] = 1'b1;  wr_cycle[14077] = 1'b0;  addr_rom[14077]='h00003654;  wr_data_rom[14077]='h00000000;
    rd_cycle[14078] = 1'b0;  wr_cycle[14078] = 1'b1;  addr_rom[14078]='h00001efc;  wr_data_rom[14078]='h00000c26;
    rd_cycle[14079] = 1'b1;  wr_cycle[14079] = 1'b0;  addr_rom[14079]='h0000305c;  wr_data_rom[14079]='h00000000;
    rd_cycle[14080] = 1'b0;  wr_cycle[14080] = 1'b1;  addr_rom[14080]='h00003fb8;  wr_data_rom[14080]='h00003ac3;
    rd_cycle[14081] = 1'b1;  wr_cycle[14081] = 1'b0;  addr_rom[14081]='h00001ee8;  wr_data_rom[14081]='h00000000;
    rd_cycle[14082] = 1'b0;  wr_cycle[14082] = 1'b1;  addr_rom[14082]='h00001cf8;  wr_data_rom[14082]='h000001f9;
    rd_cycle[14083] = 1'b1;  wr_cycle[14083] = 1'b0;  addr_rom[14083]='h000013ac;  wr_data_rom[14083]='h00000000;
    rd_cycle[14084] = 1'b1;  wr_cycle[14084] = 1'b0;  addr_rom[14084]='h00001eb0;  wr_data_rom[14084]='h00000000;
    rd_cycle[14085] = 1'b0;  wr_cycle[14085] = 1'b1;  addr_rom[14085]='h00003704;  wr_data_rom[14085]='h00003b45;
    rd_cycle[14086] = 1'b0;  wr_cycle[14086] = 1'b1;  addr_rom[14086]='h00002140;  wr_data_rom[14086]='h00002560;
    rd_cycle[14087] = 1'b0;  wr_cycle[14087] = 1'b1;  addr_rom[14087]='h00000860;  wr_data_rom[14087]='h00003493;
    rd_cycle[14088] = 1'b1;  wr_cycle[14088] = 1'b0;  addr_rom[14088]='h0000313c;  wr_data_rom[14088]='h00000000;
    rd_cycle[14089] = 1'b1;  wr_cycle[14089] = 1'b0;  addr_rom[14089]='h00001eb0;  wr_data_rom[14089]='h00000000;
    rd_cycle[14090] = 1'b1;  wr_cycle[14090] = 1'b0;  addr_rom[14090]='h00003d18;  wr_data_rom[14090]='h00000000;
    rd_cycle[14091] = 1'b0;  wr_cycle[14091] = 1'b1;  addr_rom[14091]='h00000bfc;  wr_data_rom[14091]='h0000055e;
    rd_cycle[14092] = 1'b0;  wr_cycle[14092] = 1'b1;  addr_rom[14092]='h00002860;  wr_data_rom[14092]='h00002f94;
    rd_cycle[14093] = 1'b1;  wr_cycle[14093] = 1'b0;  addr_rom[14093]='h00001598;  wr_data_rom[14093]='h00000000;
    rd_cycle[14094] = 1'b1;  wr_cycle[14094] = 1'b0;  addr_rom[14094]='h00001dec;  wr_data_rom[14094]='h00000000;
    rd_cycle[14095] = 1'b0;  wr_cycle[14095] = 1'b1;  addr_rom[14095]='h000000f8;  wr_data_rom[14095]='h00002be5;
    rd_cycle[14096] = 1'b0;  wr_cycle[14096] = 1'b1;  addr_rom[14096]='h00002f7c;  wr_data_rom[14096]='h00002fac;
    rd_cycle[14097] = 1'b0;  wr_cycle[14097] = 1'b1;  addr_rom[14097]='h000024e0;  wr_data_rom[14097]='h00002605;
    rd_cycle[14098] = 1'b1;  wr_cycle[14098] = 1'b0;  addr_rom[14098]='h00003488;  wr_data_rom[14098]='h00000000;
    rd_cycle[14099] = 1'b1;  wr_cycle[14099] = 1'b0;  addr_rom[14099]='h00001c18;  wr_data_rom[14099]='h00000000;
    rd_cycle[14100] = 1'b0;  wr_cycle[14100] = 1'b1;  addr_rom[14100]='h000008bc;  wr_data_rom[14100]='h00000ba9;
    rd_cycle[14101] = 1'b0;  wr_cycle[14101] = 1'b1;  addr_rom[14101]='h0000238c;  wr_data_rom[14101]='h000029b9;
    rd_cycle[14102] = 1'b1;  wr_cycle[14102] = 1'b0;  addr_rom[14102]='h00001fec;  wr_data_rom[14102]='h00000000;
    rd_cycle[14103] = 1'b0;  wr_cycle[14103] = 1'b1;  addr_rom[14103]='h00002ab8;  wr_data_rom[14103]='h0000181d;
    rd_cycle[14104] = 1'b1;  wr_cycle[14104] = 1'b0;  addr_rom[14104]='h00003e48;  wr_data_rom[14104]='h00000000;
    rd_cycle[14105] = 1'b1;  wr_cycle[14105] = 1'b0;  addr_rom[14105]='h00000e68;  wr_data_rom[14105]='h00000000;
    rd_cycle[14106] = 1'b1;  wr_cycle[14106] = 1'b0;  addr_rom[14106]='h0000234c;  wr_data_rom[14106]='h00000000;
    rd_cycle[14107] = 1'b1;  wr_cycle[14107] = 1'b0;  addr_rom[14107]='h000002b0;  wr_data_rom[14107]='h00000000;
    rd_cycle[14108] = 1'b1;  wr_cycle[14108] = 1'b0;  addr_rom[14108]='h00000ea4;  wr_data_rom[14108]='h00000000;
    rd_cycle[14109] = 1'b0;  wr_cycle[14109] = 1'b1;  addr_rom[14109]='h000025e0;  wr_data_rom[14109]='h000020c8;
    rd_cycle[14110] = 1'b1;  wr_cycle[14110] = 1'b0;  addr_rom[14110]='h00003d24;  wr_data_rom[14110]='h00000000;
    rd_cycle[14111] = 1'b1;  wr_cycle[14111] = 1'b0;  addr_rom[14111]='h0000234c;  wr_data_rom[14111]='h00000000;
    rd_cycle[14112] = 1'b1;  wr_cycle[14112] = 1'b0;  addr_rom[14112]='h0000212c;  wr_data_rom[14112]='h00000000;
    rd_cycle[14113] = 1'b0;  wr_cycle[14113] = 1'b1;  addr_rom[14113]='h00001798;  wr_data_rom[14113]='h0000253d;
    rd_cycle[14114] = 1'b1;  wr_cycle[14114] = 1'b0;  addr_rom[14114]='h00003b48;  wr_data_rom[14114]='h00000000;
    rd_cycle[14115] = 1'b1;  wr_cycle[14115] = 1'b0;  addr_rom[14115]='h00001cb0;  wr_data_rom[14115]='h00000000;
    rd_cycle[14116] = 1'b0;  wr_cycle[14116] = 1'b1;  addr_rom[14116]='h00001e14;  wr_data_rom[14116]='h00000436;
    rd_cycle[14117] = 1'b1;  wr_cycle[14117] = 1'b0;  addr_rom[14117]='h00000acc;  wr_data_rom[14117]='h00000000;
    rd_cycle[14118] = 1'b0;  wr_cycle[14118] = 1'b1;  addr_rom[14118]='h00000404;  wr_data_rom[14118]='h000029c6;
    rd_cycle[14119] = 1'b1;  wr_cycle[14119] = 1'b0;  addr_rom[14119]='h00001078;  wr_data_rom[14119]='h00000000;
    rd_cycle[14120] = 1'b0;  wr_cycle[14120] = 1'b1;  addr_rom[14120]='h000039b8;  wr_data_rom[14120]='h00003dd9;
    rd_cycle[14121] = 1'b0;  wr_cycle[14121] = 1'b1;  addr_rom[14121]='h00002154;  wr_data_rom[14121]='h000023b0;
    rd_cycle[14122] = 1'b1;  wr_cycle[14122] = 1'b0;  addr_rom[14122]='h00003adc;  wr_data_rom[14122]='h00000000;
    rd_cycle[14123] = 1'b1;  wr_cycle[14123] = 1'b0;  addr_rom[14123]='h000005dc;  wr_data_rom[14123]='h00000000;
    rd_cycle[14124] = 1'b0;  wr_cycle[14124] = 1'b1;  addr_rom[14124]='h000019f8;  wr_data_rom[14124]='h00003219;
    rd_cycle[14125] = 1'b1;  wr_cycle[14125] = 1'b0;  addr_rom[14125]='h00000528;  wr_data_rom[14125]='h00000000;
    rd_cycle[14126] = 1'b0;  wr_cycle[14126] = 1'b1;  addr_rom[14126]='h00001ad4;  wr_data_rom[14126]='h0000385b;
    rd_cycle[14127] = 1'b1;  wr_cycle[14127] = 1'b0;  addr_rom[14127]='h00002134;  wr_data_rom[14127]='h00000000;
    rd_cycle[14128] = 1'b1;  wr_cycle[14128] = 1'b0;  addr_rom[14128]='h00000af4;  wr_data_rom[14128]='h00000000;
    rd_cycle[14129] = 1'b1;  wr_cycle[14129] = 1'b0;  addr_rom[14129]='h00002c1c;  wr_data_rom[14129]='h00000000;
    rd_cycle[14130] = 1'b0;  wr_cycle[14130] = 1'b1;  addr_rom[14130]='h00001e50;  wr_data_rom[14130]='h00003d25;
    rd_cycle[14131] = 1'b0;  wr_cycle[14131] = 1'b1;  addr_rom[14131]='h00000dec;  wr_data_rom[14131]='h0000282d;
    rd_cycle[14132] = 1'b0;  wr_cycle[14132] = 1'b1;  addr_rom[14132]='h00000d64;  wr_data_rom[14132]='h00001a00;
    rd_cycle[14133] = 1'b1;  wr_cycle[14133] = 1'b0;  addr_rom[14133]='h00000d34;  wr_data_rom[14133]='h00000000;
    rd_cycle[14134] = 1'b1;  wr_cycle[14134] = 1'b0;  addr_rom[14134]='h00002cb4;  wr_data_rom[14134]='h00000000;
    rd_cycle[14135] = 1'b0;  wr_cycle[14135] = 1'b1;  addr_rom[14135]='h00001c40;  wr_data_rom[14135]='h000034bb;
    rd_cycle[14136] = 1'b0;  wr_cycle[14136] = 1'b1;  addr_rom[14136]='h00003e84;  wr_data_rom[14136]='h00001037;
    rd_cycle[14137] = 1'b0;  wr_cycle[14137] = 1'b1;  addr_rom[14137]='h00001bfc;  wr_data_rom[14137]='h000036a9;
    rd_cycle[14138] = 1'b1;  wr_cycle[14138] = 1'b0;  addr_rom[14138]='h0000299c;  wr_data_rom[14138]='h00000000;
    rd_cycle[14139] = 1'b0;  wr_cycle[14139] = 1'b1;  addr_rom[14139]='h00002978;  wr_data_rom[14139]='h00003fd2;
    rd_cycle[14140] = 1'b1;  wr_cycle[14140] = 1'b0;  addr_rom[14140]='h000036a0;  wr_data_rom[14140]='h00000000;
    rd_cycle[14141] = 1'b1;  wr_cycle[14141] = 1'b0;  addr_rom[14141]='h00002e94;  wr_data_rom[14141]='h00000000;
    rd_cycle[14142] = 1'b1;  wr_cycle[14142] = 1'b0;  addr_rom[14142]='h00001c40;  wr_data_rom[14142]='h00000000;
    rd_cycle[14143] = 1'b0;  wr_cycle[14143] = 1'b1;  addr_rom[14143]='h00001fa8;  wr_data_rom[14143]='h00003295;
    rd_cycle[14144] = 1'b0;  wr_cycle[14144] = 1'b1;  addr_rom[14144]='h00003750;  wr_data_rom[14144]='h000001a1;
    rd_cycle[14145] = 1'b1;  wr_cycle[14145] = 1'b0;  addr_rom[14145]='h000022d8;  wr_data_rom[14145]='h00000000;
    rd_cycle[14146] = 1'b1;  wr_cycle[14146] = 1'b0;  addr_rom[14146]='h000021d8;  wr_data_rom[14146]='h00000000;
    rd_cycle[14147] = 1'b1;  wr_cycle[14147] = 1'b0;  addr_rom[14147]='h00000f5c;  wr_data_rom[14147]='h00000000;
    rd_cycle[14148] = 1'b0;  wr_cycle[14148] = 1'b1;  addr_rom[14148]='h00000680;  wr_data_rom[14148]='h000003f4;
    rd_cycle[14149] = 1'b0;  wr_cycle[14149] = 1'b1;  addr_rom[14149]='h00002178;  wr_data_rom[14149]='h00002b31;
    rd_cycle[14150] = 1'b0;  wr_cycle[14150] = 1'b1;  addr_rom[14150]='h000030b4;  wr_data_rom[14150]='h00002bd7;
    rd_cycle[14151] = 1'b0;  wr_cycle[14151] = 1'b1;  addr_rom[14151]='h0000337c;  wr_data_rom[14151]='h00003ccd;
    rd_cycle[14152] = 1'b0;  wr_cycle[14152] = 1'b1;  addr_rom[14152]='h00003f60;  wr_data_rom[14152]='h00003cfb;
    rd_cycle[14153] = 1'b1;  wr_cycle[14153] = 1'b0;  addr_rom[14153]='h00001940;  wr_data_rom[14153]='h00000000;
    rd_cycle[14154] = 1'b0;  wr_cycle[14154] = 1'b1;  addr_rom[14154]='h000036e0;  wr_data_rom[14154]='h000018d5;
    rd_cycle[14155] = 1'b0;  wr_cycle[14155] = 1'b1;  addr_rom[14155]='h0000363c;  wr_data_rom[14155]='h00001a83;
    rd_cycle[14156] = 1'b1;  wr_cycle[14156] = 1'b0;  addr_rom[14156]='h00000ec0;  wr_data_rom[14156]='h00000000;
    rd_cycle[14157] = 1'b1;  wr_cycle[14157] = 1'b0;  addr_rom[14157]='h000003e8;  wr_data_rom[14157]='h00000000;
    rd_cycle[14158] = 1'b0;  wr_cycle[14158] = 1'b1;  addr_rom[14158]='h0000285c;  wr_data_rom[14158]='h00000c41;
    rd_cycle[14159] = 1'b0;  wr_cycle[14159] = 1'b1;  addr_rom[14159]='h00001ef8;  wr_data_rom[14159]='h00002e08;
    rd_cycle[14160] = 1'b1;  wr_cycle[14160] = 1'b0;  addr_rom[14160]='h00001d9c;  wr_data_rom[14160]='h00000000;
    rd_cycle[14161] = 1'b1;  wr_cycle[14161] = 1'b0;  addr_rom[14161]='h00000aa8;  wr_data_rom[14161]='h00000000;
    rd_cycle[14162] = 1'b0;  wr_cycle[14162] = 1'b1;  addr_rom[14162]='h00001a68;  wr_data_rom[14162]='h00001254;
    rd_cycle[14163] = 1'b1;  wr_cycle[14163] = 1'b0;  addr_rom[14163]='h0000150c;  wr_data_rom[14163]='h00000000;
    rd_cycle[14164] = 1'b1;  wr_cycle[14164] = 1'b0;  addr_rom[14164]='h00003130;  wr_data_rom[14164]='h00000000;
    rd_cycle[14165] = 1'b1;  wr_cycle[14165] = 1'b0;  addr_rom[14165]='h00001788;  wr_data_rom[14165]='h00000000;
    rd_cycle[14166] = 1'b1;  wr_cycle[14166] = 1'b0;  addr_rom[14166]='h0000275c;  wr_data_rom[14166]='h00000000;
    rd_cycle[14167] = 1'b1;  wr_cycle[14167] = 1'b0;  addr_rom[14167]='h000012d8;  wr_data_rom[14167]='h00000000;
    rd_cycle[14168] = 1'b0;  wr_cycle[14168] = 1'b1;  addr_rom[14168]='h00002098;  wr_data_rom[14168]='h000031e6;
    rd_cycle[14169] = 1'b1;  wr_cycle[14169] = 1'b0;  addr_rom[14169]='h00002a20;  wr_data_rom[14169]='h00000000;
    rd_cycle[14170] = 1'b0;  wr_cycle[14170] = 1'b1;  addr_rom[14170]='h00002610;  wr_data_rom[14170]='h0000261c;
    rd_cycle[14171] = 1'b1;  wr_cycle[14171] = 1'b0;  addr_rom[14171]='h00000404;  wr_data_rom[14171]='h00000000;
    rd_cycle[14172] = 1'b1;  wr_cycle[14172] = 1'b0;  addr_rom[14172]='h00003e10;  wr_data_rom[14172]='h00000000;
    rd_cycle[14173] = 1'b0;  wr_cycle[14173] = 1'b1;  addr_rom[14173]='h00002808;  wr_data_rom[14173]='h0000052b;
    rd_cycle[14174] = 1'b1;  wr_cycle[14174] = 1'b0;  addr_rom[14174]='h00003668;  wr_data_rom[14174]='h00000000;
    rd_cycle[14175] = 1'b1;  wr_cycle[14175] = 1'b0;  addr_rom[14175]='h00003bf0;  wr_data_rom[14175]='h00000000;
    rd_cycle[14176] = 1'b1;  wr_cycle[14176] = 1'b0;  addr_rom[14176]='h00000538;  wr_data_rom[14176]='h00000000;
    rd_cycle[14177] = 1'b1;  wr_cycle[14177] = 1'b0;  addr_rom[14177]='h00002ef4;  wr_data_rom[14177]='h00000000;
    rd_cycle[14178] = 1'b0;  wr_cycle[14178] = 1'b1;  addr_rom[14178]='h000024a4;  wr_data_rom[14178]='h00003d9e;
    rd_cycle[14179] = 1'b1;  wr_cycle[14179] = 1'b0;  addr_rom[14179]='h00001adc;  wr_data_rom[14179]='h00000000;
    rd_cycle[14180] = 1'b0;  wr_cycle[14180] = 1'b1;  addr_rom[14180]='h00002260;  wr_data_rom[14180]='h0000349e;
    rd_cycle[14181] = 1'b1;  wr_cycle[14181] = 1'b0;  addr_rom[14181]='h00000278;  wr_data_rom[14181]='h00000000;
    rd_cycle[14182] = 1'b1;  wr_cycle[14182] = 1'b0;  addr_rom[14182]='h00001944;  wr_data_rom[14182]='h00000000;
    rd_cycle[14183] = 1'b1;  wr_cycle[14183] = 1'b0;  addr_rom[14183]='h00002400;  wr_data_rom[14183]='h00000000;
    rd_cycle[14184] = 1'b0;  wr_cycle[14184] = 1'b1;  addr_rom[14184]='h00001e9c;  wr_data_rom[14184]='h00003c6f;
    rd_cycle[14185] = 1'b1;  wr_cycle[14185] = 1'b0;  addr_rom[14185]='h000021c8;  wr_data_rom[14185]='h00000000;
    rd_cycle[14186] = 1'b1;  wr_cycle[14186] = 1'b0;  addr_rom[14186]='h00002100;  wr_data_rom[14186]='h00000000;
    rd_cycle[14187] = 1'b0;  wr_cycle[14187] = 1'b1;  addr_rom[14187]='h00000ddc;  wr_data_rom[14187]='h00003900;
    rd_cycle[14188] = 1'b0;  wr_cycle[14188] = 1'b1;  addr_rom[14188]='h000031e4;  wr_data_rom[14188]='h00001d3d;
    rd_cycle[14189] = 1'b1;  wr_cycle[14189] = 1'b0;  addr_rom[14189]='h00002c94;  wr_data_rom[14189]='h00000000;
    rd_cycle[14190] = 1'b0;  wr_cycle[14190] = 1'b1;  addr_rom[14190]='h00000350;  wr_data_rom[14190]='h000023c6;
    rd_cycle[14191] = 1'b0;  wr_cycle[14191] = 1'b1;  addr_rom[14191]='h00000ef8;  wr_data_rom[14191]='h00000aea;
    rd_cycle[14192] = 1'b1;  wr_cycle[14192] = 1'b0;  addr_rom[14192]='h00001104;  wr_data_rom[14192]='h00000000;
    rd_cycle[14193] = 1'b1;  wr_cycle[14193] = 1'b0;  addr_rom[14193]='h00001500;  wr_data_rom[14193]='h00000000;
    rd_cycle[14194] = 1'b0;  wr_cycle[14194] = 1'b1;  addr_rom[14194]='h00002f80;  wr_data_rom[14194]='h00001e2c;
    rd_cycle[14195] = 1'b0;  wr_cycle[14195] = 1'b1;  addr_rom[14195]='h00003f70;  wr_data_rom[14195]='h000025d4;
    rd_cycle[14196] = 1'b1;  wr_cycle[14196] = 1'b0;  addr_rom[14196]='h00003074;  wr_data_rom[14196]='h00000000;
    rd_cycle[14197] = 1'b1;  wr_cycle[14197] = 1'b0;  addr_rom[14197]='h0000362c;  wr_data_rom[14197]='h00000000;
    rd_cycle[14198] = 1'b1;  wr_cycle[14198] = 1'b0;  addr_rom[14198]='h000003b8;  wr_data_rom[14198]='h00000000;
    rd_cycle[14199] = 1'b1;  wr_cycle[14199] = 1'b0;  addr_rom[14199]='h00000484;  wr_data_rom[14199]='h00000000;
    rd_cycle[14200] = 1'b1;  wr_cycle[14200] = 1'b0;  addr_rom[14200]='h0000328c;  wr_data_rom[14200]='h00000000;
    rd_cycle[14201] = 1'b0;  wr_cycle[14201] = 1'b1;  addr_rom[14201]='h0000081c;  wr_data_rom[14201]='h00000d6c;
    rd_cycle[14202] = 1'b0;  wr_cycle[14202] = 1'b1;  addr_rom[14202]='h0000249c;  wr_data_rom[14202]='h00002b71;
    rd_cycle[14203] = 1'b1;  wr_cycle[14203] = 1'b0;  addr_rom[14203]='h000026e8;  wr_data_rom[14203]='h00000000;
    rd_cycle[14204] = 1'b1;  wr_cycle[14204] = 1'b0;  addr_rom[14204]='h00002710;  wr_data_rom[14204]='h00000000;
    rd_cycle[14205] = 1'b1;  wr_cycle[14205] = 1'b0;  addr_rom[14205]='h00000cf4;  wr_data_rom[14205]='h00000000;
    rd_cycle[14206] = 1'b0;  wr_cycle[14206] = 1'b1;  addr_rom[14206]='h000019ec;  wr_data_rom[14206]='h0000295e;
    rd_cycle[14207] = 1'b0;  wr_cycle[14207] = 1'b1;  addr_rom[14207]='h00003064;  wr_data_rom[14207]='h000037d4;
    rd_cycle[14208] = 1'b0;  wr_cycle[14208] = 1'b1;  addr_rom[14208]='h00001108;  wr_data_rom[14208]='h00003d3c;
    rd_cycle[14209] = 1'b0;  wr_cycle[14209] = 1'b1;  addr_rom[14209]='h000022e0;  wr_data_rom[14209]='h000021f2;
    rd_cycle[14210] = 1'b0;  wr_cycle[14210] = 1'b1;  addr_rom[14210]='h00003668;  wr_data_rom[14210]='h00003be0;
    rd_cycle[14211] = 1'b0;  wr_cycle[14211] = 1'b1;  addr_rom[14211]='h00002568;  wr_data_rom[14211]='h00001e68;
    rd_cycle[14212] = 1'b0;  wr_cycle[14212] = 1'b1;  addr_rom[14212]='h00000870;  wr_data_rom[14212]='h00002964;
    rd_cycle[14213] = 1'b1;  wr_cycle[14213] = 1'b0;  addr_rom[14213]='h000009f4;  wr_data_rom[14213]='h00000000;
    rd_cycle[14214] = 1'b1;  wr_cycle[14214] = 1'b0;  addr_rom[14214]='h00002314;  wr_data_rom[14214]='h00000000;
    rd_cycle[14215] = 1'b1;  wr_cycle[14215] = 1'b0;  addr_rom[14215]='h00001c08;  wr_data_rom[14215]='h00000000;
    rd_cycle[14216] = 1'b1;  wr_cycle[14216] = 1'b0;  addr_rom[14216]='h00001788;  wr_data_rom[14216]='h00000000;
    rd_cycle[14217] = 1'b0;  wr_cycle[14217] = 1'b1;  addr_rom[14217]='h00001288;  wr_data_rom[14217]='h0000108b;
    rd_cycle[14218] = 1'b0;  wr_cycle[14218] = 1'b1;  addr_rom[14218]='h00002ec8;  wr_data_rom[14218]='h000012ac;
    rd_cycle[14219] = 1'b1;  wr_cycle[14219] = 1'b0;  addr_rom[14219]='h00000680;  wr_data_rom[14219]='h00000000;
    rd_cycle[14220] = 1'b1;  wr_cycle[14220] = 1'b0;  addr_rom[14220]='h000009a8;  wr_data_rom[14220]='h00000000;
    rd_cycle[14221] = 1'b1;  wr_cycle[14221] = 1'b0;  addr_rom[14221]='h0000120c;  wr_data_rom[14221]='h00000000;
    rd_cycle[14222] = 1'b0;  wr_cycle[14222] = 1'b1;  addr_rom[14222]='h00000aa0;  wr_data_rom[14222]='h00003382;
    rd_cycle[14223] = 1'b0;  wr_cycle[14223] = 1'b1;  addr_rom[14223]='h000031e8;  wr_data_rom[14223]='h00000f6e;
    rd_cycle[14224] = 1'b0;  wr_cycle[14224] = 1'b1;  addr_rom[14224]='h00000d54;  wr_data_rom[14224]='h000000ab;
    rd_cycle[14225] = 1'b0;  wr_cycle[14225] = 1'b1;  addr_rom[14225]='h00001044;  wr_data_rom[14225]='h00001854;
    rd_cycle[14226] = 1'b1;  wr_cycle[14226] = 1'b0;  addr_rom[14226]='h00002eb8;  wr_data_rom[14226]='h00000000;
    rd_cycle[14227] = 1'b0;  wr_cycle[14227] = 1'b1;  addr_rom[14227]='h00003264;  wr_data_rom[14227]='h00001aa2;
    rd_cycle[14228] = 1'b0;  wr_cycle[14228] = 1'b1;  addr_rom[14228]='h000002c4;  wr_data_rom[14228]='h00001df4;
    rd_cycle[14229] = 1'b0;  wr_cycle[14229] = 1'b1;  addr_rom[14229]='h00001040;  wr_data_rom[14229]='h000014d4;
    rd_cycle[14230] = 1'b0;  wr_cycle[14230] = 1'b1;  addr_rom[14230]='h00003ef4;  wr_data_rom[14230]='h00002e6e;
    rd_cycle[14231] = 1'b0;  wr_cycle[14231] = 1'b1;  addr_rom[14231]='h00002950;  wr_data_rom[14231]='h000009b8;
    rd_cycle[14232] = 1'b0;  wr_cycle[14232] = 1'b1;  addr_rom[14232]='h000001f8;  wr_data_rom[14232]='h000029da;
    rd_cycle[14233] = 1'b1;  wr_cycle[14233] = 1'b0;  addr_rom[14233]='h00000d5c;  wr_data_rom[14233]='h00000000;
    rd_cycle[14234] = 1'b0;  wr_cycle[14234] = 1'b1;  addr_rom[14234]='h00003e98;  wr_data_rom[14234]='h00001d39;
    rd_cycle[14235] = 1'b1;  wr_cycle[14235] = 1'b0;  addr_rom[14235]='h00002cf4;  wr_data_rom[14235]='h00000000;
    rd_cycle[14236] = 1'b1;  wr_cycle[14236] = 1'b0;  addr_rom[14236]='h00001f94;  wr_data_rom[14236]='h00000000;
    rd_cycle[14237] = 1'b1;  wr_cycle[14237] = 1'b0;  addr_rom[14237]='h00002960;  wr_data_rom[14237]='h00000000;
    rd_cycle[14238] = 1'b0;  wr_cycle[14238] = 1'b1;  addr_rom[14238]='h00000830;  wr_data_rom[14238]='h00001842;
    rd_cycle[14239] = 1'b0;  wr_cycle[14239] = 1'b1;  addr_rom[14239]='h00003890;  wr_data_rom[14239]='h000008da;
    rd_cycle[14240] = 1'b0;  wr_cycle[14240] = 1'b1;  addr_rom[14240]='h00002694;  wr_data_rom[14240]='h0000330f;
    rd_cycle[14241] = 1'b0;  wr_cycle[14241] = 1'b1;  addr_rom[14241]='h00000200;  wr_data_rom[14241]='h000032b2;
    rd_cycle[14242] = 1'b0;  wr_cycle[14242] = 1'b1;  addr_rom[14242]='h00003c48;  wr_data_rom[14242]='h00002d9b;
    rd_cycle[14243] = 1'b0;  wr_cycle[14243] = 1'b1;  addr_rom[14243]='h000015dc;  wr_data_rom[14243]='h00001351;
    rd_cycle[14244] = 1'b1;  wr_cycle[14244] = 1'b0;  addr_rom[14244]='h00003eec;  wr_data_rom[14244]='h00000000;
    rd_cycle[14245] = 1'b1;  wr_cycle[14245] = 1'b0;  addr_rom[14245]='h00002540;  wr_data_rom[14245]='h00000000;
    rd_cycle[14246] = 1'b0;  wr_cycle[14246] = 1'b1;  addr_rom[14246]='h00000be4;  wr_data_rom[14246]='h00002c16;
    rd_cycle[14247] = 1'b0;  wr_cycle[14247] = 1'b1;  addr_rom[14247]='h00000af4;  wr_data_rom[14247]='h00002765;
    rd_cycle[14248] = 1'b0;  wr_cycle[14248] = 1'b1;  addr_rom[14248]='h00002888;  wr_data_rom[14248]='h000025af;
    rd_cycle[14249] = 1'b1;  wr_cycle[14249] = 1'b0;  addr_rom[14249]='h00001cf4;  wr_data_rom[14249]='h00000000;
    rd_cycle[14250] = 1'b1;  wr_cycle[14250] = 1'b0;  addr_rom[14250]='h000012d4;  wr_data_rom[14250]='h00000000;
    rd_cycle[14251] = 1'b0;  wr_cycle[14251] = 1'b1;  addr_rom[14251]='h000026d8;  wr_data_rom[14251]='h0000114d;
    rd_cycle[14252] = 1'b0;  wr_cycle[14252] = 1'b1;  addr_rom[14252]='h00000428;  wr_data_rom[14252]='h00000a48;
    rd_cycle[14253] = 1'b1;  wr_cycle[14253] = 1'b0;  addr_rom[14253]='h00000f78;  wr_data_rom[14253]='h00000000;
    rd_cycle[14254] = 1'b1;  wr_cycle[14254] = 1'b0;  addr_rom[14254]='h00000a58;  wr_data_rom[14254]='h00000000;
    rd_cycle[14255] = 1'b1;  wr_cycle[14255] = 1'b0;  addr_rom[14255]='h00000348;  wr_data_rom[14255]='h00000000;
    rd_cycle[14256] = 1'b1;  wr_cycle[14256] = 1'b0;  addr_rom[14256]='h00000158;  wr_data_rom[14256]='h00000000;
    rd_cycle[14257] = 1'b1;  wr_cycle[14257] = 1'b0;  addr_rom[14257]='h00000dcc;  wr_data_rom[14257]='h00000000;
    rd_cycle[14258] = 1'b0;  wr_cycle[14258] = 1'b1;  addr_rom[14258]='h00001934;  wr_data_rom[14258]='h000007f7;
    rd_cycle[14259] = 1'b1;  wr_cycle[14259] = 1'b0;  addr_rom[14259]='h00001480;  wr_data_rom[14259]='h00000000;
    rd_cycle[14260] = 1'b1;  wr_cycle[14260] = 1'b0;  addr_rom[14260]='h00003418;  wr_data_rom[14260]='h00000000;
    rd_cycle[14261] = 1'b0;  wr_cycle[14261] = 1'b1;  addr_rom[14261]='h00000fa4;  wr_data_rom[14261]='h0000323a;
    rd_cycle[14262] = 1'b0;  wr_cycle[14262] = 1'b1;  addr_rom[14262]='h00002878;  wr_data_rom[14262]='h0000337f;
    rd_cycle[14263] = 1'b1;  wr_cycle[14263] = 1'b0;  addr_rom[14263]='h00001664;  wr_data_rom[14263]='h00000000;
    rd_cycle[14264] = 1'b0;  wr_cycle[14264] = 1'b1;  addr_rom[14264]='h00002a44;  wr_data_rom[14264]='h00001832;
    rd_cycle[14265] = 1'b0;  wr_cycle[14265] = 1'b1;  addr_rom[14265]='h00001de8;  wr_data_rom[14265]='h00000881;
    rd_cycle[14266] = 1'b1;  wr_cycle[14266] = 1'b0;  addr_rom[14266]='h00003b78;  wr_data_rom[14266]='h00000000;
    rd_cycle[14267] = 1'b1;  wr_cycle[14267] = 1'b0;  addr_rom[14267]='h00003f9c;  wr_data_rom[14267]='h00000000;
    rd_cycle[14268] = 1'b1;  wr_cycle[14268] = 1'b0;  addr_rom[14268]='h000010b4;  wr_data_rom[14268]='h00000000;
    rd_cycle[14269] = 1'b1;  wr_cycle[14269] = 1'b0;  addr_rom[14269]='h00003488;  wr_data_rom[14269]='h00000000;
    rd_cycle[14270] = 1'b0;  wr_cycle[14270] = 1'b1;  addr_rom[14270]='h00002df0;  wr_data_rom[14270]='h00001902;
    rd_cycle[14271] = 1'b0;  wr_cycle[14271] = 1'b1;  addr_rom[14271]='h00002fbc;  wr_data_rom[14271]='h0000171d;
    rd_cycle[14272] = 1'b0;  wr_cycle[14272] = 1'b1;  addr_rom[14272]='h000024fc;  wr_data_rom[14272]='h000038c6;
    rd_cycle[14273] = 1'b1;  wr_cycle[14273] = 1'b0;  addr_rom[14273]='h00002d44;  wr_data_rom[14273]='h00000000;
    rd_cycle[14274] = 1'b0;  wr_cycle[14274] = 1'b1;  addr_rom[14274]='h00003c64;  wr_data_rom[14274]='h000001ef;
    rd_cycle[14275] = 1'b0;  wr_cycle[14275] = 1'b1;  addr_rom[14275]='h000023d8;  wr_data_rom[14275]='h000021eb;
    rd_cycle[14276] = 1'b1;  wr_cycle[14276] = 1'b0;  addr_rom[14276]='h00001b20;  wr_data_rom[14276]='h00000000;
    rd_cycle[14277] = 1'b0;  wr_cycle[14277] = 1'b1;  addr_rom[14277]='h00000d38;  wr_data_rom[14277]='h00002846;
    rd_cycle[14278] = 1'b1;  wr_cycle[14278] = 1'b0;  addr_rom[14278]='h00000cf4;  wr_data_rom[14278]='h00000000;
    rd_cycle[14279] = 1'b0;  wr_cycle[14279] = 1'b1;  addr_rom[14279]='h00000558;  wr_data_rom[14279]='h00002c7f;
    rd_cycle[14280] = 1'b1;  wr_cycle[14280] = 1'b0;  addr_rom[14280]='h000002e0;  wr_data_rom[14280]='h00000000;
    rd_cycle[14281] = 1'b1;  wr_cycle[14281] = 1'b0;  addr_rom[14281]='h00002e1c;  wr_data_rom[14281]='h00000000;
    rd_cycle[14282] = 1'b0;  wr_cycle[14282] = 1'b1;  addr_rom[14282]='h00002c10;  wr_data_rom[14282]='h0000312f;
    rd_cycle[14283] = 1'b1;  wr_cycle[14283] = 1'b0;  addr_rom[14283]='h00001188;  wr_data_rom[14283]='h00000000;
    rd_cycle[14284] = 1'b1;  wr_cycle[14284] = 1'b0;  addr_rom[14284]='h000015dc;  wr_data_rom[14284]='h00000000;
    rd_cycle[14285] = 1'b0;  wr_cycle[14285] = 1'b1;  addr_rom[14285]='h00001368;  wr_data_rom[14285]='h0000014c;
    rd_cycle[14286] = 1'b1;  wr_cycle[14286] = 1'b0;  addr_rom[14286]='h000026c4;  wr_data_rom[14286]='h00000000;
    rd_cycle[14287] = 1'b1;  wr_cycle[14287] = 1'b0;  addr_rom[14287]='h00001a78;  wr_data_rom[14287]='h00000000;
    rd_cycle[14288] = 1'b0;  wr_cycle[14288] = 1'b1;  addr_rom[14288]='h000017d0;  wr_data_rom[14288]='h00001f48;
    rd_cycle[14289] = 1'b1;  wr_cycle[14289] = 1'b0;  addr_rom[14289]='h00000e7c;  wr_data_rom[14289]='h00000000;
    rd_cycle[14290] = 1'b1;  wr_cycle[14290] = 1'b0;  addr_rom[14290]='h0000110c;  wr_data_rom[14290]='h00000000;
    rd_cycle[14291] = 1'b0;  wr_cycle[14291] = 1'b1;  addr_rom[14291]='h000028d0;  wr_data_rom[14291]='h000036b9;
    rd_cycle[14292] = 1'b0;  wr_cycle[14292] = 1'b1;  addr_rom[14292]='h000027dc;  wr_data_rom[14292]='h00001bf2;
    rd_cycle[14293] = 1'b1;  wr_cycle[14293] = 1'b0;  addr_rom[14293]='h00002154;  wr_data_rom[14293]='h00000000;
    rd_cycle[14294] = 1'b1;  wr_cycle[14294] = 1'b0;  addr_rom[14294]='h00002084;  wr_data_rom[14294]='h00000000;
    rd_cycle[14295] = 1'b1;  wr_cycle[14295] = 1'b0;  addr_rom[14295]='h000028f0;  wr_data_rom[14295]='h00000000;
    rd_cycle[14296] = 1'b0;  wr_cycle[14296] = 1'b1;  addr_rom[14296]='h00003158;  wr_data_rom[14296]='h00003476;
    rd_cycle[14297] = 1'b1;  wr_cycle[14297] = 1'b0;  addr_rom[14297]='h00000b54;  wr_data_rom[14297]='h00000000;
    rd_cycle[14298] = 1'b1;  wr_cycle[14298] = 1'b0;  addr_rom[14298]='h000004ac;  wr_data_rom[14298]='h00000000;
    rd_cycle[14299] = 1'b0;  wr_cycle[14299] = 1'b1;  addr_rom[14299]='h00000ec8;  wr_data_rom[14299]='h00003706;
    rd_cycle[14300] = 1'b0;  wr_cycle[14300] = 1'b1;  addr_rom[14300]='h00003ed8;  wr_data_rom[14300]='h00000f1e;
    rd_cycle[14301] = 1'b0;  wr_cycle[14301] = 1'b1;  addr_rom[14301]='h000038c0;  wr_data_rom[14301]='h0000003a;
    rd_cycle[14302] = 1'b1;  wr_cycle[14302] = 1'b0;  addr_rom[14302]='h00000a6c;  wr_data_rom[14302]='h00000000;
    rd_cycle[14303] = 1'b1;  wr_cycle[14303] = 1'b0;  addr_rom[14303]='h000017f4;  wr_data_rom[14303]='h00000000;
    rd_cycle[14304] = 1'b0;  wr_cycle[14304] = 1'b1;  addr_rom[14304]='h00000aec;  wr_data_rom[14304]='h0000181c;
    rd_cycle[14305] = 1'b0;  wr_cycle[14305] = 1'b1;  addr_rom[14305]='h0000370c;  wr_data_rom[14305]='h000005d7;
    rd_cycle[14306] = 1'b1;  wr_cycle[14306] = 1'b0;  addr_rom[14306]='h00000700;  wr_data_rom[14306]='h00000000;
    rd_cycle[14307] = 1'b1;  wr_cycle[14307] = 1'b0;  addr_rom[14307]='h000036c8;  wr_data_rom[14307]='h00000000;
    rd_cycle[14308] = 1'b0;  wr_cycle[14308] = 1'b1;  addr_rom[14308]='h00002ed8;  wr_data_rom[14308]='h00000782;
    rd_cycle[14309] = 1'b1;  wr_cycle[14309] = 1'b0;  addr_rom[14309]='h00001218;  wr_data_rom[14309]='h00000000;
    rd_cycle[14310] = 1'b1;  wr_cycle[14310] = 1'b0;  addr_rom[14310]='h00000ea4;  wr_data_rom[14310]='h00000000;
    rd_cycle[14311] = 1'b0;  wr_cycle[14311] = 1'b1;  addr_rom[14311]='h00002ae0;  wr_data_rom[14311]='h0000236f;
    rd_cycle[14312] = 1'b1;  wr_cycle[14312] = 1'b0;  addr_rom[14312]='h00001a34;  wr_data_rom[14312]='h00000000;
    rd_cycle[14313] = 1'b1;  wr_cycle[14313] = 1'b0;  addr_rom[14313]='h000010e0;  wr_data_rom[14313]='h00000000;
    rd_cycle[14314] = 1'b1;  wr_cycle[14314] = 1'b0;  addr_rom[14314]='h000029d4;  wr_data_rom[14314]='h00000000;
    rd_cycle[14315] = 1'b0;  wr_cycle[14315] = 1'b1;  addr_rom[14315]='h000039e4;  wr_data_rom[14315]='h00000054;
    rd_cycle[14316] = 1'b0;  wr_cycle[14316] = 1'b1;  addr_rom[14316]='h00000474;  wr_data_rom[14316]='h00000ed4;
    rd_cycle[14317] = 1'b1;  wr_cycle[14317] = 1'b0;  addr_rom[14317]='h00003cec;  wr_data_rom[14317]='h00000000;
    rd_cycle[14318] = 1'b0;  wr_cycle[14318] = 1'b1;  addr_rom[14318]='h00001c84;  wr_data_rom[14318]='h000003be;
    rd_cycle[14319] = 1'b1;  wr_cycle[14319] = 1'b0;  addr_rom[14319]='h000009a8;  wr_data_rom[14319]='h00000000;
    rd_cycle[14320] = 1'b0;  wr_cycle[14320] = 1'b1;  addr_rom[14320]='h00000fb8;  wr_data_rom[14320]='h00002b1a;
    rd_cycle[14321] = 1'b0;  wr_cycle[14321] = 1'b1;  addr_rom[14321]='h00003334;  wr_data_rom[14321]='h00001f9b;
    rd_cycle[14322] = 1'b1;  wr_cycle[14322] = 1'b0;  addr_rom[14322]='h00001120;  wr_data_rom[14322]='h00000000;
    rd_cycle[14323] = 1'b0;  wr_cycle[14323] = 1'b1;  addr_rom[14323]='h00001abc;  wr_data_rom[14323]='h000020d0;
    rd_cycle[14324] = 1'b0;  wr_cycle[14324] = 1'b1;  addr_rom[14324]='h00003538;  wr_data_rom[14324]='h00003be2;
    rd_cycle[14325] = 1'b1;  wr_cycle[14325] = 1'b0;  addr_rom[14325]='h000035f4;  wr_data_rom[14325]='h00000000;
    rd_cycle[14326] = 1'b1;  wr_cycle[14326] = 1'b0;  addr_rom[14326]='h000012d0;  wr_data_rom[14326]='h00000000;
    rd_cycle[14327] = 1'b0;  wr_cycle[14327] = 1'b1;  addr_rom[14327]='h00000e84;  wr_data_rom[14327]='h00000834;
    rd_cycle[14328] = 1'b1;  wr_cycle[14328] = 1'b0;  addr_rom[14328]='h000005bc;  wr_data_rom[14328]='h00000000;
    rd_cycle[14329] = 1'b1;  wr_cycle[14329] = 1'b0;  addr_rom[14329]='h000003b0;  wr_data_rom[14329]='h00000000;
    rd_cycle[14330] = 1'b0;  wr_cycle[14330] = 1'b1;  addr_rom[14330]='h0000186c;  wr_data_rom[14330]='h00000ca0;
    rd_cycle[14331] = 1'b0;  wr_cycle[14331] = 1'b1;  addr_rom[14331]='h00001f2c;  wr_data_rom[14331]='h0000372a;
    rd_cycle[14332] = 1'b0;  wr_cycle[14332] = 1'b1;  addr_rom[14332]='h00000238;  wr_data_rom[14332]='h00003363;
    rd_cycle[14333] = 1'b0;  wr_cycle[14333] = 1'b1;  addr_rom[14333]='h00003b78;  wr_data_rom[14333]='h000012ff;
    rd_cycle[14334] = 1'b1;  wr_cycle[14334] = 1'b0;  addr_rom[14334]='h000026b0;  wr_data_rom[14334]='h00000000;
    rd_cycle[14335] = 1'b0;  wr_cycle[14335] = 1'b1;  addr_rom[14335]='h00003be4;  wr_data_rom[14335]='h00002ffc;
    rd_cycle[14336] = 1'b0;  wr_cycle[14336] = 1'b1;  addr_rom[14336]='h00002644;  wr_data_rom[14336]='h00000484;
    rd_cycle[14337] = 1'b0;  wr_cycle[14337] = 1'b1;  addr_rom[14337]='h000029bc;  wr_data_rom[14337]='h0000317d;
    rd_cycle[14338] = 1'b1;  wr_cycle[14338] = 1'b0;  addr_rom[14338]='h000021d4;  wr_data_rom[14338]='h00000000;
    rd_cycle[14339] = 1'b0;  wr_cycle[14339] = 1'b1;  addr_rom[14339]='h00003598;  wr_data_rom[14339]='h00000103;
    rd_cycle[14340] = 1'b0;  wr_cycle[14340] = 1'b1;  addr_rom[14340]='h000014b0;  wr_data_rom[14340]='h00001ca3;
    rd_cycle[14341] = 1'b1;  wr_cycle[14341] = 1'b0;  addr_rom[14341]='h00000814;  wr_data_rom[14341]='h00000000;
    rd_cycle[14342] = 1'b1;  wr_cycle[14342] = 1'b0;  addr_rom[14342]='h000016f4;  wr_data_rom[14342]='h00000000;
    rd_cycle[14343] = 1'b0;  wr_cycle[14343] = 1'b1;  addr_rom[14343]='h000008f4;  wr_data_rom[14343]='h00000b50;
    rd_cycle[14344] = 1'b0;  wr_cycle[14344] = 1'b1;  addr_rom[14344]='h00001470;  wr_data_rom[14344]='h00000b04;
    rd_cycle[14345] = 1'b0;  wr_cycle[14345] = 1'b1;  addr_rom[14345]='h00000b8c;  wr_data_rom[14345]='h000037e4;
    rd_cycle[14346] = 1'b0;  wr_cycle[14346] = 1'b1;  addr_rom[14346]='h00000b54;  wr_data_rom[14346]='h000003db;
    rd_cycle[14347] = 1'b0;  wr_cycle[14347] = 1'b1;  addr_rom[14347]='h00001930;  wr_data_rom[14347]='h000004b6;
    rd_cycle[14348] = 1'b0;  wr_cycle[14348] = 1'b1;  addr_rom[14348]='h00002784;  wr_data_rom[14348]='h00003f83;
    rd_cycle[14349] = 1'b0;  wr_cycle[14349] = 1'b1;  addr_rom[14349]='h00002d64;  wr_data_rom[14349]='h000013ac;
    rd_cycle[14350] = 1'b0;  wr_cycle[14350] = 1'b1;  addr_rom[14350]='h000008f8;  wr_data_rom[14350]='h0000119f;
    rd_cycle[14351] = 1'b0;  wr_cycle[14351] = 1'b1;  addr_rom[14351]='h0000260c;  wr_data_rom[14351]='h00003fb7;
    rd_cycle[14352] = 1'b0;  wr_cycle[14352] = 1'b1;  addr_rom[14352]='h00001c58;  wr_data_rom[14352]='h00001638;
    rd_cycle[14353] = 1'b1;  wr_cycle[14353] = 1'b0;  addr_rom[14353]='h0000297c;  wr_data_rom[14353]='h00000000;
    rd_cycle[14354] = 1'b1;  wr_cycle[14354] = 1'b0;  addr_rom[14354]='h000004e4;  wr_data_rom[14354]='h00000000;
    rd_cycle[14355] = 1'b0;  wr_cycle[14355] = 1'b1;  addr_rom[14355]='h00002dd8;  wr_data_rom[14355]='h00001a11;
    rd_cycle[14356] = 1'b0;  wr_cycle[14356] = 1'b1;  addr_rom[14356]='h00002f00;  wr_data_rom[14356]='h00001a25;
    rd_cycle[14357] = 1'b1;  wr_cycle[14357] = 1'b0;  addr_rom[14357]='h000005a4;  wr_data_rom[14357]='h00000000;
    rd_cycle[14358] = 1'b0;  wr_cycle[14358] = 1'b1;  addr_rom[14358]='h00003190;  wr_data_rom[14358]='h000012c8;
    rd_cycle[14359] = 1'b0;  wr_cycle[14359] = 1'b1;  addr_rom[14359]='h000022d0;  wr_data_rom[14359]='h0000065c;
    rd_cycle[14360] = 1'b0;  wr_cycle[14360] = 1'b1;  addr_rom[14360]='h00002504;  wr_data_rom[14360]='h0000104d;
    rd_cycle[14361] = 1'b0;  wr_cycle[14361] = 1'b1;  addr_rom[14361]='h00000cf8;  wr_data_rom[14361]='h00002c52;
    rd_cycle[14362] = 1'b1;  wr_cycle[14362] = 1'b0;  addr_rom[14362]='h000014f8;  wr_data_rom[14362]='h00000000;
    rd_cycle[14363] = 1'b0;  wr_cycle[14363] = 1'b1;  addr_rom[14363]='h00001258;  wr_data_rom[14363]='h00002ec1;
    rd_cycle[14364] = 1'b1;  wr_cycle[14364] = 1'b0;  addr_rom[14364]='h00001d78;  wr_data_rom[14364]='h00000000;
    rd_cycle[14365] = 1'b0;  wr_cycle[14365] = 1'b1;  addr_rom[14365]='h00000708;  wr_data_rom[14365]='h000018ea;
    rd_cycle[14366] = 1'b0;  wr_cycle[14366] = 1'b1;  addr_rom[14366]='h00000b4c;  wr_data_rom[14366]='h00000a0d;
    rd_cycle[14367] = 1'b1;  wr_cycle[14367] = 1'b0;  addr_rom[14367]='h00001280;  wr_data_rom[14367]='h00000000;
    rd_cycle[14368] = 1'b1;  wr_cycle[14368] = 1'b0;  addr_rom[14368]='h00001dcc;  wr_data_rom[14368]='h00000000;
    rd_cycle[14369] = 1'b1;  wr_cycle[14369] = 1'b0;  addr_rom[14369]='h000011e4;  wr_data_rom[14369]='h00000000;
    rd_cycle[14370] = 1'b1;  wr_cycle[14370] = 1'b0;  addr_rom[14370]='h0000302c;  wr_data_rom[14370]='h00000000;
    rd_cycle[14371] = 1'b0;  wr_cycle[14371] = 1'b1;  addr_rom[14371]='h00002110;  wr_data_rom[14371]='h000023ca;
    rd_cycle[14372] = 1'b0;  wr_cycle[14372] = 1'b1;  addr_rom[14372]='h00000464;  wr_data_rom[14372]='h0000275d;
    rd_cycle[14373] = 1'b0;  wr_cycle[14373] = 1'b1;  addr_rom[14373]='h0000054c;  wr_data_rom[14373]='h000021cc;
    rd_cycle[14374] = 1'b0;  wr_cycle[14374] = 1'b1;  addr_rom[14374]='h00000cdc;  wr_data_rom[14374]='h00000f10;
    rd_cycle[14375] = 1'b0;  wr_cycle[14375] = 1'b1;  addr_rom[14375]='h00002a54;  wr_data_rom[14375]='h000018eb;
    rd_cycle[14376] = 1'b1;  wr_cycle[14376] = 1'b0;  addr_rom[14376]='h00002934;  wr_data_rom[14376]='h00000000;
    rd_cycle[14377] = 1'b0;  wr_cycle[14377] = 1'b1;  addr_rom[14377]='h000005dc;  wr_data_rom[14377]='h00002c4b;
    rd_cycle[14378] = 1'b1;  wr_cycle[14378] = 1'b0;  addr_rom[14378]='h00002078;  wr_data_rom[14378]='h00000000;
    rd_cycle[14379] = 1'b1;  wr_cycle[14379] = 1'b0;  addr_rom[14379]='h00000ff4;  wr_data_rom[14379]='h00000000;
    rd_cycle[14380] = 1'b0;  wr_cycle[14380] = 1'b1;  addr_rom[14380]='h00000d84;  wr_data_rom[14380]='h00003992;
    rd_cycle[14381] = 1'b1;  wr_cycle[14381] = 1'b0;  addr_rom[14381]='h00003c24;  wr_data_rom[14381]='h00000000;
    rd_cycle[14382] = 1'b0;  wr_cycle[14382] = 1'b1;  addr_rom[14382]='h00000210;  wr_data_rom[14382]='h00000fa7;
    rd_cycle[14383] = 1'b1;  wr_cycle[14383] = 1'b0;  addr_rom[14383]='h00000a9c;  wr_data_rom[14383]='h00000000;
    rd_cycle[14384] = 1'b0;  wr_cycle[14384] = 1'b1;  addr_rom[14384]='h000039f4;  wr_data_rom[14384]='h000003da;
    rd_cycle[14385] = 1'b0;  wr_cycle[14385] = 1'b1;  addr_rom[14385]='h00001144;  wr_data_rom[14385]='h00003ab9;
    rd_cycle[14386] = 1'b1;  wr_cycle[14386] = 1'b0;  addr_rom[14386]='h000002ac;  wr_data_rom[14386]='h00000000;
    rd_cycle[14387] = 1'b1;  wr_cycle[14387] = 1'b0;  addr_rom[14387]='h00001bd0;  wr_data_rom[14387]='h00000000;
    rd_cycle[14388] = 1'b0;  wr_cycle[14388] = 1'b1;  addr_rom[14388]='h00000a04;  wr_data_rom[14388]='h00001f23;
    rd_cycle[14389] = 1'b1;  wr_cycle[14389] = 1'b0;  addr_rom[14389]='h0000368c;  wr_data_rom[14389]='h00000000;
    rd_cycle[14390] = 1'b1;  wr_cycle[14390] = 1'b0;  addr_rom[14390]='h00002450;  wr_data_rom[14390]='h00000000;
    rd_cycle[14391] = 1'b0;  wr_cycle[14391] = 1'b1;  addr_rom[14391]='h00003a7c;  wr_data_rom[14391]='h000015dc;
    rd_cycle[14392] = 1'b1;  wr_cycle[14392] = 1'b0;  addr_rom[14392]='h000022a8;  wr_data_rom[14392]='h00000000;
    rd_cycle[14393] = 1'b0;  wr_cycle[14393] = 1'b1;  addr_rom[14393]='h00002738;  wr_data_rom[14393]='h00002b1a;
    rd_cycle[14394] = 1'b0;  wr_cycle[14394] = 1'b1;  addr_rom[14394]='h00003b58;  wr_data_rom[14394]='h00001f5c;
    rd_cycle[14395] = 1'b1;  wr_cycle[14395] = 1'b0;  addr_rom[14395]='h00003374;  wr_data_rom[14395]='h00000000;
    rd_cycle[14396] = 1'b1;  wr_cycle[14396] = 1'b0;  addr_rom[14396]='h00001ea0;  wr_data_rom[14396]='h00000000;
    rd_cycle[14397] = 1'b0;  wr_cycle[14397] = 1'b1;  addr_rom[14397]='h000024e8;  wr_data_rom[14397]='h0000066d;
    rd_cycle[14398] = 1'b0;  wr_cycle[14398] = 1'b1;  addr_rom[14398]='h00001d1c;  wr_data_rom[14398]='h00000942;
    rd_cycle[14399] = 1'b1;  wr_cycle[14399] = 1'b0;  addr_rom[14399]='h000023c4;  wr_data_rom[14399]='h00000000;
    rd_cycle[14400] = 1'b0;  wr_cycle[14400] = 1'b1;  addr_rom[14400]='h000026f8;  wr_data_rom[14400]='h00000615;
    rd_cycle[14401] = 1'b1;  wr_cycle[14401] = 1'b0;  addr_rom[14401]='h000039b4;  wr_data_rom[14401]='h00000000;
    rd_cycle[14402] = 1'b0;  wr_cycle[14402] = 1'b1;  addr_rom[14402]='h00000788;  wr_data_rom[14402]='h00002e30;
    rd_cycle[14403] = 1'b1;  wr_cycle[14403] = 1'b0;  addr_rom[14403]='h000039cc;  wr_data_rom[14403]='h00000000;
    rd_cycle[14404] = 1'b0;  wr_cycle[14404] = 1'b1;  addr_rom[14404]='h00003e9c;  wr_data_rom[14404]='h00001d12;
    rd_cycle[14405] = 1'b1;  wr_cycle[14405] = 1'b0;  addr_rom[14405]='h00003998;  wr_data_rom[14405]='h00000000;
    rd_cycle[14406] = 1'b1;  wr_cycle[14406] = 1'b0;  addr_rom[14406]='h00000dbc;  wr_data_rom[14406]='h00000000;
    rd_cycle[14407] = 1'b1;  wr_cycle[14407] = 1'b0;  addr_rom[14407]='h000024d4;  wr_data_rom[14407]='h00000000;
    rd_cycle[14408] = 1'b1;  wr_cycle[14408] = 1'b0;  addr_rom[14408]='h00000748;  wr_data_rom[14408]='h00000000;
    rd_cycle[14409] = 1'b0;  wr_cycle[14409] = 1'b1;  addr_rom[14409]='h0000341c;  wr_data_rom[14409]='h00002e55;
    rd_cycle[14410] = 1'b1;  wr_cycle[14410] = 1'b0;  addr_rom[14410]='h00002b58;  wr_data_rom[14410]='h00000000;
    rd_cycle[14411] = 1'b1;  wr_cycle[14411] = 1'b0;  addr_rom[14411]='h00000ec4;  wr_data_rom[14411]='h00000000;
    rd_cycle[14412] = 1'b1;  wr_cycle[14412] = 1'b0;  addr_rom[14412]='h000001f0;  wr_data_rom[14412]='h00000000;
    rd_cycle[14413] = 1'b0;  wr_cycle[14413] = 1'b1;  addr_rom[14413]='h0000330c;  wr_data_rom[14413]='h0000165d;
    rd_cycle[14414] = 1'b0;  wr_cycle[14414] = 1'b1;  addr_rom[14414]='h00000214;  wr_data_rom[14414]='h00003c63;
    rd_cycle[14415] = 1'b1;  wr_cycle[14415] = 1'b0;  addr_rom[14415]='h00003154;  wr_data_rom[14415]='h00000000;
    rd_cycle[14416] = 1'b1;  wr_cycle[14416] = 1'b0;  addr_rom[14416]='h00000ab4;  wr_data_rom[14416]='h00000000;
    rd_cycle[14417] = 1'b1;  wr_cycle[14417] = 1'b0;  addr_rom[14417]='h00002310;  wr_data_rom[14417]='h00000000;
    rd_cycle[14418] = 1'b1;  wr_cycle[14418] = 1'b0;  addr_rom[14418]='h00001058;  wr_data_rom[14418]='h00000000;
    rd_cycle[14419] = 1'b0;  wr_cycle[14419] = 1'b1;  addr_rom[14419]='h00003428;  wr_data_rom[14419]='h0000253f;
    rd_cycle[14420] = 1'b0;  wr_cycle[14420] = 1'b1;  addr_rom[14420]='h00000800;  wr_data_rom[14420]='h0000335f;
    rd_cycle[14421] = 1'b1;  wr_cycle[14421] = 1'b0;  addr_rom[14421]='h000004cc;  wr_data_rom[14421]='h00000000;
    rd_cycle[14422] = 1'b0;  wr_cycle[14422] = 1'b1;  addr_rom[14422]='h0000168c;  wr_data_rom[14422]='h000015b4;
    rd_cycle[14423] = 1'b0;  wr_cycle[14423] = 1'b1;  addr_rom[14423]='h000002cc;  wr_data_rom[14423]='h000010cd;
    rd_cycle[14424] = 1'b1;  wr_cycle[14424] = 1'b0;  addr_rom[14424]='h00001b6c;  wr_data_rom[14424]='h00000000;
    rd_cycle[14425] = 1'b0;  wr_cycle[14425] = 1'b1;  addr_rom[14425]='h00003c5c;  wr_data_rom[14425]='h00000ec7;
    rd_cycle[14426] = 1'b0;  wr_cycle[14426] = 1'b1;  addr_rom[14426]='h00000e60;  wr_data_rom[14426]='h00001b4b;
    rd_cycle[14427] = 1'b0;  wr_cycle[14427] = 1'b1;  addr_rom[14427]='h0000392c;  wr_data_rom[14427]='h00003c09;
    rd_cycle[14428] = 1'b0;  wr_cycle[14428] = 1'b1;  addr_rom[14428]='h000006f0;  wr_data_rom[14428]='h00002d73;
    rd_cycle[14429] = 1'b1;  wr_cycle[14429] = 1'b0;  addr_rom[14429]='h00000fdc;  wr_data_rom[14429]='h00000000;
    rd_cycle[14430] = 1'b1;  wr_cycle[14430] = 1'b0;  addr_rom[14430]='h00001d70;  wr_data_rom[14430]='h00000000;
    rd_cycle[14431] = 1'b1;  wr_cycle[14431] = 1'b0;  addr_rom[14431]='h00003fb0;  wr_data_rom[14431]='h00000000;
    rd_cycle[14432] = 1'b1;  wr_cycle[14432] = 1'b0;  addr_rom[14432]='h00000df4;  wr_data_rom[14432]='h00000000;
    rd_cycle[14433] = 1'b1;  wr_cycle[14433] = 1'b0;  addr_rom[14433]='h00001bf4;  wr_data_rom[14433]='h00000000;
    rd_cycle[14434] = 1'b1;  wr_cycle[14434] = 1'b0;  addr_rom[14434]='h00003afc;  wr_data_rom[14434]='h00000000;
    rd_cycle[14435] = 1'b0;  wr_cycle[14435] = 1'b1;  addr_rom[14435]='h00001904;  wr_data_rom[14435]='h00001967;
    rd_cycle[14436] = 1'b0;  wr_cycle[14436] = 1'b1;  addr_rom[14436]='h000021c0;  wr_data_rom[14436]='h0000231d;
    rd_cycle[14437] = 1'b0;  wr_cycle[14437] = 1'b1;  addr_rom[14437]='h000011b0;  wr_data_rom[14437]='h00001137;
    rd_cycle[14438] = 1'b0;  wr_cycle[14438] = 1'b1;  addr_rom[14438]='h00002e4c;  wr_data_rom[14438]='h000035c8;
    rd_cycle[14439] = 1'b0;  wr_cycle[14439] = 1'b1;  addr_rom[14439]='h00001008;  wr_data_rom[14439]='h00001fd4;
    rd_cycle[14440] = 1'b1;  wr_cycle[14440] = 1'b0;  addr_rom[14440]='h00002c64;  wr_data_rom[14440]='h00000000;
    rd_cycle[14441] = 1'b0;  wr_cycle[14441] = 1'b1;  addr_rom[14441]='h00003218;  wr_data_rom[14441]='h00000f23;
    rd_cycle[14442] = 1'b0;  wr_cycle[14442] = 1'b1;  addr_rom[14442]='h000022b0;  wr_data_rom[14442]='h000037f7;
    rd_cycle[14443] = 1'b0;  wr_cycle[14443] = 1'b1;  addr_rom[14443]='h000020f4;  wr_data_rom[14443]='h0000130f;
    rd_cycle[14444] = 1'b1;  wr_cycle[14444] = 1'b0;  addr_rom[14444]='h000020e8;  wr_data_rom[14444]='h00000000;
    rd_cycle[14445] = 1'b1;  wr_cycle[14445] = 1'b0;  addr_rom[14445]='h000018d0;  wr_data_rom[14445]='h00000000;
    rd_cycle[14446] = 1'b0;  wr_cycle[14446] = 1'b1;  addr_rom[14446]='h00001b0c;  wr_data_rom[14446]='h00000009;
    rd_cycle[14447] = 1'b1;  wr_cycle[14447] = 1'b0;  addr_rom[14447]='h000020a4;  wr_data_rom[14447]='h00000000;
    rd_cycle[14448] = 1'b1;  wr_cycle[14448] = 1'b0;  addr_rom[14448]='h00001c90;  wr_data_rom[14448]='h00000000;
    rd_cycle[14449] = 1'b1;  wr_cycle[14449] = 1'b0;  addr_rom[14449]='h00001dd8;  wr_data_rom[14449]='h00000000;
    rd_cycle[14450] = 1'b0;  wr_cycle[14450] = 1'b1;  addr_rom[14450]='h00002610;  wr_data_rom[14450]='h00003d3b;
    rd_cycle[14451] = 1'b1;  wr_cycle[14451] = 1'b0;  addr_rom[14451]='h00000768;  wr_data_rom[14451]='h00000000;
    rd_cycle[14452] = 1'b1;  wr_cycle[14452] = 1'b0;  addr_rom[14452]='h00001690;  wr_data_rom[14452]='h00000000;
    rd_cycle[14453] = 1'b1;  wr_cycle[14453] = 1'b0;  addr_rom[14453]='h000032a4;  wr_data_rom[14453]='h00000000;
    rd_cycle[14454] = 1'b0;  wr_cycle[14454] = 1'b1;  addr_rom[14454]='h00000570;  wr_data_rom[14454]='h000015a0;
    rd_cycle[14455] = 1'b1;  wr_cycle[14455] = 1'b0;  addr_rom[14455]='h000034a4;  wr_data_rom[14455]='h00000000;
    rd_cycle[14456] = 1'b0;  wr_cycle[14456] = 1'b1;  addr_rom[14456]='h0000111c;  wr_data_rom[14456]='h0000184b;
    rd_cycle[14457] = 1'b1;  wr_cycle[14457] = 1'b0;  addr_rom[14457]='h00003e98;  wr_data_rom[14457]='h00000000;
    rd_cycle[14458] = 1'b1;  wr_cycle[14458] = 1'b0;  addr_rom[14458]='h00003cd4;  wr_data_rom[14458]='h00000000;
    rd_cycle[14459] = 1'b1;  wr_cycle[14459] = 1'b0;  addr_rom[14459]='h0000275c;  wr_data_rom[14459]='h00000000;
    rd_cycle[14460] = 1'b1;  wr_cycle[14460] = 1'b0;  addr_rom[14460]='h000036e0;  wr_data_rom[14460]='h00000000;
    rd_cycle[14461] = 1'b0;  wr_cycle[14461] = 1'b1;  addr_rom[14461]='h000024ac;  wr_data_rom[14461]='h00000a9d;
    rd_cycle[14462] = 1'b1;  wr_cycle[14462] = 1'b0;  addr_rom[14462]='h00002b8c;  wr_data_rom[14462]='h00000000;
    rd_cycle[14463] = 1'b0;  wr_cycle[14463] = 1'b1;  addr_rom[14463]='h00002a70;  wr_data_rom[14463]='h000039bb;
    rd_cycle[14464] = 1'b1;  wr_cycle[14464] = 1'b0;  addr_rom[14464]='h00003664;  wr_data_rom[14464]='h00000000;
    rd_cycle[14465] = 1'b1;  wr_cycle[14465] = 1'b0;  addr_rom[14465]='h00003464;  wr_data_rom[14465]='h00000000;
    rd_cycle[14466] = 1'b1;  wr_cycle[14466] = 1'b0;  addr_rom[14466]='h00003220;  wr_data_rom[14466]='h00000000;
    rd_cycle[14467] = 1'b1;  wr_cycle[14467] = 1'b0;  addr_rom[14467]='h0000235c;  wr_data_rom[14467]='h00000000;
    rd_cycle[14468] = 1'b1;  wr_cycle[14468] = 1'b0;  addr_rom[14468]='h00000168;  wr_data_rom[14468]='h00000000;
    rd_cycle[14469] = 1'b1;  wr_cycle[14469] = 1'b0;  addr_rom[14469]='h00001d18;  wr_data_rom[14469]='h00000000;
    rd_cycle[14470] = 1'b1;  wr_cycle[14470] = 1'b0;  addr_rom[14470]='h00002c88;  wr_data_rom[14470]='h00000000;
    rd_cycle[14471] = 1'b1;  wr_cycle[14471] = 1'b0;  addr_rom[14471]='h00002c1c;  wr_data_rom[14471]='h00000000;
    rd_cycle[14472] = 1'b1;  wr_cycle[14472] = 1'b0;  addr_rom[14472]='h0000102c;  wr_data_rom[14472]='h00000000;
    rd_cycle[14473] = 1'b0;  wr_cycle[14473] = 1'b1;  addr_rom[14473]='h000028ac;  wr_data_rom[14473]='h00003ca3;
    rd_cycle[14474] = 1'b1;  wr_cycle[14474] = 1'b0;  addr_rom[14474]='h0000075c;  wr_data_rom[14474]='h00000000;
    rd_cycle[14475] = 1'b0;  wr_cycle[14475] = 1'b1;  addr_rom[14475]='h00001724;  wr_data_rom[14475]='h0000230b;
    rd_cycle[14476] = 1'b0;  wr_cycle[14476] = 1'b1;  addr_rom[14476]='h00003038;  wr_data_rom[14476]='h00003cb5;
    rd_cycle[14477] = 1'b1;  wr_cycle[14477] = 1'b0;  addr_rom[14477]='h00001238;  wr_data_rom[14477]='h00000000;
    rd_cycle[14478] = 1'b1;  wr_cycle[14478] = 1'b0;  addr_rom[14478]='h0000185c;  wr_data_rom[14478]='h00000000;
    rd_cycle[14479] = 1'b0;  wr_cycle[14479] = 1'b1;  addr_rom[14479]='h00000478;  wr_data_rom[14479]='h00000eb7;
    rd_cycle[14480] = 1'b1;  wr_cycle[14480] = 1'b0;  addr_rom[14480]='h000032bc;  wr_data_rom[14480]='h00000000;
    rd_cycle[14481] = 1'b0;  wr_cycle[14481] = 1'b1;  addr_rom[14481]='h000004d0;  wr_data_rom[14481]='h00003f92;
    rd_cycle[14482] = 1'b1;  wr_cycle[14482] = 1'b0;  addr_rom[14482]='h00002fb8;  wr_data_rom[14482]='h00000000;
    rd_cycle[14483] = 1'b1;  wr_cycle[14483] = 1'b0;  addr_rom[14483]='h00000b6c;  wr_data_rom[14483]='h00000000;
    rd_cycle[14484] = 1'b1;  wr_cycle[14484] = 1'b0;  addr_rom[14484]='h00000254;  wr_data_rom[14484]='h00000000;
    rd_cycle[14485] = 1'b0;  wr_cycle[14485] = 1'b1;  addr_rom[14485]='h00001650;  wr_data_rom[14485]='h00002da7;
    rd_cycle[14486] = 1'b1;  wr_cycle[14486] = 1'b0;  addr_rom[14486]='h00000788;  wr_data_rom[14486]='h00000000;
    rd_cycle[14487] = 1'b0;  wr_cycle[14487] = 1'b1;  addr_rom[14487]='h00003dfc;  wr_data_rom[14487]='h00001497;
    rd_cycle[14488] = 1'b1;  wr_cycle[14488] = 1'b0;  addr_rom[14488]='h00002760;  wr_data_rom[14488]='h00000000;
    rd_cycle[14489] = 1'b1;  wr_cycle[14489] = 1'b0;  addr_rom[14489]='h00001e34;  wr_data_rom[14489]='h00000000;
    rd_cycle[14490] = 1'b1;  wr_cycle[14490] = 1'b0;  addr_rom[14490]='h00003a40;  wr_data_rom[14490]='h00000000;
    rd_cycle[14491] = 1'b1;  wr_cycle[14491] = 1'b0;  addr_rom[14491]='h0000309c;  wr_data_rom[14491]='h00000000;
    rd_cycle[14492] = 1'b0;  wr_cycle[14492] = 1'b1;  addr_rom[14492]='h00003a00;  wr_data_rom[14492]='h00002f27;
    rd_cycle[14493] = 1'b0;  wr_cycle[14493] = 1'b1;  addr_rom[14493]='h00000fcc;  wr_data_rom[14493]='h000005e6;
    rd_cycle[14494] = 1'b0;  wr_cycle[14494] = 1'b1;  addr_rom[14494]='h00003bc0;  wr_data_rom[14494]='h000022c6;
    rd_cycle[14495] = 1'b1;  wr_cycle[14495] = 1'b0;  addr_rom[14495]='h000033dc;  wr_data_rom[14495]='h00000000;
    rd_cycle[14496] = 1'b0;  wr_cycle[14496] = 1'b1;  addr_rom[14496]='h000035b4;  wr_data_rom[14496]='h0000104f;
    rd_cycle[14497] = 1'b0;  wr_cycle[14497] = 1'b1;  addr_rom[14497]='h00003bac;  wr_data_rom[14497]='h00003536;
    rd_cycle[14498] = 1'b1;  wr_cycle[14498] = 1'b0;  addr_rom[14498]='h00001fc0;  wr_data_rom[14498]='h00000000;
    rd_cycle[14499] = 1'b1;  wr_cycle[14499] = 1'b0;  addr_rom[14499]='h00001ea8;  wr_data_rom[14499]='h00000000;
    rd_cycle[14500] = 1'b1;  wr_cycle[14500] = 1'b0;  addr_rom[14500]='h00001760;  wr_data_rom[14500]='h00000000;
    rd_cycle[14501] = 1'b1;  wr_cycle[14501] = 1'b0;  addr_rom[14501]='h0000268c;  wr_data_rom[14501]='h00000000;
    rd_cycle[14502] = 1'b1;  wr_cycle[14502] = 1'b0;  addr_rom[14502]='h00000f0c;  wr_data_rom[14502]='h00000000;
    rd_cycle[14503] = 1'b1;  wr_cycle[14503] = 1'b0;  addr_rom[14503]='h000023a0;  wr_data_rom[14503]='h00000000;
    rd_cycle[14504] = 1'b0;  wr_cycle[14504] = 1'b1;  addr_rom[14504]='h000015ec;  wr_data_rom[14504]='h00000607;
    rd_cycle[14505] = 1'b0;  wr_cycle[14505] = 1'b1;  addr_rom[14505]='h0000083c;  wr_data_rom[14505]='h000008a1;
    rd_cycle[14506] = 1'b1;  wr_cycle[14506] = 1'b0;  addr_rom[14506]='h00002e68;  wr_data_rom[14506]='h00000000;
    rd_cycle[14507] = 1'b1;  wr_cycle[14507] = 1'b0;  addr_rom[14507]='h00002cf8;  wr_data_rom[14507]='h00000000;
    rd_cycle[14508] = 1'b1;  wr_cycle[14508] = 1'b0;  addr_rom[14508]='h00000900;  wr_data_rom[14508]='h00000000;
    rd_cycle[14509] = 1'b1;  wr_cycle[14509] = 1'b0;  addr_rom[14509]='h00001018;  wr_data_rom[14509]='h00000000;
    rd_cycle[14510] = 1'b0;  wr_cycle[14510] = 1'b1;  addr_rom[14510]='h00001a44;  wr_data_rom[14510]='h00003d9d;
    rd_cycle[14511] = 1'b1;  wr_cycle[14511] = 1'b0;  addr_rom[14511]='h00002598;  wr_data_rom[14511]='h00000000;
    rd_cycle[14512] = 1'b1;  wr_cycle[14512] = 1'b0;  addr_rom[14512]='h00003838;  wr_data_rom[14512]='h00000000;
    rd_cycle[14513] = 1'b0;  wr_cycle[14513] = 1'b1;  addr_rom[14513]='h000034e4;  wr_data_rom[14513]='h000007e3;
    rd_cycle[14514] = 1'b1;  wr_cycle[14514] = 1'b0;  addr_rom[14514]='h00002698;  wr_data_rom[14514]='h00000000;
    rd_cycle[14515] = 1'b1;  wr_cycle[14515] = 1'b0;  addr_rom[14515]='h000002a0;  wr_data_rom[14515]='h00000000;
    rd_cycle[14516] = 1'b1;  wr_cycle[14516] = 1'b0;  addr_rom[14516]='h0000097c;  wr_data_rom[14516]='h00000000;
    rd_cycle[14517] = 1'b1;  wr_cycle[14517] = 1'b0;  addr_rom[14517]='h000002ac;  wr_data_rom[14517]='h00000000;
    rd_cycle[14518] = 1'b1;  wr_cycle[14518] = 1'b0;  addr_rom[14518]='h00002ee8;  wr_data_rom[14518]='h00000000;
    rd_cycle[14519] = 1'b0;  wr_cycle[14519] = 1'b1;  addr_rom[14519]='h000039d8;  wr_data_rom[14519]='h00001ec0;
    rd_cycle[14520] = 1'b0;  wr_cycle[14520] = 1'b1;  addr_rom[14520]='h00003b9c;  wr_data_rom[14520]='h00003489;
    rd_cycle[14521] = 1'b0;  wr_cycle[14521] = 1'b1;  addr_rom[14521]='h00003274;  wr_data_rom[14521]='h00001dbd;
    rd_cycle[14522] = 1'b0;  wr_cycle[14522] = 1'b1;  addr_rom[14522]='h00001760;  wr_data_rom[14522]='h000031b3;
    rd_cycle[14523] = 1'b1;  wr_cycle[14523] = 1'b0;  addr_rom[14523]='h00001f84;  wr_data_rom[14523]='h00000000;
    rd_cycle[14524] = 1'b0;  wr_cycle[14524] = 1'b1;  addr_rom[14524]='h00002f68;  wr_data_rom[14524]='h00002645;
    rd_cycle[14525] = 1'b0;  wr_cycle[14525] = 1'b1;  addr_rom[14525]='h00002b04;  wr_data_rom[14525]='h0000305b;
    rd_cycle[14526] = 1'b1;  wr_cycle[14526] = 1'b0;  addr_rom[14526]='h0000105c;  wr_data_rom[14526]='h00000000;
    rd_cycle[14527] = 1'b1;  wr_cycle[14527] = 1'b0;  addr_rom[14527]='h000026d0;  wr_data_rom[14527]='h00000000;
    rd_cycle[14528] = 1'b0;  wr_cycle[14528] = 1'b1;  addr_rom[14528]='h00000070;  wr_data_rom[14528]='h00000bf0;
    rd_cycle[14529] = 1'b1;  wr_cycle[14529] = 1'b0;  addr_rom[14529]='h00002b04;  wr_data_rom[14529]='h00000000;
    rd_cycle[14530] = 1'b1;  wr_cycle[14530] = 1'b0;  addr_rom[14530]='h00001e34;  wr_data_rom[14530]='h00000000;
    rd_cycle[14531] = 1'b1;  wr_cycle[14531] = 1'b0;  addr_rom[14531]='h00001828;  wr_data_rom[14531]='h00000000;
    rd_cycle[14532] = 1'b0;  wr_cycle[14532] = 1'b1;  addr_rom[14532]='h00001368;  wr_data_rom[14532]='h0000277b;
    rd_cycle[14533] = 1'b1;  wr_cycle[14533] = 1'b0;  addr_rom[14533]='h00001ac0;  wr_data_rom[14533]='h00000000;
    rd_cycle[14534] = 1'b0;  wr_cycle[14534] = 1'b1;  addr_rom[14534]='h00001b7c;  wr_data_rom[14534]='h00000d8e;
    rd_cycle[14535] = 1'b0;  wr_cycle[14535] = 1'b1;  addr_rom[14535]='h00003cb8;  wr_data_rom[14535]='h00003908;
    rd_cycle[14536] = 1'b0;  wr_cycle[14536] = 1'b1;  addr_rom[14536]='h00003994;  wr_data_rom[14536]='h000013e9;
    rd_cycle[14537] = 1'b0;  wr_cycle[14537] = 1'b1;  addr_rom[14537]='h00000940;  wr_data_rom[14537]='h0000072c;
    rd_cycle[14538] = 1'b0;  wr_cycle[14538] = 1'b1;  addr_rom[14538]='h000032d4;  wr_data_rom[14538]='h0000209d;
    rd_cycle[14539] = 1'b0;  wr_cycle[14539] = 1'b1;  addr_rom[14539]='h00000770;  wr_data_rom[14539]='h00003493;
    rd_cycle[14540] = 1'b1;  wr_cycle[14540] = 1'b0;  addr_rom[14540]='h000012dc;  wr_data_rom[14540]='h00000000;
    rd_cycle[14541] = 1'b1;  wr_cycle[14541] = 1'b0;  addr_rom[14541]='h000021b8;  wr_data_rom[14541]='h00000000;
    rd_cycle[14542] = 1'b0;  wr_cycle[14542] = 1'b1;  addr_rom[14542]='h00000e38;  wr_data_rom[14542]='h0000111a;
    rd_cycle[14543] = 1'b0;  wr_cycle[14543] = 1'b1;  addr_rom[14543]='h000005e4;  wr_data_rom[14543]='h00001efa;
    rd_cycle[14544] = 1'b1;  wr_cycle[14544] = 1'b0;  addr_rom[14544]='h00002eb4;  wr_data_rom[14544]='h00000000;
    rd_cycle[14545] = 1'b1;  wr_cycle[14545] = 1'b0;  addr_rom[14545]='h00000a64;  wr_data_rom[14545]='h00000000;
    rd_cycle[14546] = 1'b1;  wr_cycle[14546] = 1'b0;  addr_rom[14546]='h00001c2c;  wr_data_rom[14546]='h00000000;
    rd_cycle[14547] = 1'b0;  wr_cycle[14547] = 1'b1;  addr_rom[14547]='h00002430;  wr_data_rom[14547]='h00000675;
    rd_cycle[14548] = 1'b1;  wr_cycle[14548] = 1'b0;  addr_rom[14548]='h0000379c;  wr_data_rom[14548]='h00000000;
    rd_cycle[14549] = 1'b0;  wr_cycle[14549] = 1'b1;  addr_rom[14549]='h000019d4;  wr_data_rom[14549]='h00001aa0;
    rd_cycle[14550] = 1'b0;  wr_cycle[14550] = 1'b1;  addr_rom[14550]='h00002d84;  wr_data_rom[14550]='h00000a06;
    rd_cycle[14551] = 1'b1;  wr_cycle[14551] = 1'b0;  addr_rom[14551]='h00003428;  wr_data_rom[14551]='h00000000;
    rd_cycle[14552] = 1'b0;  wr_cycle[14552] = 1'b1;  addr_rom[14552]='h00003228;  wr_data_rom[14552]='h00000431;
    rd_cycle[14553] = 1'b1;  wr_cycle[14553] = 1'b0;  addr_rom[14553]='h0000252c;  wr_data_rom[14553]='h00000000;
    rd_cycle[14554] = 1'b0;  wr_cycle[14554] = 1'b1;  addr_rom[14554]='h00000c60;  wr_data_rom[14554]='h00002de2;
    rd_cycle[14555] = 1'b1;  wr_cycle[14555] = 1'b0;  addr_rom[14555]='h00000abc;  wr_data_rom[14555]='h00000000;
    rd_cycle[14556] = 1'b1;  wr_cycle[14556] = 1'b0;  addr_rom[14556]='h000005a4;  wr_data_rom[14556]='h00000000;
    rd_cycle[14557] = 1'b0;  wr_cycle[14557] = 1'b1;  addr_rom[14557]='h00001ddc;  wr_data_rom[14557]='h00000acd;
    rd_cycle[14558] = 1'b1;  wr_cycle[14558] = 1'b0;  addr_rom[14558]='h00000534;  wr_data_rom[14558]='h00000000;
    rd_cycle[14559] = 1'b0;  wr_cycle[14559] = 1'b1;  addr_rom[14559]='h00000244;  wr_data_rom[14559]='h00002bc2;
    rd_cycle[14560] = 1'b1;  wr_cycle[14560] = 1'b0;  addr_rom[14560]='h00002bd0;  wr_data_rom[14560]='h00000000;
    rd_cycle[14561] = 1'b0;  wr_cycle[14561] = 1'b1;  addr_rom[14561]='h00000cac;  wr_data_rom[14561]='h000032e5;
    rd_cycle[14562] = 1'b1;  wr_cycle[14562] = 1'b0;  addr_rom[14562]='h00002248;  wr_data_rom[14562]='h00000000;
    rd_cycle[14563] = 1'b0;  wr_cycle[14563] = 1'b1;  addr_rom[14563]='h00001088;  wr_data_rom[14563]='h00002949;
    rd_cycle[14564] = 1'b0;  wr_cycle[14564] = 1'b1;  addr_rom[14564]='h00001a48;  wr_data_rom[14564]='h000027d3;
    rd_cycle[14565] = 1'b0;  wr_cycle[14565] = 1'b1;  addr_rom[14565]='h00000e60;  wr_data_rom[14565]='h000039f4;
    rd_cycle[14566] = 1'b0;  wr_cycle[14566] = 1'b1;  addr_rom[14566]='h00000f74;  wr_data_rom[14566]='h000024e1;
    rd_cycle[14567] = 1'b0;  wr_cycle[14567] = 1'b1;  addr_rom[14567]='h00003c2c;  wr_data_rom[14567]='h000004a3;
    rd_cycle[14568] = 1'b0;  wr_cycle[14568] = 1'b1;  addr_rom[14568]='h00003bd8;  wr_data_rom[14568]='h000031f2;
    rd_cycle[14569] = 1'b0;  wr_cycle[14569] = 1'b1;  addr_rom[14569]='h000003cc;  wr_data_rom[14569]='h00001500;
    rd_cycle[14570] = 1'b0;  wr_cycle[14570] = 1'b1;  addr_rom[14570]='h000033dc;  wr_data_rom[14570]='h00003550;
    rd_cycle[14571] = 1'b1;  wr_cycle[14571] = 1'b0;  addr_rom[14571]='h000004e0;  wr_data_rom[14571]='h00000000;
    rd_cycle[14572] = 1'b1;  wr_cycle[14572] = 1'b0;  addr_rom[14572]='h00001ba0;  wr_data_rom[14572]='h00000000;
    rd_cycle[14573] = 1'b1;  wr_cycle[14573] = 1'b0;  addr_rom[14573]='h000018b8;  wr_data_rom[14573]='h00000000;
    rd_cycle[14574] = 1'b1;  wr_cycle[14574] = 1'b0;  addr_rom[14574]='h00003a08;  wr_data_rom[14574]='h00000000;
    rd_cycle[14575] = 1'b0;  wr_cycle[14575] = 1'b1;  addr_rom[14575]='h000018fc;  wr_data_rom[14575]='h00001c67;
    rd_cycle[14576] = 1'b0;  wr_cycle[14576] = 1'b1;  addr_rom[14576]='h00002abc;  wr_data_rom[14576]='h00003bb6;
    rd_cycle[14577] = 1'b0;  wr_cycle[14577] = 1'b1;  addr_rom[14577]='h000000d4;  wr_data_rom[14577]='h00001d2e;
    rd_cycle[14578] = 1'b1;  wr_cycle[14578] = 1'b0;  addr_rom[14578]='h00003768;  wr_data_rom[14578]='h00000000;
    rd_cycle[14579] = 1'b1;  wr_cycle[14579] = 1'b0;  addr_rom[14579]='h00003410;  wr_data_rom[14579]='h00000000;
    rd_cycle[14580] = 1'b1;  wr_cycle[14580] = 1'b0;  addr_rom[14580]='h00003e98;  wr_data_rom[14580]='h00000000;
    rd_cycle[14581] = 1'b0;  wr_cycle[14581] = 1'b1;  addr_rom[14581]='h000025ac;  wr_data_rom[14581]='h00001604;
    rd_cycle[14582] = 1'b0;  wr_cycle[14582] = 1'b1;  addr_rom[14582]='h000014a8;  wr_data_rom[14582]='h00001212;
    rd_cycle[14583] = 1'b1;  wr_cycle[14583] = 1'b0;  addr_rom[14583]='h000037c8;  wr_data_rom[14583]='h00000000;
    rd_cycle[14584] = 1'b0;  wr_cycle[14584] = 1'b1;  addr_rom[14584]='h000001f0;  wr_data_rom[14584]='h00001692;
    rd_cycle[14585] = 1'b0;  wr_cycle[14585] = 1'b1;  addr_rom[14585]='h00002288;  wr_data_rom[14585]='h00003897;
    rd_cycle[14586] = 1'b0;  wr_cycle[14586] = 1'b1;  addr_rom[14586]='h000007e4;  wr_data_rom[14586]='h00003d74;
    rd_cycle[14587] = 1'b0;  wr_cycle[14587] = 1'b1;  addr_rom[14587]='h00001624;  wr_data_rom[14587]='h00002144;
    rd_cycle[14588] = 1'b0;  wr_cycle[14588] = 1'b1;  addr_rom[14588]='h0000388c;  wr_data_rom[14588]='h0000011d;
    rd_cycle[14589] = 1'b1;  wr_cycle[14589] = 1'b0;  addr_rom[14589]='h00000228;  wr_data_rom[14589]='h00000000;
    rd_cycle[14590] = 1'b1;  wr_cycle[14590] = 1'b0;  addr_rom[14590]='h0000151c;  wr_data_rom[14590]='h00000000;
    rd_cycle[14591] = 1'b0;  wr_cycle[14591] = 1'b1;  addr_rom[14591]='h00003200;  wr_data_rom[14591]='h0000296c;
    rd_cycle[14592] = 1'b0;  wr_cycle[14592] = 1'b1;  addr_rom[14592]='h00002980;  wr_data_rom[14592]='h00003bf0;
    rd_cycle[14593] = 1'b1;  wr_cycle[14593] = 1'b0;  addr_rom[14593]='h000014c4;  wr_data_rom[14593]='h00000000;
    rd_cycle[14594] = 1'b1;  wr_cycle[14594] = 1'b0;  addr_rom[14594]='h000016ac;  wr_data_rom[14594]='h00000000;
    rd_cycle[14595] = 1'b1;  wr_cycle[14595] = 1'b0;  addr_rom[14595]='h0000159c;  wr_data_rom[14595]='h00000000;
    rd_cycle[14596] = 1'b0;  wr_cycle[14596] = 1'b1;  addr_rom[14596]='h00000b50;  wr_data_rom[14596]='h00000ea3;
    rd_cycle[14597] = 1'b1;  wr_cycle[14597] = 1'b0;  addr_rom[14597]='h00000e04;  wr_data_rom[14597]='h00000000;
    rd_cycle[14598] = 1'b1;  wr_cycle[14598] = 1'b0;  addr_rom[14598]='h0000252c;  wr_data_rom[14598]='h00000000;
    rd_cycle[14599] = 1'b1;  wr_cycle[14599] = 1'b0;  addr_rom[14599]='h00000908;  wr_data_rom[14599]='h00000000;
    rd_cycle[14600] = 1'b0;  wr_cycle[14600] = 1'b1;  addr_rom[14600]='h000024f4;  wr_data_rom[14600]='h000005fc;
    rd_cycle[14601] = 1'b0;  wr_cycle[14601] = 1'b1;  addr_rom[14601]='h0000104c;  wr_data_rom[14601]='h00001bc0;
    rd_cycle[14602] = 1'b0;  wr_cycle[14602] = 1'b1;  addr_rom[14602]='h00000c6c;  wr_data_rom[14602]='h00000bc2;
    rd_cycle[14603] = 1'b1;  wr_cycle[14603] = 1'b0;  addr_rom[14603]='h00003da8;  wr_data_rom[14603]='h00000000;
    rd_cycle[14604] = 1'b1;  wr_cycle[14604] = 1'b0;  addr_rom[14604]='h00003510;  wr_data_rom[14604]='h00000000;
    rd_cycle[14605] = 1'b0;  wr_cycle[14605] = 1'b1;  addr_rom[14605]='h0000037c;  wr_data_rom[14605]='h000030fc;
    rd_cycle[14606] = 1'b0;  wr_cycle[14606] = 1'b1;  addr_rom[14606]='h00000fcc;  wr_data_rom[14606]='h00001db1;
    rd_cycle[14607] = 1'b0;  wr_cycle[14607] = 1'b1;  addr_rom[14607]='h000029ac;  wr_data_rom[14607]='h000036e5;
    rd_cycle[14608] = 1'b0;  wr_cycle[14608] = 1'b1;  addr_rom[14608]='h00002f6c;  wr_data_rom[14608]='h00002941;
    rd_cycle[14609] = 1'b0;  wr_cycle[14609] = 1'b1;  addr_rom[14609]='h00003798;  wr_data_rom[14609]='h00003b9d;
    rd_cycle[14610] = 1'b0;  wr_cycle[14610] = 1'b1;  addr_rom[14610]='h00000ea0;  wr_data_rom[14610]='h000022dc;
    rd_cycle[14611] = 1'b0;  wr_cycle[14611] = 1'b1;  addr_rom[14611]='h00002d28;  wr_data_rom[14611]='h0000025d;
    rd_cycle[14612] = 1'b0;  wr_cycle[14612] = 1'b1;  addr_rom[14612]='h00002d3c;  wr_data_rom[14612]='h000013f4;
    rd_cycle[14613] = 1'b1;  wr_cycle[14613] = 1'b0;  addr_rom[14613]='h0000073c;  wr_data_rom[14613]='h00000000;
    rd_cycle[14614] = 1'b1;  wr_cycle[14614] = 1'b0;  addr_rom[14614]='h00001ee8;  wr_data_rom[14614]='h00000000;
    rd_cycle[14615] = 1'b1;  wr_cycle[14615] = 1'b0;  addr_rom[14615]='h00000658;  wr_data_rom[14615]='h00000000;
    rd_cycle[14616] = 1'b0;  wr_cycle[14616] = 1'b1;  addr_rom[14616]='h00001a04;  wr_data_rom[14616]='h00000667;
    rd_cycle[14617] = 1'b1;  wr_cycle[14617] = 1'b0;  addr_rom[14617]='h00000738;  wr_data_rom[14617]='h00000000;
    rd_cycle[14618] = 1'b0;  wr_cycle[14618] = 1'b1;  addr_rom[14618]='h00001e54;  wr_data_rom[14618]='h000037cc;
    rd_cycle[14619] = 1'b0;  wr_cycle[14619] = 1'b1;  addr_rom[14619]='h000011a0;  wr_data_rom[14619]='h00003b5a;
    rd_cycle[14620] = 1'b0;  wr_cycle[14620] = 1'b1;  addr_rom[14620]='h00001b70;  wr_data_rom[14620]='h00000724;
    rd_cycle[14621] = 1'b0;  wr_cycle[14621] = 1'b1;  addr_rom[14621]='h0000243c;  wr_data_rom[14621]='h00000dc8;
    rd_cycle[14622] = 1'b0;  wr_cycle[14622] = 1'b1;  addr_rom[14622]='h00001d30;  wr_data_rom[14622]='h000018f6;
    rd_cycle[14623] = 1'b0;  wr_cycle[14623] = 1'b1;  addr_rom[14623]='h00001d34;  wr_data_rom[14623]='h00002ee6;
    rd_cycle[14624] = 1'b1;  wr_cycle[14624] = 1'b0;  addr_rom[14624]='h00001e7c;  wr_data_rom[14624]='h00000000;
    rd_cycle[14625] = 1'b0;  wr_cycle[14625] = 1'b1;  addr_rom[14625]='h00002c94;  wr_data_rom[14625]='h00002f8f;
    rd_cycle[14626] = 1'b0;  wr_cycle[14626] = 1'b1;  addr_rom[14626]='h000007d8;  wr_data_rom[14626]='h00003920;
    rd_cycle[14627] = 1'b1;  wr_cycle[14627] = 1'b0;  addr_rom[14627]='h00000a74;  wr_data_rom[14627]='h00000000;
    rd_cycle[14628] = 1'b1;  wr_cycle[14628] = 1'b0;  addr_rom[14628]='h00001f94;  wr_data_rom[14628]='h00000000;
    rd_cycle[14629] = 1'b1;  wr_cycle[14629] = 1'b0;  addr_rom[14629]='h00000c84;  wr_data_rom[14629]='h00000000;
    rd_cycle[14630] = 1'b0;  wr_cycle[14630] = 1'b1;  addr_rom[14630]='h00001560;  wr_data_rom[14630]='h000012f5;
    rd_cycle[14631] = 1'b0;  wr_cycle[14631] = 1'b1;  addr_rom[14631]='h00001260;  wr_data_rom[14631]='h00003e5e;
    rd_cycle[14632] = 1'b1;  wr_cycle[14632] = 1'b0;  addr_rom[14632]='h00002e70;  wr_data_rom[14632]='h00000000;
    rd_cycle[14633] = 1'b1;  wr_cycle[14633] = 1'b0;  addr_rom[14633]='h0000076c;  wr_data_rom[14633]='h00000000;
    rd_cycle[14634] = 1'b0;  wr_cycle[14634] = 1'b1;  addr_rom[14634]='h00003308;  wr_data_rom[14634]='h00003177;
    rd_cycle[14635] = 1'b0;  wr_cycle[14635] = 1'b1;  addr_rom[14635]='h00001da0;  wr_data_rom[14635]='h000020a4;
    rd_cycle[14636] = 1'b0;  wr_cycle[14636] = 1'b1;  addr_rom[14636]='h00002ab0;  wr_data_rom[14636]='h0000107f;
    rd_cycle[14637] = 1'b0;  wr_cycle[14637] = 1'b1;  addr_rom[14637]='h00001a18;  wr_data_rom[14637]='h00002d1d;
    rd_cycle[14638] = 1'b1;  wr_cycle[14638] = 1'b0;  addr_rom[14638]='h00003a48;  wr_data_rom[14638]='h00000000;
    rd_cycle[14639] = 1'b1;  wr_cycle[14639] = 1'b0;  addr_rom[14639]='h00003500;  wr_data_rom[14639]='h00000000;
    rd_cycle[14640] = 1'b1;  wr_cycle[14640] = 1'b0;  addr_rom[14640]='h000030e0;  wr_data_rom[14640]='h00000000;
    rd_cycle[14641] = 1'b1;  wr_cycle[14641] = 1'b0;  addr_rom[14641]='h00002bb4;  wr_data_rom[14641]='h00000000;
    rd_cycle[14642] = 1'b0;  wr_cycle[14642] = 1'b1;  addr_rom[14642]='h00003110;  wr_data_rom[14642]='h000017ca;
    rd_cycle[14643] = 1'b1;  wr_cycle[14643] = 1'b0;  addr_rom[14643]='h00002398;  wr_data_rom[14643]='h00000000;
    rd_cycle[14644] = 1'b0;  wr_cycle[14644] = 1'b1;  addr_rom[14644]='h00003dd8;  wr_data_rom[14644]='h0000239f;
    rd_cycle[14645] = 1'b1;  wr_cycle[14645] = 1'b0;  addr_rom[14645]='h00002e8c;  wr_data_rom[14645]='h00000000;
    rd_cycle[14646] = 1'b1;  wr_cycle[14646] = 1'b0;  addr_rom[14646]='h00001420;  wr_data_rom[14646]='h00000000;
    rd_cycle[14647] = 1'b1;  wr_cycle[14647] = 1'b0;  addr_rom[14647]='h00000e38;  wr_data_rom[14647]='h00000000;
    rd_cycle[14648] = 1'b0;  wr_cycle[14648] = 1'b1;  addr_rom[14648]='h000012a4;  wr_data_rom[14648]='h00001888;
    rd_cycle[14649] = 1'b1;  wr_cycle[14649] = 1'b0;  addr_rom[14649]='h00003274;  wr_data_rom[14649]='h00000000;
    rd_cycle[14650] = 1'b1;  wr_cycle[14650] = 1'b0;  addr_rom[14650]='h00000964;  wr_data_rom[14650]='h00000000;
    rd_cycle[14651] = 1'b0;  wr_cycle[14651] = 1'b1;  addr_rom[14651]='h00003d08;  wr_data_rom[14651]='h00000a34;
    rd_cycle[14652] = 1'b1;  wr_cycle[14652] = 1'b0;  addr_rom[14652]='h000013d0;  wr_data_rom[14652]='h00000000;
    rd_cycle[14653] = 1'b1;  wr_cycle[14653] = 1'b0;  addr_rom[14653]='h000008c8;  wr_data_rom[14653]='h00000000;
    rd_cycle[14654] = 1'b1;  wr_cycle[14654] = 1'b0;  addr_rom[14654]='h00000cf0;  wr_data_rom[14654]='h00000000;
    rd_cycle[14655] = 1'b0;  wr_cycle[14655] = 1'b1;  addr_rom[14655]='h00000230;  wr_data_rom[14655]='h000004a0;
    rd_cycle[14656] = 1'b1;  wr_cycle[14656] = 1'b0;  addr_rom[14656]='h00002ebc;  wr_data_rom[14656]='h00000000;
    rd_cycle[14657] = 1'b1;  wr_cycle[14657] = 1'b0;  addr_rom[14657]='h000011ec;  wr_data_rom[14657]='h00000000;
    rd_cycle[14658] = 1'b0;  wr_cycle[14658] = 1'b1;  addr_rom[14658]='h00001784;  wr_data_rom[14658]='h00003863;
    rd_cycle[14659] = 1'b0;  wr_cycle[14659] = 1'b1;  addr_rom[14659]='h00002054;  wr_data_rom[14659]='h00000708;
    rd_cycle[14660] = 1'b0;  wr_cycle[14660] = 1'b1;  addr_rom[14660]='h000031fc;  wr_data_rom[14660]='h00002232;
    rd_cycle[14661] = 1'b0;  wr_cycle[14661] = 1'b1;  addr_rom[14661]='h00002704;  wr_data_rom[14661]='h00000dc2;
    rd_cycle[14662] = 1'b1;  wr_cycle[14662] = 1'b0;  addr_rom[14662]='h00000404;  wr_data_rom[14662]='h00000000;
    rd_cycle[14663] = 1'b0;  wr_cycle[14663] = 1'b1;  addr_rom[14663]='h00002f38;  wr_data_rom[14663]='h00000386;
    rd_cycle[14664] = 1'b1;  wr_cycle[14664] = 1'b0;  addr_rom[14664]='h00000f94;  wr_data_rom[14664]='h00000000;
    rd_cycle[14665] = 1'b0;  wr_cycle[14665] = 1'b1;  addr_rom[14665]='h00003a88;  wr_data_rom[14665]='h000007dc;
    rd_cycle[14666] = 1'b0;  wr_cycle[14666] = 1'b1;  addr_rom[14666]='h00001738;  wr_data_rom[14666]='h00003f06;
    rd_cycle[14667] = 1'b1;  wr_cycle[14667] = 1'b0;  addr_rom[14667]='h00000760;  wr_data_rom[14667]='h00000000;
    rd_cycle[14668] = 1'b1;  wr_cycle[14668] = 1'b0;  addr_rom[14668]='h00002c18;  wr_data_rom[14668]='h00000000;
    rd_cycle[14669] = 1'b0;  wr_cycle[14669] = 1'b1;  addr_rom[14669]='h00003d78;  wr_data_rom[14669]='h0000070c;
    rd_cycle[14670] = 1'b0;  wr_cycle[14670] = 1'b1;  addr_rom[14670]='h000031d0;  wr_data_rom[14670]='h00003f31;
    rd_cycle[14671] = 1'b1;  wr_cycle[14671] = 1'b0;  addr_rom[14671]='h00003c64;  wr_data_rom[14671]='h00000000;
    rd_cycle[14672] = 1'b1;  wr_cycle[14672] = 1'b0;  addr_rom[14672]='h00003fa4;  wr_data_rom[14672]='h00000000;
    rd_cycle[14673] = 1'b0;  wr_cycle[14673] = 1'b1;  addr_rom[14673]='h00001e34;  wr_data_rom[14673]='h00001a85;
    rd_cycle[14674] = 1'b0;  wr_cycle[14674] = 1'b1;  addr_rom[14674]='h0000229c;  wr_data_rom[14674]='h00003d55;
    rd_cycle[14675] = 1'b0;  wr_cycle[14675] = 1'b1;  addr_rom[14675]='h00002240;  wr_data_rom[14675]='h000012ad;
    rd_cycle[14676] = 1'b1;  wr_cycle[14676] = 1'b0;  addr_rom[14676]='h00000320;  wr_data_rom[14676]='h00000000;
    rd_cycle[14677] = 1'b1;  wr_cycle[14677] = 1'b0;  addr_rom[14677]='h000034ac;  wr_data_rom[14677]='h00000000;
    rd_cycle[14678] = 1'b0;  wr_cycle[14678] = 1'b1;  addr_rom[14678]='h00003740;  wr_data_rom[14678]='h0000378a;
    rd_cycle[14679] = 1'b0;  wr_cycle[14679] = 1'b1;  addr_rom[14679]='h0000309c;  wr_data_rom[14679]='h0000071a;
    rd_cycle[14680] = 1'b0;  wr_cycle[14680] = 1'b1;  addr_rom[14680]='h000026ac;  wr_data_rom[14680]='h0000217a;
    rd_cycle[14681] = 1'b1;  wr_cycle[14681] = 1'b0;  addr_rom[14681]='h00000070;  wr_data_rom[14681]='h00000000;
    rd_cycle[14682] = 1'b1;  wr_cycle[14682] = 1'b0;  addr_rom[14682]='h0000233c;  wr_data_rom[14682]='h00000000;
    rd_cycle[14683] = 1'b0;  wr_cycle[14683] = 1'b1;  addr_rom[14683]='h0000343c;  wr_data_rom[14683]='h0000355d;
    rd_cycle[14684] = 1'b1;  wr_cycle[14684] = 1'b0;  addr_rom[14684]='h000007c8;  wr_data_rom[14684]='h00000000;
    rd_cycle[14685] = 1'b0;  wr_cycle[14685] = 1'b1;  addr_rom[14685]='h00000fa8;  wr_data_rom[14685]='h00002581;
    rd_cycle[14686] = 1'b1;  wr_cycle[14686] = 1'b0;  addr_rom[14686]='h00000928;  wr_data_rom[14686]='h00000000;
    rd_cycle[14687] = 1'b1;  wr_cycle[14687] = 1'b0;  addr_rom[14687]='h00003c74;  wr_data_rom[14687]='h00000000;
    rd_cycle[14688] = 1'b0;  wr_cycle[14688] = 1'b1;  addr_rom[14688]='h000002a4;  wr_data_rom[14688]='h0000372f;
    rd_cycle[14689] = 1'b1;  wr_cycle[14689] = 1'b0;  addr_rom[14689]='h00003180;  wr_data_rom[14689]='h00000000;
    rd_cycle[14690] = 1'b0;  wr_cycle[14690] = 1'b1;  addr_rom[14690]='h00002b24;  wr_data_rom[14690]='h00001037;
    rd_cycle[14691] = 1'b1;  wr_cycle[14691] = 1'b0;  addr_rom[14691]='h00001f48;  wr_data_rom[14691]='h00000000;
    rd_cycle[14692] = 1'b1;  wr_cycle[14692] = 1'b0;  addr_rom[14692]='h00002f58;  wr_data_rom[14692]='h00000000;
    rd_cycle[14693] = 1'b0;  wr_cycle[14693] = 1'b1;  addr_rom[14693]='h00002178;  wr_data_rom[14693]='h0000039d;
    rd_cycle[14694] = 1'b1;  wr_cycle[14694] = 1'b0;  addr_rom[14694]='h00000b88;  wr_data_rom[14694]='h00000000;
    rd_cycle[14695] = 1'b1;  wr_cycle[14695] = 1'b0;  addr_rom[14695]='h00000a8c;  wr_data_rom[14695]='h00000000;
    rd_cycle[14696] = 1'b1;  wr_cycle[14696] = 1'b0;  addr_rom[14696]='h000028ec;  wr_data_rom[14696]='h00000000;
    rd_cycle[14697] = 1'b1;  wr_cycle[14697] = 1'b0;  addr_rom[14697]='h00002a98;  wr_data_rom[14697]='h00000000;
    rd_cycle[14698] = 1'b1;  wr_cycle[14698] = 1'b0;  addr_rom[14698]='h00002944;  wr_data_rom[14698]='h00000000;
    rd_cycle[14699] = 1'b1;  wr_cycle[14699] = 1'b0;  addr_rom[14699]='h00003a4c;  wr_data_rom[14699]='h00000000;
    rd_cycle[14700] = 1'b1;  wr_cycle[14700] = 1'b0;  addr_rom[14700]='h00000780;  wr_data_rom[14700]='h00000000;
    rd_cycle[14701] = 1'b1;  wr_cycle[14701] = 1'b0;  addr_rom[14701]='h00001e60;  wr_data_rom[14701]='h00000000;
    rd_cycle[14702] = 1'b0;  wr_cycle[14702] = 1'b1;  addr_rom[14702]='h00003a54;  wr_data_rom[14702]='h00003dd8;
    rd_cycle[14703] = 1'b0;  wr_cycle[14703] = 1'b1;  addr_rom[14703]='h000014a4;  wr_data_rom[14703]='h00000eb4;
    rd_cycle[14704] = 1'b0;  wr_cycle[14704] = 1'b1;  addr_rom[14704]='h00003ecc;  wr_data_rom[14704]='h00003e87;
    rd_cycle[14705] = 1'b0;  wr_cycle[14705] = 1'b1;  addr_rom[14705]='h000019ec;  wr_data_rom[14705]='h000032ce;
    rd_cycle[14706] = 1'b1;  wr_cycle[14706] = 1'b0;  addr_rom[14706]='h00002370;  wr_data_rom[14706]='h00000000;
    rd_cycle[14707] = 1'b1;  wr_cycle[14707] = 1'b0;  addr_rom[14707]='h0000133c;  wr_data_rom[14707]='h00000000;
    rd_cycle[14708] = 1'b1;  wr_cycle[14708] = 1'b0;  addr_rom[14708]='h00003a18;  wr_data_rom[14708]='h00000000;
    rd_cycle[14709] = 1'b0;  wr_cycle[14709] = 1'b1;  addr_rom[14709]='h000030e8;  wr_data_rom[14709]='h00002041;
    rd_cycle[14710] = 1'b1;  wr_cycle[14710] = 1'b0;  addr_rom[14710]='h00003084;  wr_data_rom[14710]='h00000000;
    rd_cycle[14711] = 1'b0;  wr_cycle[14711] = 1'b1;  addr_rom[14711]='h00000fd0;  wr_data_rom[14711]='h00001876;
    rd_cycle[14712] = 1'b0;  wr_cycle[14712] = 1'b1;  addr_rom[14712]='h000007d4;  wr_data_rom[14712]='h00003050;
    rd_cycle[14713] = 1'b0;  wr_cycle[14713] = 1'b1;  addr_rom[14713]='h00002d38;  wr_data_rom[14713]='h00000c39;
    rd_cycle[14714] = 1'b1;  wr_cycle[14714] = 1'b0;  addr_rom[14714]='h00000bf4;  wr_data_rom[14714]='h00000000;
    rd_cycle[14715] = 1'b1;  wr_cycle[14715] = 1'b0;  addr_rom[14715]='h00003060;  wr_data_rom[14715]='h00000000;
    rd_cycle[14716] = 1'b0;  wr_cycle[14716] = 1'b1;  addr_rom[14716]='h000008d0;  wr_data_rom[14716]='h00001140;
    rd_cycle[14717] = 1'b1;  wr_cycle[14717] = 1'b0;  addr_rom[14717]='h00002128;  wr_data_rom[14717]='h00000000;
    rd_cycle[14718] = 1'b0;  wr_cycle[14718] = 1'b1;  addr_rom[14718]='h000002c0;  wr_data_rom[14718]='h00001088;
    rd_cycle[14719] = 1'b0;  wr_cycle[14719] = 1'b1;  addr_rom[14719]='h00000434;  wr_data_rom[14719]='h00000848;
    rd_cycle[14720] = 1'b1;  wr_cycle[14720] = 1'b0;  addr_rom[14720]='h000002f8;  wr_data_rom[14720]='h00000000;
    rd_cycle[14721] = 1'b1;  wr_cycle[14721] = 1'b0;  addr_rom[14721]='h000021f8;  wr_data_rom[14721]='h00000000;
    rd_cycle[14722] = 1'b0;  wr_cycle[14722] = 1'b1;  addr_rom[14722]='h00002d38;  wr_data_rom[14722]='h0000212c;
    rd_cycle[14723] = 1'b0;  wr_cycle[14723] = 1'b1;  addr_rom[14723]='h00002910;  wr_data_rom[14723]='h0000276f;
    rd_cycle[14724] = 1'b0;  wr_cycle[14724] = 1'b1;  addr_rom[14724]='h00000e90;  wr_data_rom[14724]='h00000a18;
    rd_cycle[14725] = 1'b0;  wr_cycle[14725] = 1'b1;  addr_rom[14725]='h00000450;  wr_data_rom[14725]='h00002ce5;
    rd_cycle[14726] = 1'b1;  wr_cycle[14726] = 1'b0;  addr_rom[14726]='h00003730;  wr_data_rom[14726]='h00000000;
    rd_cycle[14727] = 1'b1;  wr_cycle[14727] = 1'b0;  addr_rom[14727]='h000018e0;  wr_data_rom[14727]='h00000000;
    rd_cycle[14728] = 1'b1;  wr_cycle[14728] = 1'b0;  addr_rom[14728]='h0000145c;  wr_data_rom[14728]='h00000000;
    rd_cycle[14729] = 1'b1;  wr_cycle[14729] = 1'b0;  addr_rom[14729]='h00002020;  wr_data_rom[14729]='h00000000;
    rd_cycle[14730] = 1'b0;  wr_cycle[14730] = 1'b1;  addr_rom[14730]='h000026f0;  wr_data_rom[14730]='h0000098c;
    rd_cycle[14731] = 1'b1;  wr_cycle[14731] = 1'b0;  addr_rom[14731]='h0000276c;  wr_data_rom[14731]='h00000000;
    rd_cycle[14732] = 1'b1;  wr_cycle[14732] = 1'b0;  addr_rom[14732]='h00002f40;  wr_data_rom[14732]='h00000000;
    rd_cycle[14733] = 1'b1;  wr_cycle[14733] = 1'b0;  addr_rom[14733]='h000010c8;  wr_data_rom[14733]='h00000000;
    rd_cycle[14734] = 1'b0;  wr_cycle[14734] = 1'b1;  addr_rom[14734]='h00000944;  wr_data_rom[14734]='h00003bc2;
    rd_cycle[14735] = 1'b0;  wr_cycle[14735] = 1'b1;  addr_rom[14735]='h00002cdc;  wr_data_rom[14735]='h000015e1;
    rd_cycle[14736] = 1'b0;  wr_cycle[14736] = 1'b1;  addr_rom[14736]='h00003998;  wr_data_rom[14736]='h00003d4f;
    rd_cycle[14737] = 1'b0;  wr_cycle[14737] = 1'b1;  addr_rom[14737]='h00000674;  wr_data_rom[14737]='h000025e7;
    rd_cycle[14738] = 1'b1;  wr_cycle[14738] = 1'b0;  addr_rom[14738]='h00000398;  wr_data_rom[14738]='h00000000;
    rd_cycle[14739] = 1'b0;  wr_cycle[14739] = 1'b1;  addr_rom[14739]='h00000c98;  wr_data_rom[14739]='h00003345;
    rd_cycle[14740] = 1'b0;  wr_cycle[14740] = 1'b1;  addr_rom[14740]='h00000988;  wr_data_rom[14740]='h00003c86;
    rd_cycle[14741] = 1'b0;  wr_cycle[14741] = 1'b1;  addr_rom[14741]='h000017b4;  wr_data_rom[14741]='h000001b0;
    rd_cycle[14742] = 1'b0;  wr_cycle[14742] = 1'b1;  addr_rom[14742]='h00001870;  wr_data_rom[14742]='h00000210;
    rd_cycle[14743] = 1'b0;  wr_cycle[14743] = 1'b1;  addr_rom[14743]='h0000340c;  wr_data_rom[14743]='h0000092d;
    rd_cycle[14744] = 1'b0;  wr_cycle[14744] = 1'b1;  addr_rom[14744]='h000015f4;  wr_data_rom[14744]='h00001f48;
    rd_cycle[14745] = 1'b0;  wr_cycle[14745] = 1'b1;  addr_rom[14745]='h00001b40;  wr_data_rom[14745]='h000001af;
    rd_cycle[14746] = 1'b1;  wr_cycle[14746] = 1'b0;  addr_rom[14746]='h000015a4;  wr_data_rom[14746]='h00000000;
    rd_cycle[14747] = 1'b0;  wr_cycle[14747] = 1'b1;  addr_rom[14747]='h00001bec;  wr_data_rom[14747]='h000027a9;
    rd_cycle[14748] = 1'b0;  wr_cycle[14748] = 1'b1;  addr_rom[14748]='h0000149c;  wr_data_rom[14748]='h00000066;
    rd_cycle[14749] = 1'b1;  wr_cycle[14749] = 1'b0;  addr_rom[14749]='h00000f50;  wr_data_rom[14749]='h00000000;
    rd_cycle[14750] = 1'b0;  wr_cycle[14750] = 1'b1;  addr_rom[14750]='h00002d18;  wr_data_rom[14750]='h0000142c;
    rd_cycle[14751] = 1'b1;  wr_cycle[14751] = 1'b0;  addr_rom[14751]='h00003794;  wr_data_rom[14751]='h00000000;
    rd_cycle[14752] = 1'b1;  wr_cycle[14752] = 1'b0;  addr_rom[14752]='h000012b8;  wr_data_rom[14752]='h00000000;
    rd_cycle[14753] = 1'b1;  wr_cycle[14753] = 1'b0;  addr_rom[14753]='h000015b8;  wr_data_rom[14753]='h00000000;
    rd_cycle[14754] = 1'b1;  wr_cycle[14754] = 1'b0;  addr_rom[14754]='h0000007c;  wr_data_rom[14754]='h00000000;
    rd_cycle[14755] = 1'b1;  wr_cycle[14755] = 1'b0;  addr_rom[14755]='h000018ac;  wr_data_rom[14755]='h00000000;
    rd_cycle[14756] = 1'b0;  wr_cycle[14756] = 1'b1;  addr_rom[14756]='h00000f28;  wr_data_rom[14756]='h00001ed1;
    rd_cycle[14757] = 1'b1;  wr_cycle[14757] = 1'b0;  addr_rom[14757]='h00001748;  wr_data_rom[14757]='h00000000;
    rd_cycle[14758] = 1'b0;  wr_cycle[14758] = 1'b1;  addr_rom[14758]='h00000380;  wr_data_rom[14758]='h00000640;
    rd_cycle[14759] = 1'b1;  wr_cycle[14759] = 1'b0;  addr_rom[14759]='h00001ac4;  wr_data_rom[14759]='h00000000;
    rd_cycle[14760] = 1'b0;  wr_cycle[14760] = 1'b1;  addr_rom[14760]='h000011ac;  wr_data_rom[14760]='h00003755;
    rd_cycle[14761] = 1'b0;  wr_cycle[14761] = 1'b1;  addr_rom[14761]='h00002cd4;  wr_data_rom[14761]='h000011ca;
    rd_cycle[14762] = 1'b1;  wr_cycle[14762] = 1'b0;  addr_rom[14762]='h00001730;  wr_data_rom[14762]='h00000000;
    rd_cycle[14763] = 1'b1;  wr_cycle[14763] = 1'b0;  addr_rom[14763]='h00003884;  wr_data_rom[14763]='h00000000;
    rd_cycle[14764] = 1'b1;  wr_cycle[14764] = 1'b0;  addr_rom[14764]='h00001414;  wr_data_rom[14764]='h00000000;
    rd_cycle[14765] = 1'b0;  wr_cycle[14765] = 1'b1;  addr_rom[14765]='h00000c64;  wr_data_rom[14765]='h00003712;
    rd_cycle[14766] = 1'b1;  wr_cycle[14766] = 1'b0;  addr_rom[14766]='h00002e3c;  wr_data_rom[14766]='h00000000;
    rd_cycle[14767] = 1'b1;  wr_cycle[14767] = 1'b0;  addr_rom[14767]='h00001824;  wr_data_rom[14767]='h00000000;
    rd_cycle[14768] = 1'b0;  wr_cycle[14768] = 1'b1;  addr_rom[14768]='h00003058;  wr_data_rom[14768]='h0000124d;
    rd_cycle[14769] = 1'b0;  wr_cycle[14769] = 1'b1;  addr_rom[14769]='h00000a20;  wr_data_rom[14769]='h00002d31;
    rd_cycle[14770] = 1'b0;  wr_cycle[14770] = 1'b1;  addr_rom[14770]='h00000df8;  wr_data_rom[14770]='h00002beb;
    rd_cycle[14771] = 1'b1;  wr_cycle[14771] = 1'b0;  addr_rom[14771]='h000032f0;  wr_data_rom[14771]='h00000000;
    rd_cycle[14772] = 1'b0;  wr_cycle[14772] = 1'b1;  addr_rom[14772]='h000011a4;  wr_data_rom[14772]='h00002743;
    rd_cycle[14773] = 1'b1;  wr_cycle[14773] = 1'b0;  addr_rom[14773]='h0000084c;  wr_data_rom[14773]='h00000000;
    rd_cycle[14774] = 1'b1;  wr_cycle[14774] = 1'b0;  addr_rom[14774]='h00001388;  wr_data_rom[14774]='h00000000;
    rd_cycle[14775] = 1'b0;  wr_cycle[14775] = 1'b1;  addr_rom[14775]='h00002408;  wr_data_rom[14775]='h000009c4;
    rd_cycle[14776] = 1'b1;  wr_cycle[14776] = 1'b0;  addr_rom[14776]='h0000269c;  wr_data_rom[14776]='h00000000;
    rd_cycle[14777] = 1'b0;  wr_cycle[14777] = 1'b1;  addr_rom[14777]='h0000175c;  wr_data_rom[14777]='h00002449;
    rd_cycle[14778] = 1'b0;  wr_cycle[14778] = 1'b1;  addr_rom[14778]='h000008d0;  wr_data_rom[14778]='h000033f5;
    rd_cycle[14779] = 1'b1;  wr_cycle[14779] = 1'b0;  addr_rom[14779]='h00003558;  wr_data_rom[14779]='h00000000;
    rd_cycle[14780] = 1'b0;  wr_cycle[14780] = 1'b1;  addr_rom[14780]='h00001cc8;  wr_data_rom[14780]='h00001b41;
    rd_cycle[14781] = 1'b1;  wr_cycle[14781] = 1'b0;  addr_rom[14781]='h000020a4;  wr_data_rom[14781]='h00000000;
    rd_cycle[14782] = 1'b0;  wr_cycle[14782] = 1'b1;  addr_rom[14782]='h000014c8;  wr_data_rom[14782]='h000030b3;
    rd_cycle[14783] = 1'b0;  wr_cycle[14783] = 1'b1;  addr_rom[14783]='h000023dc;  wr_data_rom[14783]='h00001133;
    rd_cycle[14784] = 1'b1;  wr_cycle[14784] = 1'b0;  addr_rom[14784]='h00001f3c;  wr_data_rom[14784]='h00000000;
    rd_cycle[14785] = 1'b1;  wr_cycle[14785] = 1'b0;  addr_rom[14785]='h000023b0;  wr_data_rom[14785]='h00000000;
    rd_cycle[14786] = 1'b1;  wr_cycle[14786] = 1'b0;  addr_rom[14786]='h00003ba8;  wr_data_rom[14786]='h00000000;
    rd_cycle[14787] = 1'b0;  wr_cycle[14787] = 1'b1;  addr_rom[14787]='h00003aa4;  wr_data_rom[14787]='h00000f3d;
    rd_cycle[14788] = 1'b1;  wr_cycle[14788] = 1'b0;  addr_rom[14788]='h00002aa4;  wr_data_rom[14788]='h00000000;
    rd_cycle[14789] = 1'b0;  wr_cycle[14789] = 1'b1;  addr_rom[14789]='h00002d54;  wr_data_rom[14789]='h00000be8;
    rd_cycle[14790] = 1'b0;  wr_cycle[14790] = 1'b1;  addr_rom[14790]='h00003cf8;  wr_data_rom[14790]='h000033dc;
    rd_cycle[14791] = 1'b0;  wr_cycle[14791] = 1'b1;  addr_rom[14791]='h00001c30;  wr_data_rom[14791]='h00000f00;
    rd_cycle[14792] = 1'b1;  wr_cycle[14792] = 1'b0;  addr_rom[14792]='h00003fac;  wr_data_rom[14792]='h00000000;
    rd_cycle[14793] = 1'b0;  wr_cycle[14793] = 1'b1;  addr_rom[14793]='h00003bfc;  wr_data_rom[14793]='h00000bd2;
    rd_cycle[14794] = 1'b0;  wr_cycle[14794] = 1'b1;  addr_rom[14794]='h00001078;  wr_data_rom[14794]='h0000259a;
    rd_cycle[14795] = 1'b1;  wr_cycle[14795] = 1'b0;  addr_rom[14795]='h00003198;  wr_data_rom[14795]='h00000000;
    rd_cycle[14796] = 1'b0;  wr_cycle[14796] = 1'b1;  addr_rom[14796]='h00002d18;  wr_data_rom[14796]='h000039f0;
    rd_cycle[14797] = 1'b0;  wr_cycle[14797] = 1'b1;  addr_rom[14797]='h000016ac;  wr_data_rom[14797]='h00003f1f;
    rd_cycle[14798] = 1'b1;  wr_cycle[14798] = 1'b0;  addr_rom[14798]='h000011d4;  wr_data_rom[14798]='h00000000;
    rd_cycle[14799] = 1'b1;  wr_cycle[14799] = 1'b0;  addr_rom[14799]='h00001d6c;  wr_data_rom[14799]='h00000000;
    rd_cycle[14800] = 1'b0;  wr_cycle[14800] = 1'b1;  addr_rom[14800]='h00003af8;  wr_data_rom[14800]='h00003dec;
    rd_cycle[14801] = 1'b0;  wr_cycle[14801] = 1'b1;  addr_rom[14801]='h00001d8c;  wr_data_rom[14801]='h0000253d;
    rd_cycle[14802] = 1'b1;  wr_cycle[14802] = 1'b0;  addr_rom[14802]='h000032f0;  wr_data_rom[14802]='h00000000;
    rd_cycle[14803] = 1'b0;  wr_cycle[14803] = 1'b1;  addr_rom[14803]='h000023bc;  wr_data_rom[14803]='h00003266;
    rd_cycle[14804] = 1'b1;  wr_cycle[14804] = 1'b0;  addr_rom[14804]='h00003b84;  wr_data_rom[14804]='h00000000;
    rd_cycle[14805] = 1'b1;  wr_cycle[14805] = 1'b0;  addr_rom[14805]='h00002614;  wr_data_rom[14805]='h00000000;
    rd_cycle[14806] = 1'b0;  wr_cycle[14806] = 1'b1;  addr_rom[14806]='h00002bfc;  wr_data_rom[14806]='h00003044;
    rd_cycle[14807] = 1'b0;  wr_cycle[14807] = 1'b1;  addr_rom[14807]='h00002bd0;  wr_data_rom[14807]='h00001fe6;
    rd_cycle[14808] = 1'b1;  wr_cycle[14808] = 1'b0;  addr_rom[14808]='h00003d34;  wr_data_rom[14808]='h00000000;
    rd_cycle[14809] = 1'b0;  wr_cycle[14809] = 1'b1;  addr_rom[14809]='h000028d0;  wr_data_rom[14809]='h000018fe;
    rd_cycle[14810] = 1'b0;  wr_cycle[14810] = 1'b1;  addr_rom[14810]='h00003c90;  wr_data_rom[14810]='h00002fdf;
    rd_cycle[14811] = 1'b0;  wr_cycle[14811] = 1'b1;  addr_rom[14811]='h000010e0;  wr_data_rom[14811]='h000025bc;
    rd_cycle[14812] = 1'b1;  wr_cycle[14812] = 1'b0;  addr_rom[14812]='h000012e8;  wr_data_rom[14812]='h00000000;
    rd_cycle[14813] = 1'b1;  wr_cycle[14813] = 1'b0;  addr_rom[14813]='h00002958;  wr_data_rom[14813]='h00000000;
    rd_cycle[14814] = 1'b0;  wr_cycle[14814] = 1'b1;  addr_rom[14814]='h000033dc;  wr_data_rom[14814]='h000003f7;
    rd_cycle[14815] = 1'b1;  wr_cycle[14815] = 1'b0;  addr_rom[14815]='h00001c04;  wr_data_rom[14815]='h00000000;
    rd_cycle[14816] = 1'b0;  wr_cycle[14816] = 1'b1;  addr_rom[14816]='h00003604;  wr_data_rom[14816]='h0000372f;
    rd_cycle[14817] = 1'b0;  wr_cycle[14817] = 1'b1;  addr_rom[14817]='h00001bd4;  wr_data_rom[14817]='h0000007d;
    rd_cycle[14818] = 1'b0;  wr_cycle[14818] = 1'b1;  addr_rom[14818]='h00000fc4;  wr_data_rom[14818]='h00003f4a;
    rd_cycle[14819] = 1'b0;  wr_cycle[14819] = 1'b1;  addr_rom[14819]='h0000153c;  wr_data_rom[14819]='h00003c34;
    rd_cycle[14820] = 1'b1;  wr_cycle[14820] = 1'b0;  addr_rom[14820]='h00001918;  wr_data_rom[14820]='h00000000;
    rd_cycle[14821] = 1'b0;  wr_cycle[14821] = 1'b1;  addr_rom[14821]='h00002fd8;  wr_data_rom[14821]='h00000c09;
    rd_cycle[14822] = 1'b1;  wr_cycle[14822] = 1'b0;  addr_rom[14822]='h00000818;  wr_data_rom[14822]='h00000000;
    rd_cycle[14823] = 1'b1;  wr_cycle[14823] = 1'b0;  addr_rom[14823]='h00001f80;  wr_data_rom[14823]='h00000000;
    rd_cycle[14824] = 1'b0;  wr_cycle[14824] = 1'b1;  addr_rom[14824]='h000004a0;  wr_data_rom[14824]='h0000112d;
    rd_cycle[14825] = 1'b1;  wr_cycle[14825] = 1'b0;  addr_rom[14825]='h00001378;  wr_data_rom[14825]='h00000000;
    rd_cycle[14826] = 1'b1;  wr_cycle[14826] = 1'b0;  addr_rom[14826]='h00001ea4;  wr_data_rom[14826]='h00000000;
    rd_cycle[14827] = 1'b1;  wr_cycle[14827] = 1'b0;  addr_rom[14827]='h00003894;  wr_data_rom[14827]='h00000000;
    rd_cycle[14828] = 1'b1;  wr_cycle[14828] = 1'b0;  addr_rom[14828]='h00003b7c;  wr_data_rom[14828]='h00000000;
    rd_cycle[14829] = 1'b1;  wr_cycle[14829] = 1'b0;  addr_rom[14829]='h000032f8;  wr_data_rom[14829]='h00000000;
    rd_cycle[14830] = 1'b0;  wr_cycle[14830] = 1'b1;  addr_rom[14830]='h0000034c;  wr_data_rom[14830]='h00003b29;
    rd_cycle[14831] = 1'b1;  wr_cycle[14831] = 1'b0;  addr_rom[14831]='h00001b48;  wr_data_rom[14831]='h00000000;
    rd_cycle[14832] = 1'b1;  wr_cycle[14832] = 1'b0;  addr_rom[14832]='h00002820;  wr_data_rom[14832]='h00000000;
    rd_cycle[14833] = 1'b1;  wr_cycle[14833] = 1'b0;  addr_rom[14833]='h00003868;  wr_data_rom[14833]='h00000000;
    rd_cycle[14834] = 1'b0;  wr_cycle[14834] = 1'b1;  addr_rom[14834]='h00003814;  wr_data_rom[14834]='h00002b36;
    rd_cycle[14835] = 1'b0;  wr_cycle[14835] = 1'b1;  addr_rom[14835]='h0000059c;  wr_data_rom[14835]='h000021eb;
    rd_cycle[14836] = 1'b1;  wr_cycle[14836] = 1'b0;  addr_rom[14836]='h00003ce4;  wr_data_rom[14836]='h00000000;
    rd_cycle[14837] = 1'b1;  wr_cycle[14837] = 1'b0;  addr_rom[14837]='h00001644;  wr_data_rom[14837]='h00000000;
    rd_cycle[14838] = 1'b1;  wr_cycle[14838] = 1'b0;  addr_rom[14838]='h00003d74;  wr_data_rom[14838]='h00000000;
    rd_cycle[14839] = 1'b1;  wr_cycle[14839] = 1'b0;  addr_rom[14839]='h00000660;  wr_data_rom[14839]='h00000000;
    rd_cycle[14840] = 1'b1;  wr_cycle[14840] = 1'b0;  addr_rom[14840]='h00001d84;  wr_data_rom[14840]='h00000000;
    rd_cycle[14841] = 1'b0;  wr_cycle[14841] = 1'b1;  addr_rom[14841]='h000022e0;  wr_data_rom[14841]='h00003f46;
    rd_cycle[14842] = 1'b1;  wr_cycle[14842] = 1'b0;  addr_rom[14842]='h00003ef0;  wr_data_rom[14842]='h00000000;
    rd_cycle[14843] = 1'b1;  wr_cycle[14843] = 1'b0;  addr_rom[14843]='h000004d4;  wr_data_rom[14843]='h00000000;
    rd_cycle[14844] = 1'b0;  wr_cycle[14844] = 1'b1;  addr_rom[14844]='h00003700;  wr_data_rom[14844]='h00000cc6;
    rd_cycle[14845] = 1'b0;  wr_cycle[14845] = 1'b1;  addr_rom[14845]='h000036f8;  wr_data_rom[14845]='h00002cdc;
    rd_cycle[14846] = 1'b0;  wr_cycle[14846] = 1'b1;  addr_rom[14846]='h00001f14;  wr_data_rom[14846]='h00003fdd;
    rd_cycle[14847] = 1'b1;  wr_cycle[14847] = 1'b0;  addr_rom[14847]='h0000171c;  wr_data_rom[14847]='h00000000;
    rd_cycle[14848] = 1'b1;  wr_cycle[14848] = 1'b0;  addr_rom[14848]='h00001fa8;  wr_data_rom[14848]='h00000000;
    rd_cycle[14849] = 1'b0;  wr_cycle[14849] = 1'b1;  addr_rom[14849]='h0000012c;  wr_data_rom[14849]='h000027a7;
    rd_cycle[14850] = 1'b0;  wr_cycle[14850] = 1'b1;  addr_rom[14850]='h000031b0;  wr_data_rom[14850]='h000012bd;
    rd_cycle[14851] = 1'b1;  wr_cycle[14851] = 1'b0;  addr_rom[14851]='h00002890;  wr_data_rom[14851]='h00000000;
    rd_cycle[14852] = 1'b1;  wr_cycle[14852] = 1'b0;  addr_rom[14852]='h000005a8;  wr_data_rom[14852]='h00000000;
    rd_cycle[14853] = 1'b0;  wr_cycle[14853] = 1'b1;  addr_rom[14853]='h000010f0;  wr_data_rom[14853]='h00001d19;
    rd_cycle[14854] = 1'b1;  wr_cycle[14854] = 1'b0;  addr_rom[14854]='h00002204;  wr_data_rom[14854]='h00000000;
    rd_cycle[14855] = 1'b1;  wr_cycle[14855] = 1'b0;  addr_rom[14855]='h000039a4;  wr_data_rom[14855]='h00000000;
    rd_cycle[14856] = 1'b1;  wr_cycle[14856] = 1'b0;  addr_rom[14856]='h000019f8;  wr_data_rom[14856]='h00000000;
    rd_cycle[14857] = 1'b1;  wr_cycle[14857] = 1'b0;  addr_rom[14857]='h00000d48;  wr_data_rom[14857]='h00000000;
    rd_cycle[14858] = 1'b1;  wr_cycle[14858] = 1'b0;  addr_rom[14858]='h000030dc;  wr_data_rom[14858]='h00000000;
    rd_cycle[14859] = 1'b1;  wr_cycle[14859] = 1'b0;  addr_rom[14859]='h00000164;  wr_data_rom[14859]='h00000000;
    rd_cycle[14860] = 1'b0;  wr_cycle[14860] = 1'b1;  addr_rom[14860]='h00003dfc;  wr_data_rom[14860]='h00001790;
    rd_cycle[14861] = 1'b0;  wr_cycle[14861] = 1'b1;  addr_rom[14861]='h0000098c;  wr_data_rom[14861]='h000026da;
    rd_cycle[14862] = 1'b0;  wr_cycle[14862] = 1'b1;  addr_rom[14862]='h000031cc;  wr_data_rom[14862]='h00001c9d;
    rd_cycle[14863] = 1'b1;  wr_cycle[14863] = 1'b0;  addr_rom[14863]='h00002434;  wr_data_rom[14863]='h00000000;
    rd_cycle[14864] = 1'b0;  wr_cycle[14864] = 1'b1;  addr_rom[14864]='h0000254c;  wr_data_rom[14864]='h000015de;
    rd_cycle[14865] = 1'b0;  wr_cycle[14865] = 1'b1;  addr_rom[14865]='h00003004;  wr_data_rom[14865]='h000011ff;
    rd_cycle[14866] = 1'b0;  wr_cycle[14866] = 1'b1;  addr_rom[14866]='h00001614;  wr_data_rom[14866]='h000029d7;
    rd_cycle[14867] = 1'b0;  wr_cycle[14867] = 1'b1;  addr_rom[14867]='h000029b8;  wr_data_rom[14867]='h00000998;
    rd_cycle[14868] = 1'b0;  wr_cycle[14868] = 1'b1;  addr_rom[14868]='h00002c6c;  wr_data_rom[14868]='h00003ef7;
    rd_cycle[14869] = 1'b0;  wr_cycle[14869] = 1'b1;  addr_rom[14869]='h00003894;  wr_data_rom[14869]='h0000150e;
    rd_cycle[14870] = 1'b1;  wr_cycle[14870] = 1'b0;  addr_rom[14870]='h00002030;  wr_data_rom[14870]='h00000000;
    rd_cycle[14871] = 1'b1;  wr_cycle[14871] = 1'b0;  addr_rom[14871]='h000017c0;  wr_data_rom[14871]='h00000000;
    rd_cycle[14872] = 1'b0;  wr_cycle[14872] = 1'b1;  addr_rom[14872]='h00000f00;  wr_data_rom[14872]='h0000353b;
    rd_cycle[14873] = 1'b0;  wr_cycle[14873] = 1'b1;  addr_rom[14873]='h00003bdc;  wr_data_rom[14873]='h00000c49;
    rd_cycle[14874] = 1'b0;  wr_cycle[14874] = 1'b1;  addr_rom[14874]='h00002e54;  wr_data_rom[14874]='h00000429;
    rd_cycle[14875] = 1'b1;  wr_cycle[14875] = 1'b0;  addr_rom[14875]='h000006fc;  wr_data_rom[14875]='h00000000;
    rd_cycle[14876] = 1'b1;  wr_cycle[14876] = 1'b0;  addr_rom[14876]='h00002fd4;  wr_data_rom[14876]='h00000000;
    rd_cycle[14877] = 1'b0;  wr_cycle[14877] = 1'b1;  addr_rom[14877]='h000025c4;  wr_data_rom[14877]='h00003647;
    rd_cycle[14878] = 1'b1;  wr_cycle[14878] = 1'b0;  addr_rom[14878]='h00002760;  wr_data_rom[14878]='h00000000;
    rd_cycle[14879] = 1'b0;  wr_cycle[14879] = 1'b1;  addr_rom[14879]='h000005f8;  wr_data_rom[14879]='h00000e22;
    rd_cycle[14880] = 1'b1;  wr_cycle[14880] = 1'b0;  addr_rom[14880]='h00001f3c;  wr_data_rom[14880]='h00000000;
    rd_cycle[14881] = 1'b1;  wr_cycle[14881] = 1'b0;  addr_rom[14881]='h00003d00;  wr_data_rom[14881]='h00000000;
    rd_cycle[14882] = 1'b1;  wr_cycle[14882] = 1'b0;  addr_rom[14882]='h00001868;  wr_data_rom[14882]='h00000000;
    rd_cycle[14883] = 1'b0;  wr_cycle[14883] = 1'b1;  addr_rom[14883]='h00000404;  wr_data_rom[14883]='h00001b94;
    rd_cycle[14884] = 1'b0;  wr_cycle[14884] = 1'b1;  addr_rom[14884]='h00001348;  wr_data_rom[14884]='h00003497;
    rd_cycle[14885] = 1'b0;  wr_cycle[14885] = 1'b1;  addr_rom[14885]='h00002d4c;  wr_data_rom[14885]='h000014ba;
    rd_cycle[14886] = 1'b1;  wr_cycle[14886] = 1'b0;  addr_rom[14886]='h00000230;  wr_data_rom[14886]='h00000000;
    rd_cycle[14887] = 1'b0;  wr_cycle[14887] = 1'b1;  addr_rom[14887]='h00003770;  wr_data_rom[14887]='h00003841;
    rd_cycle[14888] = 1'b1;  wr_cycle[14888] = 1'b0;  addr_rom[14888]='h000024dc;  wr_data_rom[14888]='h00000000;
    rd_cycle[14889] = 1'b0;  wr_cycle[14889] = 1'b1;  addr_rom[14889]='h00002124;  wr_data_rom[14889]='h00001478;
    rd_cycle[14890] = 1'b0;  wr_cycle[14890] = 1'b1;  addr_rom[14890]='h00001e18;  wr_data_rom[14890]='h00003a7f;
    rd_cycle[14891] = 1'b1;  wr_cycle[14891] = 1'b0;  addr_rom[14891]='h00000db0;  wr_data_rom[14891]='h00000000;
    rd_cycle[14892] = 1'b0;  wr_cycle[14892] = 1'b1;  addr_rom[14892]='h000028a0;  wr_data_rom[14892]='h00000ea0;
    rd_cycle[14893] = 1'b1;  wr_cycle[14893] = 1'b0;  addr_rom[14893]='h0000138c;  wr_data_rom[14893]='h00000000;
    rd_cycle[14894] = 1'b0;  wr_cycle[14894] = 1'b1;  addr_rom[14894]='h00000b54;  wr_data_rom[14894]='h00002c3b;
    rd_cycle[14895] = 1'b0;  wr_cycle[14895] = 1'b1;  addr_rom[14895]='h00001ab0;  wr_data_rom[14895]='h000000ff;
    rd_cycle[14896] = 1'b1;  wr_cycle[14896] = 1'b0;  addr_rom[14896]='h000008dc;  wr_data_rom[14896]='h00000000;
    rd_cycle[14897] = 1'b0;  wr_cycle[14897] = 1'b1;  addr_rom[14897]='h00002b2c;  wr_data_rom[14897]='h000014b0;
    rd_cycle[14898] = 1'b1;  wr_cycle[14898] = 1'b0;  addr_rom[14898]='h0000235c;  wr_data_rom[14898]='h00000000;
    rd_cycle[14899] = 1'b0;  wr_cycle[14899] = 1'b1;  addr_rom[14899]='h00003350;  wr_data_rom[14899]='h000026ba;
    rd_cycle[14900] = 1'b0;  wr_cycle[14900] = 1'b1;  addr_rom[14900]='h0000292c;  wr_data_rom[14900]='h00001312;
    rd_cycle[14901] = 1'b0;  wr_cycle[14901] = 1'b1;  addr_rom[14901]='h00002f94;  wr_data_rom[14901]='h00003d3b;
    rd_cycle[14902] = 1'b0;  wr_cycle[14902] = 1'b1;  addr_rom[14902]='h00001548;  wr_data_rom[14902]='h0000179d;
    rd_cycle[14903] = 1'b1;  wr_cycle[14903] = 1'b0;  addr_rom[14903]='h00000c44;  wr_data_rom[14903]='h00000000;
    rd_cycle[14904] = 1'b0;  wr_cycle[14904] = 1'b1;  addr_rom[14904]='h00003c64;  wr_data_rom[14904]='h00001914;
    rd_cycle[14905] = 1'b0;  wr_cycle[14905] = 1'b1;  addr_rom[14905]='h00000b18;  wr_data_rom[14905]='h00000be5;
    rd_cycle[14906] = 1'b0;  wr_cycle[14906] = 1'b1;  addr_rom[14906]='h00000fb8;  wr_data_rom[14906]='h00000f2a;
    rd_cycle[14907] = 1'b0;  wr_cycle[14907] = 1'b1;  addr_rom[14907]='h00003af4;  wr_data_rom[14907]='h00000a71;
    rd_cycle[14908] = 1'b1;  wr_cycle[14908] = 1'b0;  addr_rom[14908]='h00002da8;  wr_data_rom[14908]='h00000000;
    rd_cycle[14909] = 1'b0;  wr_cycle[14909] = 1'b1;  addr_rom[14909]='h000013e8;  wr_data_rom[14909]='h000039db;
    rd_cycle[14910] = 1'b1;  wr_cycle[14910] = 1'b0;  addr_rom[14910]='h00002bbc;  wr_data_rom[14910]='h00000000;
    rd_cycle[14911] = 1'b1;  wr_cycle[14911] = 1'b0;  addr_rom[14911]='h00001fd4;  wr_data_rom[14911]='h00000000;
    rd_cycle[14912] = 1'b0;  wr_cycle[14912] = 1'b1;  addr_rom[14912]='h00002080;  wr_data_rom[14912]='h0000112a;
    rd_cycle[14913] = 1'b1;  wr_cycle[14913] = 1'b0;  addr_rom[14913]='h000027b8;  wr_data_rom[14913]='h00000000;
    rd_cycle[14914] = 1'b1;  wr_cycle[14914] = 1'b0;  addr_rom[14914]='h00000fb0;  wr_data_rom[14914]='h00000000;
    rd_cycle[14915] = 1'b1;  wr_cycle[14915] = 1'b0;  addr_rom[14915]='h0000015c;  wr_data_rom[14915]='h00000000;
    rd_cycle[14916] = 1'b0;  wr_cycle[14916] = 1'b1;  addr_rom[14916]='h0000358c;  wr_data_rom[14916]='h000015f7;
    rd_cycle[14917] = 1'b0;  wr_cycle[14917] = 1'b1;  addr_rom[14917]='h00000250;  wr_data_rom[14917]='h00002101;
    rd_cycle[14918] = 1'b1;  wr_cycle[14918] = 1'b0;  addr_rom[14918]='h00001774;  wr_data_rom[14918]='h00000000;
    rd_cycle[14919] = 1'b0;  wr_cycle[14919] = 1'b1;  addr_rom[14919]='h00000874;  wr_data_rom[14919]='h0000209c;
    rd_cycle[14920] = 1'b0;  wr_cycle[14920] = 1'b1;  addr_rom[14920]='h00003544;  wr_data_rom[14920]='h000000fb;
    rd_cycle[14921] = 1'b1;  wr_cycle[14921] = 1'b0;  addr_rom[14921]='h00000008;  wr_data_rom[14921]='h00000000;
    rd_cycle[14922] = 1'b1;  wr_cycle[14922] = 1'b0;  addr_rom[14922]='h000010a8;  wr_data_rom[14922]='h00000000;
    rd_cycle[14923] = 1'b1;  wr_cycle[14923] = 1'b0;  addr_rom[14923]='h00003680;  wr_data_rom[14923]='h00000000;
    rd_cycle[14924] = 1'b0;  wr_cycle[14924] = 1'b1;  addr_rom[14924]='h00002960;  wr_data_rom[14924]='h00000a8a;
    rd_cycle[14925] = 1'b1;  wr_cycle[14925] = 1'b0;  addr_rom[14925]='h0000264c;  wr_data_rom[14925]='h00000000;
    rd_cycle[14926] = 1'b0;  wr_cycle[14926] = 1'b1;  addr_rom[14926]='h000006ec;  wr_data_rom[14926]='h000004a2;
    rd_cycle[14927] = 1'b1;  wr_cycle[14927] = 1'b0;  addr_rom[14927]='h000000c0;  wr_data_rom[14927]='h00000000;
    rd_cycle[14928] = 1'b1;  wr_cycle[14928] = 1'b0;  addr_rom[14928]='h000007b4;  wr_data_rom[14928]='h00000000;
    rd_cycle[14929] = 1'b0;  wr_cycle[14929] = 1'b1;  addr_rom[14929]='h00002844;  wr_data_rom[14929]='h00000133;
    rd_cycle[14930] = 1'b0;  wr_cycle[14930] = 1'b1;  addr_rom[14930]='h000038f4;  wr_data_rom[14930]='h000017e2;
    rd_cycle[14931] = 1'b0;  wr_cycle[14931] = 1'b1;  addr_rom[14931]='h00001eb0;  wr_data_rom[14931]='h000006e7;
    rd_cycle[14932] = 1'b1;  wr_cycle[14932] = 1'b0;  addr_rom[14932]='h00002018;  wr_data_rom[14932]='h00000000;
    rd_cycle[14933] = 1'b0;  wr_cycle[14933] = 1'b1;  addr_rom[14933]='h00000964;  wr_data_rom[14933]='h000037d5;
    rd_cycle[14934] = 1'b0;  wr_cycle[14934] = 1'b1;  addr_rom[14934]='h00001b68;  wr_data_rom[14934]='h000003a8;
    rd_cycle[14935] = 1'b1;  wr_cycle[14935] = 1'b0;  addr_rom[14935]='h00002b60;  wr_data_rom[14935]='h00000000;
    rd_cycle[14936] = 1'b1;  wr_cycle[14936] = 1'b0;  addr_rom[14936]='h00003bf4;  wr_data_rom[14936]='h00000000;
    rd_cycle[14937] = 1'b0;  wr_cycle[14937] = 1'b1;  addr_rom[14937]='h00001254;  wr_data_rom[14937]='h000006a8;
    rd_cycle[14938] = 1'b0;  wr_cycle[14938] = 1'b1;  addr_rom[14938]='h000019d8;  wr_data_rom[14938]='h00003417;
    rd_cycle[14939] = 1'b0;  wr_cycle[14939] = 1'b1;  addr_rom[14939]='h00001dc8;  wr_data_rom[14939]='h00001314;
    rd_cycle[14940] = 1'b1;  wr_cycle[14940] = 1'b0;  addr_rom[14940]='h000018d0;  wr_data_rom[14940]='h00000000;
    rd_cycle[14941] = 1'b1;  wr_cycle[14941] = 1'b0;  addr_rom[14941]='h00002588;  wr_data_rom[14941]='h00000000;
    rd_cycle[14942] = 1'b0;  wr_cycle[14942] = 1'b1;  addr_rom[14942]='h00001de0;  wr_data_rom[14942]='h00001ca4;
    rd_cycle[14943] = 1'b0;  wr_cycle[14943] = 1'b1;  addr_rom[14943]='h00000cf8;  wr_data_rom[14943]='h0000235b;
    rd_cycle[14944] = 1'b1;  wr_cycle[14944] = 1'b0;  addr_rom[14944]='h00003e0c;  wr_data_rom[14944]='h00000000;
    rd_cycle[14945] = 1'b0;  wr_cycle[14945] = 1'b1;  addr_rom[14945]='h0000222c;  wr_data_rom[14945]='h0000048d;
    rd_cycle[14946] = 1'b0;  wr_cycle[14946] = 1'b1;  addr_rom[14946]='h00000e14;  wr_data_rom[14946]='h00001bd9;
    rd_cycle[14947] = 1'b1;  wr_cycle[14947] = 1'b0;  addr_rom[14947]='h000015c4;  wr_data_rom[14947]='h00000000;
    rd_cycle[14948] = 1'b1;  wr_cycle[14948] = 1'b0;  addr_rom[14948]='h000038dc;  wr_data_rom[14948]='h00000000;
    rd_cycle[14949] = 1'b1;  wr_cycle[14949] = 1'b0;  addr_rom[14949]='h00003008;  wr_data_rom[14949]='h00000000;
    rd_cycle[14950] = 1'b0;  wr_cycle[14950] = 1'b1;  addr_rom[14950]='h000007f0;  wr_data_rom[14950]='h00002de4;
    rd_cycle[14951] = 1'b1;  wr_cycle[14951] = 1'b0;  addr_rom[14951]='h00002670;  wr_data_rom[14951]='h00000000;
    rd_cycle[14952] = 1'b1;  wr_cycle[14952] = 1'b0;  addr_rom[14952]='h00002168;  wr_data_rom[14952]='h00000000;
    rd_cycle[14953] = 1'b0;  wr_cycle[14953] = 1'b1;  addr_rom[14953]='h00003874;  wr_data_rom[14953]='h00000ae2;
    rd_cycle[14954] = 1'b1;  wr_cycle[14954] = 1'b0;  addr_rom[14954]='h00000f78;  wr_data_rom[14954]='h00000000;
    rd_cycle[14955] = 1'b1;  wr_cycle[14955] = 1'b0;  addr_rom[14955]='h00001974;  wr_data_rom[14955]='h00000000;
    rd_cycle[14956] = 1'b0;  wr_cycle[14956] = 1'b1;  addr_rom[14956]='h00002584;  wr_data_rom[14956]='h0000348e;
    rd_cycle[14957] = 1'b0;  wr_cycle[14957] = 1'b1;  addr_rom[14957]='h00002704;  wr_data_rom[14957]='h00000317;
    rd_cycle[14958] = 1'b0;  wr_cycle[14958] = 1'b1;  addr_rom[14958]='h00000ecc;  wr_data_rom[14958]='h00000056;
    rd_cycle[14959] = 1'b1;  wr_cycle[14959] = 1'b0;  addr_rom[14959]='h00000c9c;  wr_data_rom[14959]='h00000000;
    rd_cycle[14960] = 1'b1;  wr_cycle[14960] = 1'b0;  addr_rom[14960]='h00003aa8;  wr_data_rom[14960]='h00000000;
    rd_cycle[14961] = 1'b1;  wr_cycle[14961] = 1'b0;  addr_rom[14961]='h000038dc;  wr_data_rom[14961]='h00000000;
    rd_cycle[14962] = 1'b1;  wr_cycle[14962] = 1'b0;  addr_rom[14962]='h00003d3c;  wr_data_rom[14962]='h00000000;
    rd_cycle[14963] = 1'b0;  wr_cycle[14963] = 1'b1;  addr_rom[14963]='h00001ae8;  wr_data_rom[14963]='h00001118;
    rd_cycle[14964] = 1'b0;  wr_cycle[14964] = 1'b1;  addr_rom[14964]='h00000194;  wr_data_rom[14964]='h000007dd;
    rd_cycle[14965] = 1'b0;  wr_cycle[14965] = 1'b1;  addr_rom[14965]='h0000097c;  wr_data_rom[14965]='h0000260a;
    rd_cycle[14966] = 1'b0;  wr_cycle[14966] = 1'b1;  addr_rom[14966]='h000018dc;  wr_data_rom[14966]='h00002721;
    rd_cycle[14967] = 1'b1;  wr_cycle[14967] = 1'b0;  addr_rom[14967]='h000012f0;  wr_data_rom[14967]='h00000000;
    rd_cycle[14968] = 1'b1;  wr_cycle[14968] = 1'b0;  addr_rom[14968]='h00002878;  wr_data_rom[14968]='h00000000;
    rd_cycle[14969] = 1'b0;  wr_cycle[14969] = 1'b1;  addr_rom[14969]='h00000434;  wr_data_rom[14969]='h00003378;
    rd_cycle[14970] = 1'b1;  wr_cycle[14970] = 1'b0;  addr_rom[14970]='h00003c7c;  wr_data_rom[14970]='h00000000;
    rd_cycle[14971] = 1'b0;  wr_cycle[14971] = 1'b1;  addr_rom[14971]='h000006bc;  wr_data_rom[14971]='h00000e01;
    rd_cycle[14972] = 1'b0;  wr_cycle[14972] = 1'b1;  addr_rom[14972]='h00000e04;  wr_data_rom[14972]='h00000ba1;
    rd_cycle[14973] = 1'b1;  wr_cycle[14973] = 1'b0;  addr_rom[14973]='h000024b4;  wr_data_rom[14973]='h00000000;
    rd_cycle[14974] = 1'b1;  wr_cycle[14974] = 1'b0;  addr_rom[14974]='h00000d28;  wr_data_rom[14974]='h00000000;
    rd_cycle[14975] = 1'b0;  wr_cycle[14975] = 1'b1;  addr_rom[14975]='h00002784;  wr_data_rom[14975]='h00002487;
    rd_cycle[14976] = 1'b0;  wr_cycle[14976] = 1'b1;  addr_rom[14976]='h00003a58;  wr_data_rom[14976]='h00001ec5;
    rd_cycle[14977] = 1'b1;  wr_cycle[14977] = 1'b0;  addr_rom[14977]='h00002588;  wr_data_rom[14977]='h00000000;
    rd_cycle[14978] = 1'b1;  wr_cycle[14978] = 1'b0;  addr_rom[14978]='h00003a64;  wr_data_rom[14978]='h00000000;
    rd_cycle[14979] = 1'b1;  wr_cycle[14979] = 1'b0;  addr_rom[14979]='h00003c94;  wr_data_rom[14979]='h00000000;
    rd_cycle[14980] = 1'b0;  wr_cycle[14980] = 1'b1;  addr_rom[14980]='h00001b3c;  wr_data_rom[14980]='h000037b6;
    rd_cycle[14981] = 1'b1;  wr_cycle[14981] = 1'b0;  addr_rom[14981]='h000002b4;  wr_data_rom[14981]='h00000000;
    rd_cycle[14982] = 1'b0;  wr_cycle[14982] = 1'b1;  addr_rom[14982]='h000025a4;  wr_data_rom[14982]='h00001bd0;
    rd_cycle[14983] = 1'b0;  wr_cycle[14983] = 1'b1;  addr_rom[14983]='h00002194;  wr_data_rom[14983]='h00003320;
    rd_cycle[14984] = 1'b0;  wr_cycle[14984] = 1'b1;  addr_rom[14984]='h00000700;  wr_data_rom[14984]='h00000529;
    rd_cycle[14985] = 1'b1;  wr_cycle[14985] = 1'b0;  addr_rom[14985]='h00001aec;  wr_data_rom[14985]='h00000000;
    rd_cycle[14986] = 1'b1;  wr_cycle[14986] = 1'b0;  addr_rom[14986]='h00000bdc;  wr_data_rom[14986]='h00000000;
    rd_cycle[14987] = 1'b0;  wr_cycle[14987] = 1'b1;  addr_rom[14987]='h00000930;  wr_data_rom[14987]='h00000809;
    rd_cycle[14988] = 1'b1;  wr_cycle[14988] = 1'b0;  addr_rom[14988]='h00001528;  wr_data_rom[14988]='h00000000;
    rd_cycle[14989] = 1'b0;  wr_cycle[14989] = 1'b1;  addr_rom[14989]='h000029c0;  wr_data_rom[14989]='h00002b0a;
    rd_cycle[14990] = 1'b0;  wr_cycle[14990] = 1'b1;  addr_rom[14990]='h000022b4;  wr_data_rom[14990]='h00003c4e;
    rd_cycle[14991] = 1'b0;  wr_cycle[14991] = 1'b1;  addr_rom[14991]='h00003450;  wr_data_rom[14991]='h00001cd9;
    rd_cycle[14992] = 1'b1;  wr_cycle[14992] = 1'b0;  addr_rom[14992]='h000022c0;  wr_data_rom[14992]='h00000000;
    rd_cycle[14993] = 1'b0;  wr_cycle[14993] = 1'b1;  addr_rom[14993]='h000034fc;  wr_data_rom[14993]='h00003868;
    rd_cycle[14994] = 1'b0;  wr_cycle[14994] = 1'b1;  addr_rom[14994]='h00003b84;  wr_data_rom[14994]='h00002556;
    rd_cycle[14995] = 1'b1;  wr_cycle[14995] = 1'b0;  addr_rom[14995]='h0000169c;  wr_data_rom[14995]='h00000000;
    rd_cycle[14996] = 1'b0;  wr_cycle[14996] = 1'b1;  addr_rom[14996]='h00001ea0;  wr_data_rom[14996]='h00003804;
    rd_cycle[14997] = 1'b1;  wr_cycle[14997] = 1'b0;  addr_rom[14997]='h00003df4;  wr_data_rom[14997]='h00000000;
    rd_cycle[14998] = 1'b1;  wr_cycle[14998] = 1'b0;  addr_rom[14998]='h000012f8;  wr_data_rom[14998]='h00000000;
    rd_cycle[14999] = 1'b0;  wr_cycle[14999] = 1'b1;  addr_rom[14999]='h000006f8;  wr_data_rom[14999]='h00002083;
    rd_cycle[15000] = 1'b1;  wr_cycle[15000] = 1'b0;  addr_rom[15000]='h00000790;  wr_data_rom[15000]='h00000000;
    rd_cycle[15001] = 1'b0;  wr_cycle[15001] = 1'b1;  addr_rom[15001]='h000016d8;  wr_data_rom[15001]='h00000cd4;
    rd_cycle[15002] = 1'b0;  wr_cycle[15002] = 1'b1;  addr_rom[15002]='h000016d4;  wr_data_rom[15002]='h0000043f;
    rd_cycle[15003] = 1'b0;  wr_cycle[15003] = 1'b1;  addr_rom[15003]='h00002de4;  wr_data_rom[15003]='h00001966;
    rd_cycle[15004] = 1'b0;  wr_cycle[15004] = 1'b1;  addr_rom[15004]='h0000117c;  wr_data_rom[15004]='h00000dd5;
    rd_cycle[15005] = 1'b0;  wr_cycle[15005] = 1'b1;  addr_rom[15005]='h00000bec;  wr_data_rom[15005]='h00003c18;
    rd_cycle[15006] = 1'b0;  wr_cycle[15006] = 1'b1;  addr_rom[15006]='h00002474;  wr_data_rom[15006]='h00001417;
    rd_cycle[15007] = 1'b1;  wr_cycle[15007] = 1'b0;  addr_rom[15007]='h00000af0;  wr_data_rom[15007]='h00000000;
    rd_cycle[15008] = 1'b0;  wr_cycle[15008] = 1'b1;  addr_rom[15008]='h00001bd4;  wr_data_rom[15008]='h00002f0a;
    rd_cycle[15009] = 1'b0;  wr_cycle[15009] = 1'b1;  addr_rom[15009]='h00003298;  wr_data_rom[15009]='h0000114b;
    rd_cycle[15010] = 1'b1;  wr_cycle[15010] = 1'b0;  addr_rom[15010]='h00002cec;  wr_data_rom[15010]='h00000000;
    rd_cycle[15011] = 1'b1;  wr_cycle[15011] = 1'b0;  addr_rom[15011]='h00002f8c;  wr_data_rom[15011]='h00000000;
    rd_cycle[15012] = 1'b0;  wr_cycle[15012] = 1'b1;  addr_rom[15012]='h000039c4;  wr_data_rom[15012]='h00003a8d;
    rd_cycle[15013] = 1'b0;  wr_cycle[15013] = 1'b1;  addr_rom[15013]='h000003e0;  wr_data_rom[15013]='h00003703;
    rd_cycle[15014] = 1'b1;  wr_cycle[15014] = 1'b0;  addr_rom[15014]='h000019f8;  wr_data_rom[15014]='h00000000;
    rd_cycle[15015] = 1'b0;  wr_cycle[15015] = 1'b1;  addr_rom[15015]='h00003dd8;  wr_data_rom[15015]='h00003e83;
    rd_cycle[15016] = 1'b0;  wr_cycle[15016] = 1'b1;  addr_rom[15016]='h00001878;  wr_data_rom[15016]='h00001d12;
    rd_cycle[15017] = 1'b1;  wr_cycle[15017] = 1'b0;  addr_rom[15017]='h000014ac;  wr_data_rom[15017]='h00000000;
    rd_cycle[15018] = 1'b1;  wr_cycle[15018] = 1'b0;  addr_rom[15018]='h000009e8;  wr_data_rom[15018]='h00000000;
    rd_cycle[15019] = 1'b1;  wr_cycle[15019] = 1'b0;  addr_rom[15019]='h00000254;  wr_data_rom[15019]='h00000000;
    rd_cycle[15020] = 1'b1;  wr_cycle[15020] = 1'b0;  addr_rom[15020]='h000030cc;  wr_data_rom[15020]='h00000000;
    rd_cycle[15021] = 1'b0;  wr_cycle[15021] = 1'b1;  addr_rom[15021]='h0000047c;  wr_data_rom[15021]='h00000752;
    rd_cycle[15022] = 1'b0;  wr_cycle[15022] = 1'b1;  addr_rom[15022]='h00003520;  wr_data_rom[15022]='h000027d5;
    rd_cycle[15023] = 1'b0;  wr_cycle[15023] = 1'b1;  addr_rom[15023]='h00001944;  wr_data_rom[15023]='h0000090f;
    rd_cycle[15024] = 1'b1;  wr_cycle[15024] = 1'b0;  addr_rom[15024]='h00001c1c;  wr_data_rom[15024]='h00000000;
    rd_cycle[15025] = 1'b0;  wr_cycle[15025] = 1'b1;  addr_rom[15025]='h00002fa8;  wr_data_rom[15025]='h000017cf;
    rd_cycle[15026] = 1'b0;  wr_cycle[15026] = 1'b1;  addr_rom[15026]='h00003290;  wr_data_rom[15026]='h0000266f;
    rd_cycle[15027] = 1'b0;  wr_cycle[15027] = 1'b1;  addr_rom[15027]='h00001cfc;  wr_data_rom[15027]='h00000f49;
    rd_cycle[15028] = 1'b1;  wr_cycle[15028] = 1'b0;  addr_rom[15028]='h0000254c;  wr_data_rom[15028]='h00000000;
    rd_cycle[15029] = 1'b0;  wr_cycle[15029] = 1'b1;  addr_rom[15029]='h00002080;  wr_data_rom[15029]='h00000398;
    rd_cycle[15030] = 1'b0;  wr_cycle[15030] = 1'b1;  addr_rom[15030]='h000033cc;  wr_data_rom[15030]='h00002b8b;
    rd_cycle[15031] = 1'b1;  wr_cycle[15031] = 1'b0;  addr_rom[15031]='h00001a74;  wr_data_rom[15031]='h00000000;
    rd_cycle[15032] = 1'b1;  wr_cycle[15032] = 1'b0;  addr_rom[15032]='h000018dc;  wr_data_rom[15032]='h00000000;
    rd_cycle[15033] = 1'b0;  wr_cycle[15033] = 1'b1;  addr_rom[15033]='h0000195c;  wr_data_rom[15033]='h0000217f;
    rd_cycle[15034] = 1'b1;  wr_cycle[15034] = 1'b0;  addr_rom[15034]='h00000584;  wr_data_rom[15034]='h00000000;
    rd_cycle[15035] = 1'b1;  wr_cycle[15035] = 1'b0;  addr_rom[15035]='h00000184;  wr_data_rom[15035]='h00000000;
    rd_cycle[15036] = 1'b0;  wr_cycle[15036] = 1'b1;  addr_rom[15036]='h00002498;  wr_data_rom[15036]='h00003ddf;
    rd_cycle[15037] = 1'b0;  wr_cycle[15037] = 1'b1;  addr_rom[15037]='h000025ec;  wr_data_rom[15037]='h0000202e;
    rd_cycle[15038] = 1'b0;  wr_cycle[15038] = 1'b1;  addr_rom[15038]='h00001cb8;  wr_data_rom[15038]='h00001baf;
    rd_cycle[15039] = 1'b0;  wr_cycle[15039] = 1'b1;  addr_rom[15039]='h00003c44;  wr_data_rom[15039]='h00002580;
    rd_cycle[15040] = 1'b1;  wr_cycle[15040] = 1'b0;  addr_rom[15040]='h00002088;  wr_data_rom[15040]='h00000000;
    rd_cycle[15041] = 1'b0;  wr_cycle[15041] = 1'b1;  addr_rom[15041]='h0000290c;  wr_data_rom[15041]='h000025ec;
    rd_cycle[15042] = 1'b1;  wr_cycle[15042] = 1'b0;  addr_rom[15042]='h000037f8;  wr_data_rom[15042]='h00000000;
    rd_cycle[15043] = 1'b1;  wr_cycle[15043] = 1'b0;  addr_rom[15043]='h00001b84;  wr_data_rom[15043]='h00000000;
    rd_cycle[15044] = 1'b1;  wr_cycle[15044] = 1'b0;  addr_rom[15044]='h00002054;  wr_data_rom[15044]='h00000000;
    rd_cycle[15045] = 1'b0;  wr_cycle[15045] = 1'b1;  addr_rom[15045]='h0000344c;  wr_data_rom[15045]='h00002c61;
    rd_cycle[15046] = 1'b0;  wr_cycle[15046] = 1'b1;  addr_rom[15046]='h00001f18;  wr_data_rom[15046]='h00001de6;
    rd_cycle[15047] = 1'b1;  wr_cycle[15047] = 1'b0;  addr_rom[15047]='h00002bd4;  wr_data_rom[15047]='h00000000;
    rd_cycle[15048] = 1'b0;  wr_cycle[15048] = 1'b1;  addr_rom[15048]='h00002d00;  wr_data_rom[15048]='h0000321f;
    rd_cycle[15049] = 1'b0;  wr_cycle[15049] = 1'b1;  addr_rom[15049]='h00002fb8;  wr_data_rom[15049]='h00001648;
    rd_cycle[15050] = 1'b1;  wr_cycle[15050] = 1'b0;  addr_rom[15050]='h00002bac;  wr_data_rom[15050]='h00000000;
    rd_cycle[15051] = 1'b1;  wr_cycle[15051] = 1'b0;  addr_rom[15051]='h00001680;  wr_data_rom[15051]='h00000000;
    rd_cycle[15052] = 1'b1;  wr_cycle[15052] = 1'b0;  addr_rom[15052]='h00002d30;  wr_data_rom[15052]='h00000000;
    rd_cycle[15053] = 1'b1;  wr_cycle[15053] = 1'b0;  addr_rom[15053]='h00000d38;  wr_data_rom[15053]='h00000000;
    rd_cycle[15054] = 1'b1;  wr_cycle[15054] = 1'b0;  addr_rom[15054]='h00003a74;  wr_data_rom[15054]='h00000000;
    rd_cycle[15055] = 1'b0;  wr_cycle[15055] = 1'b1;  addr_rom[15055]='h00001938;  wr_data_rom[15055]='h000036aa;
    rd_cycle[15056] = 1'b1;  wr_cycle[15056] = 1'b0;  addr_rom[15056]='h00003970;  wr_data_rom[15056]='h00000000;
    rd_cycle[15057] = 1'b1;  wr_cycle[15057] = 1'b0;  addr_rom[15057]='h00002c0c;  wr_data_rom[15057]='h00000000;
    rd_cycle[15058] = 1'b0;  wr_cycle[15058] = 1'b1;  addr_rom[15058]='h00000f74;  wr_data_rom[15058]='h000009e9;
    rd_cycle[15059] = 1'b1;  wr_cycle[15059] = 1'b0;  addr_rom[15059]='h00001e54;  wr_data_rom[15059]='h00000000;
    rd_cycle[15060] = 1'b1;  wr_cycle[15060] = 1'b0;  addr_rom[15060]='h00001d70;  wr_data_rom[15060]='h00000000;
    rd_cycle[15061] = 1'b1;  wr_cycle[15061] = 1'b0;  addr_rom[15061]='h000037f4;  wr_data_rom[15061]='h00000000;
    rd_cycle[15062] = 1'b0;  wr_cycle[15062] = 1'b1;  addr_rom[15062]='h000021ec;  wr_data_rom[15062]='h0000193e;
    rd_cycle[15063] = 1'b0;  wr_cycle[15063] = 1'b1;  addr_rom[15063]='h00001c64;  wr_data_rom[15063]='h000006b7;
    rd_cycle[15064] = 1'b0;  wr_cycle[15064] = 1'b1;  addr_rom[15064]='h00000740;  wr_data_rom[15064]='h000028a4;
    rd_cycle[15065] = 1'b0;  wr_cycle[15065] = 1'b1;  addr_rom[15065]='h000025b0;  wr_data_rom[15065]='h00001be7;
    rd_cycle[15066] = 1'b0;  wr_cycle[15066] = 1'b1;  addr_rom[15066]='h00001130;  wr_data_rom[15066]='h00003001;
    rd_cycle[15067] = 1'b0;  wr_cycle[15067] = 1'b1;  addr_rom[15067]='h00000668;  wr_data_rom[15067]='h000024eb;
    rd_cycle[15068] = 1'b1;  wr_cycle[15068] = 1'b0;  addr_rom[15068]='h00002bd8;  wr_data_rom[15068]='h00000000;
    rd_cycle[15069] = 1'b0;  wr_cycle[15069] = 1'b1;  addr_rom[15069]='h00001d94;  wr_data_rom[15069]='h00001957;
    rd_cycle[15070] = 1'b1;  wr_cycle[15070] = 1'b0;  addr_rom[15070]='h000034fc;  wr_data_rom[15070]='h00000000;
    rd_cycle[15071] = 1'b1;  wr_cycle[15071] = 1'b0;  addr_rom[15071]='h00001f48;  wr_data_rom[15071]='h00000000;
    rd_cycle[15072] = 1'b0;  wr_cycle[15072] = 1'b1;  addr_rom[15072]='h00003a1c;  wr_data_rom[15072]='h000008b5;
    rd_cycle[15073] = 1'b1;  wr_cycle[15073] = 1'b0;  addr_rom[15073]='h00000260;  wr_data_rom[15073]='h00000000;
    rd_cycle[15074] = 1'b1;  wr_cycle[15074] = 1'b0;  addr_rom[15074]='h00000628;  wr_data_rom[15074]='h00000000;
    rd_cycle[15075] = 1'b0;  wr_cycle[15075] = 1'b1;  addr_rom[15075]='h00001c54;  wr_data_rom[15075]='h00003afd;
    rd_cycle[15076] = 1'b0;  wr_cycle[15076] = 1'b1;  addr_rom[15076]='h000009c8;  wr_data_rom[15076]='h00001544;
    rd_cycle[15077] = 1'b1;  wr_cycle[15077] = 1'b0;  addr_rom[15077]='h0000136c;  wr_data_rom[15077]='h00000000;
    rd_cycle[15078] = 1'b1;  wr_cycle[15078] = 1'b0;  addr_rom[15078]='h00003a94;  wr_data_rom[15078]='h00000000;
    rd_cycle[15079] = 1'b1;  wr_cycle[15079] = 1'b0;  addr_rom[15079]='h00001a48;  wr_data_rom[15079]='h00000000;
    rd_cycle[15080] = 1'b0;  wr_cycle[15080] = 1'b1;  addr_rom[15080]='h00000198;  wr_data_rom[15080]='h00000cb2;
    rd_cycle[15081] = 1'b0;  wr_cycle[15081] = 1'b1;  addr_rom[15081]='h00003734;  wr_data_rom[15081]='h00000b62;
    rd_cycle[15082] = 1'b1;  wr_cycle[15082] = 1'b0;  addr_rom[15082]='h000023bc;  wr_data_rom[15082]='h00000000;
    rd_cycle[15083] = 1'b1;  wr_cycle[15083] = 1'b0;  addr_rom[15083]='h00002e34;  wr_data_rom[15083]='h00000000;
    rd_cycle[15084] = 1'b1;  wr_cycle[15084] = 1'b0;  addr_rom[15084]='h000005ac;  wr_data_rom[15084]='h00000000;
    rd_cycle[15085] = 1'b0;  wr_cycle[15085] = 1'b1;  addr_rom[15085]='h00000e44;  wr_data_rom[15085]='h00001ec5;
    rd_cycle[15086] = 1'b1;  wr_cycle[15086] = 1'b0;  addr_rom[15086]='h00003644;  wr_data_rom[15086]='h00000000;
    rd_cycle[15087] = 1'b1;  wr_cycle[15087] = 1'b0;  addr_rom[15087]='h000023fc;  wr_data_rom[15087]='h00000000;
    rd_cycle[15088] = 1'b0;  wr_cycle[15088] = 1'b1;  addr_rom[15088]='h00000274;  wr_data_rom[15088]='h0000344c;
    rd_cycle[15089] = 1'b1;  wr_cycle[15089] = 1'b0;  addr_rom[15089]='h00003474;  wr_data_rom[15089]='h00000000;
    rd_cycle[15090] = 1'b0;  wr_cycle[15090] = 1'b1;  addr_rom[15090]='h00003300;  wr_data_rom[15090]='h00002abb;
    rd_cycle[15091] = 1'b0;  wr_cycle[15091] = 1'b1;  addr_rom[15091]='h00003994;  wr_data_rom[15091]='h00001070;
    rd_cycle[15092] = 1'b0;  wr_cycle[15092] = 1'b1;  addr_rom[15092]='h00003560;  wr_data_rom[15092]='h000023ae;
    rd_cycle[15093] = 1'b1;  wr_cycle[15093] = 1'b0;  addr_rom[15093]='h000005dc;  wr_data_rom[15093]='h00000000;
    rd_cycle[15094] = 1'b0;  wr_cycle[15094] = 1'b1;  addr_rom[15094]='h00000b84;  wr_data_rom[15094]='h000021ca;
    rd_cycle[15095] = 1'b1;  wr_cycle[15095] = 1'b0;  addr_rom[15095]='h00001dcc;  wr_data_rom[15095]='h00000000;
    rd_cycle[15096] = 1'b0;  wr_cycle[15096] = 1'b1;  addr_rom[15096]='h00003e04;  wr_data_rom[15096]='h0000263d;
    rd_cycle[15097] = 1'b0;  wr_cycle[15097] = 1'b1;  addr_rom[15097]='h00001ae8;  wr_data_rom[15097]='h000034a8;
    rd_cycle[15098] = 1'b1;  wr_cycle[15098] = 1'b0;  addr_rom[15098]='h00003a78;  wr_data_rom[15098]='h00000000;
    rd_cycle[15099] = 1'b0;  wr_cycle[15099] = 1'b1;  addr_rom[15099]='h00003e84;  wr_data_rom[15099]='h00000238;
    rd_cycle[15100] = 1'b0;  wr_cycle[15100] = 1'b1;  addr_rom[15100]='h00001518;  wr_data_rom[15100]='h000031c7;
    rd_cycle[15101] = 1'b1;  wr_cycle[15101] = 1'b0;  addr_rom[15101]='h0000037c;  wr_data_rom[15101]='h00000000;
    rd_cycle[15102] = 1'b1;  wr_cycle[15102] = 1'b0;  addr_rom[15102]='h00000bc4;  wr_data_rom[15102]='h00000000;
    rd_cycle[15103] = 1'b0;  wr_cycle[15103] = 1'b1;  addr_rom[15103]='h00002d5c;  wr_data_rom[15103]='h0000288b;
    rd_cycle[15104] = 1'b1;  wr_cycle[15104] = 1'b0;  addr_rom[15104]='h00000a40;  wr_data_rom[15104]='h00000000;
    rd_cycle[15105] = 1'b0;  wr_cycle[15105] = 1'b1;  addr_rom[15105]='h000036d8;  wr_data_rom[15105]='h00003d02;
    rd_cycle[15106] = 1'b0;  wr_cycle[15106] = 1'b1;  addr_rom[15106]='h000011a4;  wr_data_rom[15106]='h00000bf5;
    rd_cycle[15107] = 1'b0;  wr_cycle[15107] = 1'b1;  addr_rom[15107]='h00002e50;  wr_data_rom[15107]='h00001be3;
    rd_cycle[15108] = 1'b1;  wr_cycle[15108] = 1'b0;  addr_rom[15108]='h000001e0;  wr_data_rom[15108]='h00000000;
    rd_cycle[15109] = 1'b1;  wr_cycle[15109] = 1'b0;  addr_rom[15109]='h00003ba0;  wr_data_rom[15109]='h00000000;
    rd_cycle[15110] = 1'b0;  wr_cycle[15110] = 1'b1;  addr_rom[15110]='h00002900;  wr_data_rom[15110]='h00003277;
    rd_cycle[15111] = 1'b0;  wr_cycle[15111] = 1'b1;  addr_rom[15111]='h00001b24;  wr_data_rom[15111]='h00002e68;
    rd_cycle[15112] = 1'b0;  wr_cycle[15112] = 1'b1;  addr_rom[15112]='h00002f78;  wr_data_rom[15112]='h00000cc9;
    rd_cycle[15113] = 1'b1;  wr_cycle[15113] = 1'b0;  addr_rom[15113]='h00002608;  wr_data_rom[15113]='h00000000;
    rd_cycle[15114] = 1'b1;  wr_cycle[15114] = 1'b0;  addr_rom[15114]='h000032c4;  wr_data_rom[15114]='h00000000;
    rd_cycle[15115] = 1'b1;  wr_cycle[15115] = 1'b0;  addr_rom[15115]='h000024a8;  wr_data_rom[15115]='h00000000;
    rd_cycle[15116] = 1'b0;  wr_cycle[15116] = 1'b1;  addr_rom[15116]='h00000194;  wr_data_rom[15116]='h000033cc;
    rd_cycle[15117] = 1'b1;  wr_cycle[15117] = 1'b0;  addr_rom[15117]='h00000634;  wr_data_rom[15117]='h00000000;
    rd_cycle[15118] = 1'b1;  wr_cycle[15118] = 1'b0;  addr_rom[15118]='h00000300;  wr_data_rom[15118]='h00000000;
    rd_cycle[15119] = 1'b0;  wr_cycle[15119] = 1'b1;  addr_rom[15119]='h00000bd4;  wr_data_rom[15119]='h00002223;
    rd_cycle[15120] = 1'b0;  wr_cycle[15120] = 1'b1;  addr_rom[15120]='h00003960;  wr_data_rom[15120]='h000017f7;
    rd_cycle[15121] = 1'b1;  wr_cycle[15121] = 1'b0;  addr_rom[15121]='h00001c9c;  wr_data_rom[15121]='h00000000;
    rd_cycle[15122] = 1'b0;  wr_cycle[15122] = 1'b1;  addr_rom[15122]='h00001b6c;  wr_data_rom[15122]='h0000347e;
    rd_cycle[15123] = 1'b0;  wr_cycle[15123] = 1'b1;  addr_rom[15123]='h00001028;  wr_data_rom[15123]='h0000325c;
    rd_cycle[15124] = 1'b1;  wr_cycle[15124] = 1'b0;  addr_rom[15124]='h00000cf0;  wr_data_rom[15124]='h00000000;
    rd_cycle[15125] = 1'b1;  wr_cycle[15125] = 1'b0;  addr_rom[15125]='h00000434;  wr_data_rom[15125]='h00000000;
    rd_cycle[15126] = 1'b0;  wr_cycle[15126] = 1'b1;  addr_rom[15126]='h00003afc;  wr_data_rom[15126]='h00003870;
    rd_cycle[15127] = 1'b0;  wr_cycle[15127] = 1'b1;  addr_rom[15127]='h0000299c;  wr_data_rom[15127]='h00002343;
    rd_cycle[15128] = 1'b0;  wr_cycle[15128] = 1'b1;  addr_rom[15128]='h00000610;  wr_data_rom[15128]='h00003ff3;
    rd_cycle[15129] = 1'b1;  wr_cycle[15129] = 1'b0;  addr_rom[15129]='h000019a8;  wr_data_rom[15129]='h00000000;
    rd_cycle[15130] = 1'b0;  wr_cycle[15130] = 1'b1;  addr_rom[15130]='h00001018;  wr_data_rom[15130]='h000002be;
    rd_cycle[15131] = 1'b0;  wr_cycle[15131] = 1'b1;  addr_rom[15131]='h00001470;  wr_data_rom[15131]='h00000bd0;
    rd_cycle[15132] = 1'b1;  wr_cycle[15132] = 1'b0;  addr_rom[15132]='h00001d94;  wr_data_rom[15132]='h00000000;
    rd_cycle[15133] = 1'b1;  wr_cycle[15133] = 1'b0;  addr_rom[15133]='h000032d4;  wr_data_rom[15133]='h00000000;
    rd_cycle[15134] = 1'b1;  wr_cycle[15134] = 1'b0;  addr_rom[15134]='h0000055c;  wr_data_rom[15134]='h00000000;
    rd_cycle[15135] = 1'b1;  wr_cycle[15135] = 1'b0;  addr_rom[15135]='h00002c88;  wr_data_rom[15135]='h00000000;
    rd_cycle[15136] = 1'b1;  wr_cycle[15136] = 1'b0;  addr_rom[15136]='h00001304;  wr_data_rom[15136]='h00000000;
    rd_cycle[15137] = 1'b1;  wr_cycle[15137] = 1'b0;  addr_rom[15137]='h00003c74;  wr_data_rom[15137]='h00000000;
    rd_cycle[15138] = 1'b1;  wr_cycle[15138] = 1'b0;  addr_rom[15138]='h00001c68;  wr_data_rom[15138]='h00000000;
    rd_cycle[15139] = 1'b1;  wr_cycle[15139] = 1'b0;  addr_rom[15139]='h00003304;  wr_data_rom[15139]='h00000000;
    rd_cycle[15140] = 1'b1;  wr_cycle[15140] = 1'b0;  addr_rom[15140]='h00003eb4;  wr_data_rom[15140]='h00000000;
    rd_cycle[15141] = 1'b1;  wr_cycle[15141] = 1'b0;  addr_rom[15141]='h00001a4c;  wr_data_rom[15141]='h00000000;
    rd_cycle[15142] = 1'b1;  wr_cycle[15142] = 1'b0;  addr_rom[15142]='h00003418;  wr_data_rom[15142]='h00000000;
    rd_cycle[15143] = 1'b0;  wr_cycle[15143] = 1'b1;  addr_rom[15143]='h000002e4;  wr_data_rom[15143]='h0000090f;
    rd_cycle[15144] = 1'b1;  wr_cycle[15144] = 1'b0;  addr_rom[15144]='h00003b2c;  wr_data_rom[15144]='h00000000;
    rd_cycle[15145] = 1'b1;  wr_cycle[15145] = 1'b0;  addr_rom[15145]='h00002e94;  wr_data_rom[15145]='h00000000;
    rd_cycle[15146] = 1'b1;  wr_cycle[15146] = 1'b0;  addr_rom[15146]='h000017fc;  wr_data_rom[15146]='h00000000;
    rd_cycle[15147] = 1'b0;  wr_cycle[15147] = 1'b1;  addr_rom[15147]='h0000168c;  wr_data_rom[15147]='h000033bc;
    rd_cycle[15148] = 1'b1;  wr_cycle[15148] = 1'b0;  addr_rom[15148]='h00000b24;  wr_data_rom[15148]='h00000000;
    rd_cycle[15149] = 1'b1;  wr_cycle[15149] = 1'b0;  addr_rom[15149]='h000008a4;  wr_data_rom[15149]='h00000000;
    rd_cycle[15150] = 1'b0;  wr_cycle[15150] = 1'b1;  addr_rom[15150]='h00002ff4;  wr_data_rom[15150]='h000032cc;
    rd_cycle[15151] = 1'b1;  wr_cycle[15151] = 1'b0;  addr_rom[15151]='h00000a0c;  wr_data_rom[15151]='h00000000;
    rd_cycle[15152] = 1'b0;  wr_cycle[15152] = 1'b1;  addr_rom[15152]='h00001430;  wr_data_rom[15152]='h00003114;
    rd_cycle[15153] = 1'b1;  wr_cycle[15153] = 1'b0;  addr_rom[15153]='h000034cc;  wr_data_rom[15153]='h00000000;
    rd_cycle[15154] = 1'b0;  wr_cycle[15154] = 1'b1;  addr_rom[15154]='h00001060;  wr_data_rom[15154]='h00003dac;
    rd_cycle[15155] = 1'b1;  wr_cycle[15155] = 1'b0;  addr_rom[15155]='h00003a38;  wr_data_rom[15155]='h00000000;
    rd_cycle[15156] = 1'b1;  wr_cycle[15156] = 1'b0;  addr_rom[15156]='h00000cb8;  wr_data_rom[15156]='h00000000;
    rd_cycle[15157] = 1'b0;  wr_cycle[15157] = 1'b1;  addr_rom[15157]='h00002a08;  wr_data_rom[15157]='h000031c2;
    rd_cycle[15158] = 1'b1;  wr_cycle[15158] = 1'b0;  addr_rom[15158]='h000005c0;  wr_data_rom[15158]='h00000000;
    rd_cycle[15159] = 1'b0;  wr_cycle[15159] = 1'b1;  addr_rom[15159]='h00000528;  wr_data_rom[15159]='h0000222c;
    rd_cycle[15160] = 1'b0;  wr_cycle[15160] = 1'b1;  addr_rom[15160]='h0000288c;  wr_data_rom[15160]='h00001d76;
    rd_cycle[15161] = 1'b1;  wr_cycle[15161] = 1'b0;  addr_rom[15161]='h000004b0;  wr_data_rom[15161]='h00000000;
    rd_cycle[15162] = 1'b0;  wr_cycle[15162] = 1'b1;  addr_rom[15162]='h00000278;  wr_data_rom[15162]='h00002bf2;
    rd_cycle[15163] = 1'b0;  wr_cycle[15163] = 1'b1;  addr_rom[15163]='h00002614;  wr_data_rom[15163]='h000003b7;
    rd_cycle[15164] = 1'b1;  wr_cycle[15164] = 1'b0;  addr_rom[15164]='h00001698;  wr_data_rom[15164]='h00000000;
    rd_cycle[15165] = 1'b0;  wr_cycle[15165] = 1'b1;  addr_rom[15165]='h000036d8;  wr_data_rom[15165]='h000026c4;
    rd_cycle[15166] = 1'b0;  wr_cycle[15166] = 1'b1;  addr_rom[15166]='h00000d2c;  wr_data_rom[15166]='h000008f8;
    rd_cycle[15167] = 1'b1;  wr_cycle[15167] = 1'b0;  addr_rom[15167]='h000032f8;  wr_data_rom[15167]='h00000000;
    rd_cycle[15168] = 1'b1;  wr_cycle[15168] = 1'b0;  addr_rom[15168]='h00003aac;  wr_data_rom[15168]='h00000000;
    rd_cycle[15169] = 1'b1;  wr_cycle[15169] = 1'b0;  addr_rom[15169]='h000019b4;  wr_data_rom[15169]='h00000000;
    rd_cycle[15170] = 1'b0;  wr_cycle[15170] = 1'b1;  addr_rom[15170]='h00000090;  wr_data_rom[15170]='h00002b8e;
    rd_cycle[15171] = 1'b1;  wr_cycle[15171] = 1'b0;  addr_rom[15171]='h0000343c;  wr_data_rom[15171]='h00000000;
    rd_cycle[15172] = 1'b1;  wr_cycle[15172] = 1'b0;  addr_rom[15172]='h000000e8;  wr_data_rom[15172]='h00000000;
    rd_cycle[15173] = 1'b1;  wr_cycle[15173] = 1'b0;  addr_rom[15173]='h00000264;  wr_data_rom[15173]='h00000000;
    rd_cycle[15174] = 1'b0;  wr_cycle[15174] = 1'b1;  addr_rom[15174]='h00000af8;  wr_data_rom[15174]='h00002544;
    rd_cycle[15175] = 1'b0;  wr_cycle[15175] = 1'b1;  addr_rom[15175]='h00001580;  wr_data_rom[15175]='h00001e9f;
    rd_cycle[15176] = 1'b0;  wr_cycle[15176] = 1'b1;  addr_rom[15176]='h000006f8;  wr_data_rom[15176]='h00000c99;
    rd_cycle[15177] = 1'b1;  wr_cycle[15177] = 1'b0;  addr_rom[15177]='h00002974;  wr_data_rom[15177]='h00000000;
    rd_cycle[15178] = 1'b0;  wr_cycle[15178] = 1'b1;  addr_rom[15178]='h0000142c;  wr_data_rom[15178]='h00000fbd;
    rd_cycle[15179] = 1'b1;  wr_cycle[15179] = 1'b0;  addr_rom[15179]='h00000f04;  wr_data_rom[15179]='h00000000;
    rd_cycle[15180] = 1'b1;  wr_cycle[15180] = 1'b0;  addr_rom[15180]='h00001c34;  wr_data_rom[15180]='h00000000;
    rd_cycle[15181] = 1'b1;  wr_cycle[15181] = 1'b0;  addr_rom[15181]='h000027fc;  wr_data_rom[15181]='h00000000;
    rd_cycle[15182] = 1'b1;  wr_cycle[15182] = 1'b0;  addr_rom[15182]='h000027d8;  wr_data_rom[15182]='h00000000;
    rd_cycle[15183] = 1'b1;  wr_cycle[15183] = 1'b0;  addr_rom[15183]='h000000c8;  wr_data_rom[15183]='h00000000;
    rd_cycle[15184] = 1'b1;  wr_cycle[15184] = 1'b0;  addr_rom[15184]='h000013c0;  wr_data_rom[15184]='h00000000;
    rd_cycle[15185] = 1'b0;  wr_cycle[15185] = 1'b1;  addr_rom[15185]='h00001f08;  wr_data_rom[15185]='h0000000d;
    rd_cycle[15186] = 1'b1;  wr_cycle[15186] = 1'b0;  addr_rom[15186]='h000012f8;  wr_data_rom[15186]='h00000000;
    rd_cycle[15187] = 1'b1;  wr_cycle[15187] = 1'b0;  addr_rom[15187]='h00002524;  wr_data_rom[15187]='h00000000;
    rd_cycle[15188] = 1'b0;  wr_cycle[15188] = 1'b1;  addr_rom[15188]='h000029e8;  wr_data_rom[15188]='h00003fac;
    rd_cycle[15189] = 1'b0;  wr_cycle[15189] = 1'b1;  addr_rom[15189]='h000022ec;  wr_data_rom[15189]='h000027b2;
    rd_cycle[15190] = 1'b0;  wr_cycle[15190] = 1'b1;  addr_rom[15190]='h000017c4;  wr_data_rom[15190]='h000016e7;
    rd_cycle[15191] = 1'b0;  wr_cycle[15191] = 1'b1;  addr_rom[15191]='h00003ff8;  wr_data_rom[15191]='h00002176;
    rd_cycle[15192] = 1'b1;  wr_cycle[15192] = 1'b0;  addr_rom[15192]='h00003d70;  wr_data_rom[15192]='h00000000;
    rd_cycle[15193] = 1'b1;  wr_cycle[15193] = 1'b0;  addr_rom[15193]='h00003b60;  wr_data_rom[15193]='h00000000;
    rd_cycle[15194] = 1'b0;  wr_cycle[15194] = 1'b1;  addr_rom[15194]='h00000538;  wr_data_rom[15194]='h0000223d;
    rd_cycle[15195] = 1'b0;  wr_cycle[15195] = 1'b1;  addr_rom[15195]='h00003888;  wr_data_rom[15195]='h0000253e;
    rd_cycle[15196] = 1'b0;  wr_cycle[15196] = 1'b1;  addr_rom[15196]='h0000166c;  wr_data_rom[15196]='h000016d3;
    rd_cycle[15197] = 1'b1;  wr_cycle[15197] = 1'b0;  addr_rom[15197]='h00002648;  wr_data_rom[15197]='h00000000;
    rd_cycle[15198] = 1'b0;  wr_cycle[15198] = 1'b1;  addr_rom[15198]='h000020ec;  wr_data_rom[15198]='h00003aea;
    rd_cycle[15199] = 1'b1;  wr_cycle[15199] = 1'b0;  addr_rom[15199]='h00003034;  wr_data_rom[15199]='h00000000;
    rd_cycle[15200] = 1'b1;  wr_cycle[15200] = 1'b0;  addr_rom[15200]='h000038f4;  wr_data_rom[15200]='h00000000;
    rd_cycle[15201] = 1'b1;  wr_cycle[15201] = 1'b0;  addr_rom[15201]='h00000650;  wr_data_rom[15201]='h00000000;
    rd_cycle[15202] = 1'b1;  wr_cycle[15202] = 1'b0;  addr_rom[15202]='h0000130c;  wr_data_rom[15202]='h00000000;
    rd_cycle[15203] = 1'b0;  wr_cycle[15203] = 1'b1;  addr_rom[15203]='h00002fa4;  wr_data_rom[15203]='h000013e0;
    rd_cycle[15204] = 1'b0;  wr_cycle[15204] = 1'b1;  addr_rom[15204]='h00001450;  wr_data_rom[15204]='h00001c5b;
    rd_cycle[15205] = 1'b0;  wr_cycle[15205] = 1'b1;  addr_rom[15205]='h00000e64;  wr_data_rom[15205]='h00002295;
    rd_cycle[15206] = 1'b1;  wr_cycle[15206] = 1'b0;  addr_rom[15206]='h00000a74;  wr_data_rom[15206]='h00000000;
    rd_cycle[15207] = 1'b0;  wr_cycle[15207] = 1'b1;  addr_rom[15207]='h00000014;  wr_data_rom[15207]='h00000fc1;
    rd_cycle[15208] = 1'b0;  wr_cycle[15208] = 1'b1;  addr_rom[15208]='h00002504;  wr_data_rom[15208]='h000016f7;
    rd_cycle[15209] = 1'b1;  wr_cycle[15209] = 1'b0;  addr_rom[15209]='h000002a4;  wr_data_rom[15209]='h00000000;
    rd_cycle[15210] = 1'b0;  wr_cycle[15210] = 1'b1;  addr_rom[15210]='h00001240;  wr_data_rom[15210]='h000003ae;
    rd_cycle[15211] = 1'b0;  wr_cycle[15211] = 1'b1;  addr_rom[15211]='h000025d8;  wr_data_rom[15211]='h000035f7;
    rd_cycle[15212] = 1'b0;  wr_cycle[15212] = 1'b1;  addr_rom[15212]='h00002138;  wr_data_rom[15212]='h00001322;
    rd_cycle[15213] = 1'b0;  wr_cycle[15213] = 1'b1;  addr_rom[15213]='h00001fc0;  wr_data_rom[15213]='h00001cdc;
    rd_cycle[15214] = 1'b1;  wr_cycle[15214] = 1'b0;  addr_rom[15214]='h0000022c;  wr_data_rom[15214]='h00000000;
    rd_cycle[15215] = 1'b1;  wr_cycle[15215] = 1'b0;  addr_rom[15215]='h00001660;  wr_data_rom[15215]='h00000000;
    rd_cycle[15216] = 1'b0;  wr_cycle[15216] = 1'b1;  addr_rom[15216]='h00002ff4;  wr_data_rom[15216]='h00003fe9;
    rd_cycle[15217] = 1'b0;  wr_cycle[15217] = 1'b1;  addr_rom[15217]='h00003b24;  wr_data_rom[15217]='h0000040a;
    rd_cycle[15218] = 1'b1;  wr_cycle[15218] = 1'b0;  addr_rom[15218]='h00001b3c;  wr_data_rom[15218]='h00000000;
    rd_cycle[15219] = 1'b0;  wr_cycle[15219] = 1'b1;  addr_rom[15219]='h0000285c;  wr_data_rom[15219]='h00003b86;
    rd_cycle[15220] = 1'b1;  wr_cycle[15220] = 1'b0;  addr_rom[15220]='h000004ec;  wr_data_rom[15220]='h00000000;
    rd_cycle[15221] = 1'b1;  wr_cycle[15221] = 1'b0;  addr_rom[15221]='h00002c68;  wr_data_rom[15221]='h00000000;
    rd_cycle[15222] = 1'b1;  wr_cycle[15222] = 1'b0;  addr_rom[15222]='h00001fb4;  wr_data_rom[15222]='h00000000;
    rd_cycle[15223] = 1'b1;  wr_cycle[15223] = 1'b0;  addr_rom[15223]='h00001e7c;  wr_data_rom[15223]='h00000000;
    rd_cycle[15224] = 1'b1;  wr_cycle[15224] = 1'b0;  addr_rom[15224]='h00002a80;  wr_data_rom[15224]='h00000000;
    rd_cycle[15225] = 1'b0;  wr_cycle[15225] = 1'b1;  addr_rom[15225]='h00001bc8;  wr_data_rom[15225]='h00003007;
    rd_cycle[15226] = 1'b1;  wr_cycle[15226] = 1'b0;  addr_rom[15226]='h00002da0;  wr_data_rom[15226]='h00000000;
    rd_cycle[15227] = 1'b0;  wr_cycle[15227] = 1'b1;  addr_rom[15227]='h00002510;  wr_data_rom[15227]='h00000686;
    rd_cycle[15228] = 1'b0;  wr_cycle[15228] = 1'b1;  addr_rom[15228]='h00002854;  wr_data_rom[15228]='h00003a8d;
    rd_cycle[15229] = 1'b1;  wr_cycle[15229] = 1'b0;  addr_rom[15229]='h00003bd0;  wr_data_rom[15229]='h00000000;
    rd_cycle[15230] = 1'b0;  wr_cycle[15230] = 1'b1;  addr_rom[15230]='h00001984;  wr_data_rom[15230]='h00002978;
    rd_cycle[15231] = 1'b0;  wr_cycle[15231] = 1'b1;  addr_rom[15231]='h00001c28;  wr_data_rom[15231]='h00002385;
    rd_cycle[15232] = 1'b0;  wr_cycle[15232] = 1'b1;  addr_rom[15232]='h00000328;  wr_data_rom[15232]='h00001dc4;
    rd_cycle[15233] = 1'b0;  wr_cycle[15233] = 1'b1;  addr_rom[15233]='h00001680;  wr_data_rom[15233]='h00001f89;
    rd_cycle[15234] = 1'b0;  wr_cycle[15234] = 1'b1;  addr_rom[15234]='h00001158;  wr_data_rom[15234]='h000010f5;
    rd_cycle[15235] = 1'b0;  wr_cycle[15235] = 1'b1;  addr_rom[15235]='h000022c4;  wr_data_rom[15235]='h000020ac;
    rd_cycle[15236] = 1'b1;  wr_cycle[15236] = 1'b0;  addr_rom[15236]='h00003004;  wr_data_rom[15236]='h00000000;
    rd_cycle[15237] = 1'b1;  wr_cycle[15237] = 1'b0;  addr_rom[15237]='h00003f44;  wr_data_rom[15237]='h00000000;
    rd_cycle[15238] = 1'b0;  wr_cycle[15238] = 1'b1;  addr_rom[15238]='h000024b0;  wr_data_rom[15238]='h000016e9;
    rd_cycle[15239] = 1'b0;  wr_cycle[15239] = 1'b1;  addr_rom[15239]='h00002df8;  wr_data_rom[15239]='h0000207b;
    rd_cycle[15240] = 1'b0;  wr_cycle[15240] = 1'b1;  addr_rom[15240]='h000012cc;  wr_data_rom[15240]='h0000131a;
    rd_cycle[15241] = 1'b0;  wr_cycle[15241] = 1'b1;  addr_rom[15241]='h00001ff0;  wr_data_rom[15241]='h0000011b;
    rd_cycle[15242] = 1'b1;  wr_cycle[15242] = 1'b0;  addr_rom[15242]='h000009a8;  wr_data_rom[15242]='h00000000;
    rd_cycle[15243] = 1'b0;  wr_cycle[15243] = 1'b1;  addr_rom[15243]='h00000e90;  wr_data_rom[15243]='h00002dec;
    rd_cycle[15244] = 1'b0;  wr_cycle[15244] = 1'b1;  addr_rom[15244]='h00003e88;  wr_data_rom[15244]='h00002353;
    rd_cycle[15245] = 1'b0;  wr_cycle[15245] = 1'b1;  addr_rom[15245]='h0000303c;  wr_data_rom[15245]='h00000ea0;
    rd_cycle[15246] = 1'b1;  wr_cycle[15246] = 1'b0;  addr_rom[15246]='h00001e60;  wr_data_rom[15246]='h00000000;
    rd_cycle[15247] = 1'b1;  wr_cycle[15247] = 1'b0;  addr_rom[15247]='h00003c4c;  wr_data_rom[15247]='h00000000;
    rd_cycle[15248] = 1'b1;  wr_cycle[15248] = 1'b0;  addr_rom[15248]='h00003254;  wr_data_rom[15248]='h00000000;
    rd_cycle[15249] = 1'b0;  wr_cycle[15249] = 1'b1;  addr_rom[15249]='h00003750;  wr_data_rom[15249]='h00000670;
    rd_cycle[15250] = 1'b0;  wr_cycle[15250] = 1'b1;  addr_rom[15250]='h00002464;  wr_data_rom[15250]='h00001a7c;
    rd_cycle[15251] = 1'b1;  wr_cycle[15251] = 1'b0;  addr_rom[15251]='h0000027c;  wr_data_rom[15251]='h00000000;
    rd_cycle[15252] = 1'b1;  wr_cycle[15252] = 1'b0;  addr_rom[15252]='h000019b4;  wr_data_rom[15252]='h00000000;
    rd_cycle[15253] = 1'b0;  wr_cycle[15253] = 1'b1;  addr_rom[15253]='h00001e54;  wr_data_rom[15253]='h00001dad;
    rd_cycle[15254] = 1'b0;  wr_cycle[15254] = 1'b1;  addr_rom[15254]='h00001fac;  wr_data_rom[15254]='h0000025d;
    rd_cycle[15255] = 1'b0;  wr_cycle[15255] = 1'b1;  addr_rom[15255]='h00000bb8;  wr_data_rom[15255]='h00001a93;
    rd_cycle[15256] = 1'b1;  wr_cycle[15256] = 1'b0;  addr_rom[15256]='h00002ff4;  wr_data_rom[15256]='h00000000;
    rd_cycle[15257] = 1'b1;  wr_cycle[15257] = 1'b0;  addr_rom[15257]='h0000001c;  wr_data_rom[15257]='h00000000;
    rd_cycle[15258] = 1'b0;  wr_cycle[15258] = 1'b1;  addr_rom[15258]='h00003650;  wr_data_rom[15258]='h000017b9;
    rd_cycle[15259] = 1'b0;  wr_cycle[15259] = 1'b1;  addr_rom[15259]='h0000007c;  wr_data_rom[15259]='h00000f0a;
    rd_cycle[15260] = 1'b1;  wr_cycle[15260] = 1'b0;  addr_rom[15260]='h00002eac;  wr_data_rom[15260]='h00000000;
    rd_cycle[15261] = 1'b0;  wr_cycle[15261] = 1'b1;  addr_rom[15261]='h00003378;  wr_data_rom[15261]='h00002a60;
    rd_cycle[15262] = 1'b1;  wr_cycle[15262] = 1'b0;  addr_rom[15262]='h0000273c;  wr_data_rom[15262]='h00000000;
    rd_cycle[15263] = 1'b0;  wr_cycle[15263] = 1'b1;  addr_rom[15263]='h00003960;  wr_data_rom[15263]='h00003c6f;
    rd_cycle[15264] = 1'b0;  wr_cycle[15264] = 1'b1;  addr_rom[15264]='h00001e80;  wr_data_rom[15264]='h000037d8;
    rd_cycle[15265] = 1'b0;  wr_cycle[15265] = 1'b1;  addr_rom[15265]='h0000001c;  wr_data_rom[15265]='h00000f46;
    rd_cycle[15266] = 1'b0;  wr_cycle[15266] = 1'b1;  addr_rom[15266]='h00000698;  wr_data_rom[15266]='h00000631;
    rd_cycle[15267] = 1'b0;  wr_cycle[15267] = 1'b1;  addr_rom[15267]='h000008dc;  wr_data_rom[15267]='h0000053f;
    rd_cycle[15268] = 1'b1;  wr_cycle[15268] = 1'b0;  addr_rom[15268]='h000015a0;  wr_data_rom[15268]='h00000000;
    rd_cycle[15269] = 1'b0;  wr_cycle[15269] = 1'b1;  addr_rom[15269]='h00000f94;  wr_data_rom[15269]='h00001ff0;
    rd_cycle[15270] = 1'b0;  wr_cycle[15270] = 1'b1;  addr_rom[15270]='h00000810;  wr_data_rom[15270]='h00003596;
    rd_cycle[15271] = 1'b0;  wr_cycle[15271] = 1'b1;  addr_rom[15271]='h000001a0;  wr_data_rom[15271]='h00001cc4;
    rd_cycle[15272] = 1'b1;  wr_cycle[15272] = 1'b0;  addr_rom[15272]='h00000894;  wr_data_rom[15272]='h00000000;
    rd_cycle[15273] = 1'b0;  wr_cycle[15273] = 1'b1;  addr_rom[15273]='h000002bc;  wr_data_rom[15273]='h00003b3c;
    rd_cycle[15274] = 1'b1;  wr_cycle[15274] = 1'b0;  addr_rom[15274]='h00002998;  wr_data_rom[15274]='h00000000;
    rd_cycle[15275] = 1'b0;  wr_cycle[15275] = 1'b1;  addr_rom[15275]='h0000100c;  wr_data_rom[15275]='h00000165;
    rd_cycle[15276] = 1'b1;  wr_cycle[15276] = 1'b0;  addr_rom[15276]='h000002f8;  wr_data_rom[15276]='h00000000;
    rd_cycle[15277] = 1'b1;  wr_cycle[15277] = 1'b0;  addr_rom[15277]='h0000307c;  wr_data_rom[15277]='h00000000;
    rd_cycle[15278] = 1'b0;  wr_cycle[15278] = 1'b1;  addr_rom[15278]='h00002314;  wr_data_rom[15278]='h00003440;
    rd_cycle[15279] = 1'b1;  wr_cycle[15279] = 1'b0;  addr_rom[15279]='h00000110;  wr_data_rom[15279]='h00000000;
    rd_cycle[15280] = 1'b1;  wr_cycle[15280] = 1'b0;  addr_rom[15280]='h000035f8;  wr_data_rom[15280]='h00000000;
    rd_cycle[15281] = 1'b1;  wr_cycle[15281] = 1'b0;  addr_rom[15281]='h00000364;  wr_data_rom[15281]='h00000000;
    rd_cycle[15282] = 1'b1;  wr_cycle[15282] = 1'b0;  addr_rom[15282]='h000030a8;  wr_data_rom[15282]='h00000000;
    rd_cycle[15283] = 1'b1;  wr_cycle[15283] = 1'b0;  addr_rom[15283]='h00001c1c;  wr_data_rom[15283]='h00000000;
    rd_cycle[15284] = 1'b1;  wr_cycle[15284] = 1'b0;  addr_rom[15284]='h000023e0;  wr_data_rom[15284]='h00000000;
    rd_cycle[15285] = 1'b1;  wr_cycle[15285] = 1'b0;  addr_rom[15285]='h00002c44;  wr_data_rom[15285]='h00000000;
    rd_cycle[15286] = 1'b0;  wr_cycle[15286] = 1'b1;  addr_rom[15286]='h000016cc;  wr_data_rom[15286]='h00001299;
    rd_cycle[15287] = 1'b1;  wr_cycle[15287] = 1'b0;  addr_rom[15287]='h000004a0;  wr_data_rom[15287]='h00000000;
    rd_cycle[15288] = 1'b0;  wr_cycle[15288] = 1'b1;  addr_rom[15288]='h0000044c;  wr_data_rom[15288]='h00001bc2;
    rd_cycle[15289] = 1'b0;  wr_cycle[15289] = 1'b1;  addr_rom[15289]='h000015d0;  wr_data_rom[15289]='h00003fa2;
    rd_cycle[15290] = 1'b1;  wr_cycle[15290] = 1'b0;  addr_rom[15290]='h00001da4;  wr_data_rom[15290]='h00000000;
    rd_cycle[15291] = 1'b1;  wr_cycle[15291] = 1'b0;  addr_rom[15291]='h00001b5c;  wr_data_rom[15291]='h00000000;
    rd_cycle[15292] = 1'b0;  wr_cycle[15292] = 1'b1;  addr_rom[15292]='h00000b24;  wr_data_rom[15292]='h00003781;
    rd_cycle[15293] = 1'b0;  wr_cycle[15293] = 1'b1;  addr_rom[15293]='h00001b08;  wr_data_rom[15293]='h000007e0;
    rd_cycle[15294] = 1'b0;  wr_cycle[15294] = 1'b1;  addr_rom[15294]='h00001da0;  wr_data_rom[15294]='h00000fc9;
    rd_cycle[15295] = 1'b1;  wr_cycle[15295] = 1'b0;  addr_rom[15295]='h000005c8;  wr_data_rom[15295]='h00000000;
    rd_cycle[15296] = 1'b0;  wr_cycle[15296] = 1'b1;  addr_rom[15296]='h00001a50;  wr_data_rom[15296]='h00001408;
    rd_cycle[15297] = 1'b0;  wr_cycle[15297] = 1'b1;  addr_rom[15297]='h0000122c;  wr_data_rom[15297]='h00003606;
    rd_cycle[15298] = 1'b0;  wr_cycle[15298] = 1'b1;  addr_rom[15298]='h00001870;  wr_data_rom[15298]='h000020a8;
    rd_cycle[15299] = 1'b1;  wr_cycle[15299] = 1'b0;  addr_rom[15299]='h00002510;  wr_data_rom[15299]='h00000000;
    rd_cycle[15300] = 1'b1;  wr_cycle[15300] = 1'b0;  addr_rom[15300]='h00002d50;  wr_data_rom[15300]='h00000000;
    rd_cycle[15301] = 1'b1;  wr_cycle[15301] = 1'b0;  addr_rom[15301]='h000014ec;  wr_data_rom[15301]='h00000000;
    rd_cycle[15302] = 1'b1;  wr_cycle[15302] = 1'b0;  addr_rom[15302]='h00001418;  wr_data_rom[15302]='h00000000;
    rd_cycle[15303] = 1'b0;  wr_cycle[15303] = 1'b1;  addr_rom[15303]='h00000254;  wr_data_rom[15303]='h00002e8e;
    rd_cycle[15304] = 1'b0;  wr_cycle[15304] = 1'b1;  addr_rom[15304]='h0000221c;  wr_data_rom[15304]='h00002878;
    rd_cycle[15305] = 1'b0;  wr_cycle[15305] = 1'b1;  addr_rom[15305]='h0000094c;  wr_data_rom[15305]='h00003bd1;
    rd_cycle[15306] = 1'b1;  wr_cycle[15306] = 1'b0;  addr_rom[15306]='h00003790;  wr_data_rom[15306]='h00000000;
    rd_cycle[15307] = 1'b0;  wr_cycle[15307] = 1'b1;  addr_rom[15307]='h00001540;  wr_data_rom[15307]='h00002227;
    rd_cycle[15308] = 1'b0;  wr_cycle[15308] = 1'b1;  addr_rom[15308]='h00001a40;  wr_data_rom[15308]='h00002bff;
    rd_cycle[15309] = 1'b0;  wr_cycle[15309] = 1'b1;  addr_rom[15309]='h00000b18;  wr_data_rom[15309]='h000010af;
    rd_cycle[15310] = 1'b0;  wr_cycle[15310] = 1'b1;  addr_rom[15310]='h00002f5c;  wr_data_rom[15310]='h00002a8d;
    rd_cycle[15311] = 1'b0;  wr_cycle[15311] = 1'b1;  addr_rom[15311]='h00003f70;  wr_data_rom[15311]='h000016cf;
    rd_cycle[15312] = 1'b1;  wr_cycle[15312] = 1'b0;  addr_rom[15312]='h00000978;  wr_data_rom[15312]='h00000000;
    rd_cycle[15313] = 1'b1;  wr_cycle[15313] = 1'b0;  addr_rom[15313]='h00002a0c;  wr_data_rom[15313]='h00000000;
    rd_cycle[15314] = 1'b1;  wr_cycle[15314] = 1'b0;  addr_rom[15314]='h00003278;  wr_data_rom[15314]='h00000000;
    rd_cycle[15315] = 1'b1;  wr_cycle[15315] = 1'b0;  addr_rom[15315]='h000007a0;  wr_data_rom[15315]='h00000000;
    rd_cycle[15316] = 1'b1;  wr_cycle[15316] = 1'b0;  addr_rom[15316]='h00000db8;  wr_data_rom[15316]='h00000000;
    rd_cycle[15317] = 1'b1;  wr_cycle[15317] = 1'b0;  addr_rom[15317]='h00001950;  wr_data_rom[15317]='h00000000;
    rd_cycle[15318] = 1'b1;  wr_cycle[15318] = 1'b0;  addr_rom[15318]='h00000524;  wr_data_rom[15318]='h00000000;
    rd_cycle[15319] = 1'b1;  wr_cycle[15319] = 1'b0;  addr_rom[15319]='h000025e0;  wr_data_rom[15319]='h00000000;
    rd_cycle[15320] = 1'b1;  wr_cycle[15320] = 1'b0;  addr_rom[15320]='h000007f4;  wr_data_rom[15320]='h00000000;
    rd_cycle[15321] = 1'b1;  wr_cycle[15321] = 1'b0;  addr_rom[15321]='h000016d4;  wr_data_rom[15321]='h00000000;
    rd_cycle[15322] = 1'b1;  wr_cycle[15322] = 1'b0;  addr_rom[15322]='h00001018;  wr_data_rom[15322]='h00000000;
    rd_cycle[15323] = 1'b1;  wr_cycle[15323] = 1'b0;  addr_rom[15323]='h00002780;  wr_data_rom[15323]='h00000000;
    rd_cycle[15324] = 1'b1;  wr_cycle[15324] = 1'b0;  addr_rom[15324]='h00003280;  wr_data_rom[15324]='h00000000;
    rd_cycle[15325] = 1'b1;  wr_cycle[15325] = 1'b0;  addr_rom[15325]='h00003498;  wr_data_rom[15325]='h00000000;
    rd_cycle[15326] = 1'b1;  wr_cycle[15326] = 1'b0;  addr_rom[15326]='h0000059c;  wr_data_rom[15326]='h00000000;
    rd_cycle[15327] = 1'b1;  wr_cycle[15327] = 1'b0;  addr_rom[15327]='h00002194;  wr_data_rom[15327]='h00000000;
    rd_cycle[15328] = 1'b1;  wr_cycle[15328] = 1'b0;  addr_rom[15328]='h000018fc;  wr_data_rom[15328]='h00000000;
    rd_cycle[15329] = 1'b0;  wr_cycle[15329] = 1'b1;  addr_rom[15329]='h00002a28;  wr_data_rom[15329]='h00001c57;
    rd_cycle[15330] = 1'b1;  wr_cycle[15330] = 1'b0;  addr_rom[15330]='h00002db4;  wr_data_rom[15330]='h00000000;
    rd_cycle[15331] = 1'b1;  wr_cycle[15331] = 1'b0;  addr_rom[15331]='h00003b40;  wr_data_rom[15331]='h00000000;
    rd_cycle[15332] = 1'b0;  wr_cycle[15332] = 1'b1;  addr_rom[15332]='h00003a38;  wr_data_rom[15332]='h0000260d;
    rd_cycle[15333] = 1'b0;  wr_cycle[15333] = 1'b1;  addr_rom[15333]='h00001060;  wr_data_rom[15333]='h00003491;
    rd_cycle[15334] = 1'b0;  wr_cycle[15334] = 1'b1;  addr_rom[15334]='h000016a0;  wr_data_rom[15334]='h00003ff7;
    rd_cycle[15335] = 1'b1;  wr_cycle[15335] = 1'b0;  addr_rom[15335]='h00003180;  wr_data_rom[15335]='h00000000;
    rd_cycle[15336] = 1'b0;  wr_cycle[15336] = 1'b1;  addr_rom[15336]='h0000082c;  wr_data_rom[15336]='h00001d2d;
    rd_cycle[15337] = 1'b1;  wr_cycle[15337] = 1'b0;  addr_rom[15337]='h00001d7c;  wr_data_rom[15337]='h00000000;
    rd_cycle[15338] = 1'b1;  wr_cycle[15338] = 1'b0;  addr_rom[15338]='h000000fc;  wr_data_rom[15338]='h00000000;
    rd_cycle[15339] = 1'b0;  wr_cycle[15339] = 1'b1;  addr_rom[15339]='h000018c8;  wr_data_rom[15339]='h000012e6;
    rd_cycle[15340] = 1'b0;  wr_cycle[15340] = 1'b1;  addr_rom[15340]='h00002a4c;  wr_data_rom[15340]='h000023ff;
    rd_cycle[15341] = 1'b0;  wr_cycle[15341] = 1'b1;  addr_rom[15341]='h0000292c;  wr_data_rom[15341]='h00003ab7;
    rd_cycle[15342] = 1'b1;  wr_cycle[15342] = 1'b0;  addr_rom[15342]='h00002550;  wr_data_rom[15342]='h00000000;
    rd_cycle[15343] = 1'b1;  wr_cycle[15343] = 1'b0;  addr_rom[15343]='h00000bf0;  wr_data_rom[15343]='h00000000;
    rd_cycle[15344] = 1'b0;  wr_cycle[15344] = 1'b1;  addr_rom[15344]='h00003b04;  wr_data_rom[15344]='h000000c1;
    rd_cycle[15345] = 1'b1;  wr_cycle[15345] = 1'b0;  addr_rom[15345]='h000019f4;  wr_data_rom[15345]='h00000000;
    rd_cycle[15346] = 1'b1;  wr_cycle[15346] = 1'b0;  addr_rom[15346]='h00001b34;  wr_data_rom[15346]='h00000000;
    rd_cycle[15347] = 1'b0;  wr_cycle[15347] = 1'b1;  addr_rom[15347]='h0000089c;  wr_data_rom[15347]='h00000f09;
    rd_cycle[15348] = 1'b0;  wr_cycle[15348] = 1'b1;  addr_rom[15348]='h00002fdc;  wr_data_rom[15348]='h00001b88;
    rd_cycle[15349] = 1'b0;  wr_cycle[15349] = 1'b1;  addr_rom[15349]='h00000114;  wr_data_rom[15349]='h000029c8;
    rd_cycle[15350] = 1'b1;  wr_cycle[15350] = 1'b0;  addr_rom[15350]='h00001034;  wr_data_rom[15350]='h00000000;
    rd_cycle[15351] = 1'b1;  wr_cycle[15351] = 1'b0;  addr_rom[15351]='h00002d38;  wr_data_rom[15351]='h00000000;
    rd_cycle[15352] = 1'b0;  wr_cycle[15352] = 1'b1;  addr_rom[15352]='h000034e8;  wr_data_rom[15352]='h00001b57;
    rd_cycle[15353] = 1'b0;  wr_cycle[15353] = 1'b1;  addr_rom[15353]='h00002180;  wr_data_rom[15353]='h00002f44;
    rd_cycle[15354] = 1'b0;  wr_cycle[15354] = 1'b1;  addr_rom[15354]='h00003ff8;  wr_data_rom[15354]='h00001a1f;
    rd_cycle[15355] = 1'b0;  wr_cycle[15355] = 1'b1;  addr_rom[15355]='h00000870;  wr_data_rom[15355]='h00002063;
    rd_cycle[15356] = 1'b0;  wr_cycle[15356] = 1'b1;  addr_rom[15356]='h000000d0;  wr_data_rom[15356]='h00000c13;
    rd_cycle[15357] = 1'b0;  wr_cycle[15357] = 1'b1;  addr_rom[15357]='h000028fc;  wr_data_rom[15357]='h00002c8e;
    rd_cycle[15358] = 1'b0;  wr_cycle[15358] = 1'b1;  addr_rom[15358]='h00002f48;  wr_data_rom[15358]='h000006f9;
    rd_cycle[15359] = 1'b1;  wr_cycle[15359] = 1'b0;  addr_rom[15359]='h00000654;  wr_data_rom[15359]='h00000000;
    rd_cycle[15360] = 1'b1;  wr_cycle[15360] = 1'b0;  addr_rom[15360]='h000012dc;  wr_data_rom[15360]='h00000000;
    rd_cycle[15361] = 1'b0;  wr_cycle[15361] = 1'b1;  addr_rom[15361]='h00002280;  wr_data_rom[15361]='h000019a8;
    rd_cycle[15362] = 1'b1;  wr_cycle[15362] = 1'b0;  addr_rom[15362]='h00002854;  wr_data_rom[15362]='h00000000;
    rd_cycle[15363] = 1'b0;  wr_cycle[15363] = 1'b1;  addr_rom[15363]='h000016e0;  wr_data_rom[15363]='h000008b8;
    rd_cycle[15364] = 1'b0;  wr_cycle[15364] = 1'b1;  addr_rom[15364]='h00000144;  wr_data_rom[15364]='h0000038b;
    rd_cycle[15365] = 1'b1;  wr_cycle[15365] = 1'b0;  addr_rom[15365]='h000038a8;  wr_data_rom[15365]='h00000000;
    rd_cycle[15366] = 1'b1;  wr_cycle[15366] = 1'b0;  addr_rom[15366]='h00001eb4;  wr_data_rom[15366]='h00000000;
    rd_cycle[15367] = 1'b1;  wr_cycle[15367] = 1'b0;  addr_rom[15367]='h000018d0;  wr_data_rom[15367]='h00000000;
    rd_cycle[15368] = 1'b1;  wr_cycle[15368] = 1'b0;  addr_rom[15368]='h00003e44;  wr_data_rom[15368]='h00000000;
    rd_cycle[15369] = 1'b1;  wr_cycle[15369] = 1'b0;  addr_rom[15369]='h00001608;  wr_data_rom[15369]='h00000000;
    rd_cycle[15370] = 1'b0;  wr_cycle[15370] = 1'b1;  addr_rom[15370]='h0000204c;  wr_data_rom[15370]='h000031f8;
    rd_cycle[15371] = 1'b0;  wr_cycle[15371] = 1'b1;  addr_rom[15371]='h00003f6c;  wr_data_rom[15371]='h00003965;
    rd_cycle[15372] = 1'b1;  wr_cycle[15372] = 1'b0;  addr_rom[15372]='h00002b98;  wr_data_rom[15372]='h00000000;
    rd_cycle[15373] = 1'b0;  wr_cycle[15373] = 1'b1;  addr_rom[15373]='h00003214;  wr_data_rom[15373]='h00003a00;
    rd_cycle[15374] = 1'b1;  wr_cycle[15374] = 1'b0;  addr_rom[15374]='h00002d58;  wr_data_rom[15374]='h00000000;
    rd_cycle[15375] = 1'b1;  wr_cycle[15375] = 1'b0;  addr_rom[15375]='h00003260;  wr_data_rom[15375]='h00000000;
    rd_cycle[15376] = 1'b1;  wr_cycle[15376] = 1'b0;  addr_rom[15376]='h00000958;  wr_data_rom[15376]='h00000000;
    rd_cycle[15377] = 1'b0;  wr_cycle[15377] = 1'b1;  addr_rom[15377]='h00002a00;  wr_data_rom[15377]='h00000c09;
    rd_cycle[15378] = 1'b1;  wr_cycle[15378] = 1'b0;  addr_rom[15378]='h00001990;  wr_data_rom[15378]='h00000000;
    rd_cycle[15379] = 1'b1;  wr_cycle[15379] = 1'b0;  addr_rom[15379]='h00000cbc;  wr_data_rom[15379]='h00000000;
    rd_cycle[15380] = 1'b1;  wr_cycle[15380] = 1'b0;  addr_rom[15380]='h00000c94;  wr_data_rom[15380]='h00000000;
    rd_cycle[15381] = 1'b1;  wr_cycle[15381] = 1'b0;  addr_rom[15381]='h000027ec;  wr_data_rom[15381]='h00000000;
    rd_cycle[15382] = 1'b1;  wr_cycle[15382] = 1'b0;  addr_rom[15382]='h00001c70;  wr_data_rom[15382]='h00000000;
    rd_cycle[15383] = 1'b1;  wr_cycle[15383] = 1'b0;  addr_rom[15383]='h00003604;  wr_data_rom[15383]='h00000000;
    rd_cycle[15384] = 1'b1;  wr_cycle[15384] = 1'b0;  addr_rom[15384]='h00000044;  wr_data_rom[15384]='h00000000;
    rd_cycle[15385] = 1'b0;  wr_cycle[15385] = 1'b1;  addr_rom[15385]='h00000b00;  wr_data_rom[15385]='h00002673;
    rd_cycle[15386] = 1'b0;  wr_cycle[15386] = 1'b1;  addr_rom[15386]='h00003ec4;  wr_data_rom[15386]='h000011ef;
    rd_cycle[15387] = 1'b0;  wr_cycle[15387] = 1'b1;  addr_rom[15387]='h00003e7c;  wr_data_rom[15387]='h00003d09;
    rd_cycle[15388] = 1'b1;  wr_cycle[15388] = 1'b0;  addr_rom[15388]='h00002494;  wr_data_rom[15388]='h00000000;
    rd_cycle[15389] = 1'b1;  wr_cycle[15389] = 1'b0;  addr_rom[15389]='h00002f38;  wr_data_rom[15389]='h00000000;
    rd_cycle[15390] = 1'b0;  wr_cycle[15390] = 1'b1;  addr_rom[15390]='h00000bc4;  wr_data_rom[15390]='h0000179c;
    rd_cycle[15391] = 1'b0;  wr_cycle[15391] = 1'b1;  addr_rom[15391]='h0000358c;  wr_data_rom[15391]='h00000d1a;
    rd_cycle[15392] = 1'b0;  wr_cycle[15392] = 1'b1;  addr_rom[15392]='h0000289c;  wr_data_rom[15392]='h000036f9;
    rd_cycle[15393] = 1'b0;  wr_cycle[15393] = 1'b1;  addr_rom[15393]='h000002fc;  wr_data_rom[15393]='h000037ad;
    rd_cycle[15394] = 1'b0;  wr_cycle[15394] = 1'b1;  addr_rom[15394]='h000010c0;  wr_data_rom[15394]='h0000166a;
    rd_cycle[15395] = 1'b0;  wr_cycle[15395] = 1'b1;  addr_rom[15395]='h00000208;  wr_data_rom[15395]='h00002281;
    rd_cycle[15396] = 1'b0;  wr_cycle[15396] = 1'b1;  addr_rom[15396]='h00002bac;  wr_data_rom[15396]='h000032d4;
    rd_cycle[15397] = 1'b0;  wr_cycle[15397] = 1'b1;  addr_rom[15397]='h00000160;  wr_data_rom[15397]='h00001406;
    rd_cycle[15398] = 1'b0;  wr_cycle[15398] = 1'b1;  addr_rom[15398]='h000029ac;  wr_data_rom[15398]='h00003806;
    rd_cycle[15399] = 1'b1;  wr_cycle[15399] = 1'b0;  addr_rom[15399]='h00000d74;  wr_data_rom[15399]='h00000000;
    rd_cycle[15400] = 1'b1;  wr_cycle[15400] = 1'b0;  addr_rom[15400]='h000034f0;  wr_data_rom[15400]='h00000000;
    rd_cycle[15401] = 1'b1;  wr_cycle[15401] = 1'b0;  addr_rom[15401]='h000038c4;  wr_data_rom[15401]='h00000000;
    rd_cycle[15402] = 1'b0;  wr_cycle[15402] = 1'b1;  addr_rom[15402]='h0000248c;  wr_data_rom[15402]='h00000447;
    rd_cycle[15403] = 1'b0;  wr_cycle[15403] = 1'b1;  addr_rom[15403]='h00000118;  wr_data_rom[15403]='h00002c53;
    rd_cycle[15404] = 1'b1;  wr_cycle[15404] = 1'b0;  addr_rom[15404]='h00002a4c;  wr_data_rom[15404]='h00000000;
    rd_cycle[15405] = 1'b1;  wr_cycle[15405] = 1'b0;  addr_rom[15405]='h00001e1c;  wr_data_rom[15405]='h00000000;
    rd_cycle[15406] = 1'b1;  wr_cycle[15406] = 1'b0;  addr_rom[15406]='h00002c70;  wr_data_rom[15406]='h00000000;
    rd_cycle[15407] = 1'b0;  wr_cycle[15407] = 1'b1;  addr_rom[15407]='h00002780;  wr_data_rom[15407]='h0000186c;
    rd_cycle[15408] = 1'b0;  wr_cycle[15408] = 1'b1;  addr_rom[15408]='h0000003c;  wr_data_rom[15408]='h00002d7d;
    rd_cycle[15409] = 1'b0;  wr_cycle[15409] = 1'b1;  addr_rom[15409]='h00002bf4;  wr_data_rom[15409]='h00001a90;
    rd_cycle[15410] = 1'b1;  wr_cycle[15410] = 1'b0;  addr_rom[15410]='h000019e0;  wr_data_rom[15410]='h00000000;
    rd_cycle[15411] = 1'b1;  wr_cycle[15411] = 1'b0;  addr_rom[15411]='h000020e8;  wr_data_rom[15411]='h00000000;
    rd_cycle[15412] = 1'b0;  wr_cycle[15412] = 1'b1;  addr_rom[15412]='h00001528;  wr_data_rom[15412]='h000039ec;
    rd_cycle[15413] = 1'b1;  wr_cycle[15413] = 1'b0;  addr_rom[15413]='h00003a5c;  wr_data_rom[15413]='h00000000;
    rd_cycle[15414] = 1'b0;  wr_cycle[15414] = 1'b1;  addr_rom[15414]='h000028b0;  wr_data_rom[15414]='h00001f70;
    rd_cycle[15415] = 1'b1;  wr_cycle[15415] = 1'b0;  addr_rom[15415]='h00003138;  wr_data_rom[15415]='h00000000;
    rd_cycle[15416] = 1'b0;  wr_cycle[15416] = 1'b1;  addr_rom[15416]='h00000054;  wr_data_rom[15416]='h00001bee;
    rd_cycle[15417] = 1'b1;  wr_cycle[15417] = 1'b0;  addr_rom[15417]='h00000784;  wr_data_rom[15417]='h00000000;
    rd_cycle[15418] = 1'b0;  wr_cycle[15418] = 1'b1;  addr_rom[15418]='h000020a8;  wr_data_rom[15418]='h0000174e;
    rd_cycle[15419] = 1'b1;  wr_cycle[15419] = 1'b0;  addr_rom[15419]='h0000199c;  wr_data_rom[15419]='h00000000;
    rd_cycle[15420] = 1'b0;  wr_cycle[15420] = 1'b1;  addr_rom[15420]='h00002784;  wr_data_rom[15420]='h00002017;
    rd_cycle[15421] = 1'b0;  wr_cycle[15421] = 1'b1;  addr_rom[15421]='h00001db4;  wr_data_rom[15421]='h00001f0c;
    rd_cycle[15422] = 1'b0;  wr_cycle[15422] = 1'b1;  addr_rom[15422]='h00000a80;  wr_data_rom[15422]='h00002d1b;
    rd_cycle[15423] = 1'b1;  wr_cycle[15423] = 1'b0;  addr_rom[15423]='h00002eac;  wr_data_rom[15423]='h00000000;
    rd_cycle[15424] = 1'b0;  wr_cycle[15424] = 1'b1;  addr_rom[15424]='h000033d4;  wr_data_rom[15424]='h000003d9;
    rd_cycle[15425] = 1'b1;  wr_cycle[15425] = 1'b0;  addr_rom[15425]='h00002d84;  wr_data_rom[15425]='h00000000;
    rd_cycle[15426] = 1'b0;  wr_cycle[15426] = 1'b1;  addr_rom[15426]='h000022a4;  wr_data_rom[15426]='h0000221d;
    rd_cycle[15427] = 1'b1;  wr_cycle[15427] = 1'b0;  addr_rom[15427]='h0000376c;  wr_data_rom[15427]='h00000000;
    rd_cycle[15428] = 1'b1;  wr_cycle[15428] = 1'b0;  addr_rom[15428]='h0000214c;  wr_data_rom[15428]='h00000000;
    rd_cycle[15429] = 1'b0;  wr_cycle[15429] = 1'b1;  addr_rom[15429]='h000020a8;  wr_data_rom[15429]='h00001254;
    rd_cycle[15430] = 1'b1;  wr_cycle[15430] = 1'b0;  addr_rom[15430]='h00003fbc;  wr_data_rom[15430]='h00000000;
    rd_cycle[15431] = 1'b1;  wr_cycle[15431] = 1'b0;  addr_rom[15431]='h00000ae8;  wr_data_rom[15431]='h00000000;
    rd_cycle[15432] = 1'b0;  wr_cycle[15432] = 1'b1;  addr_rom[15432]='h000007e4;  wr_data_rom[15432]='h00001100;
    rd_cycle[15433] = 1'b1;  wr_cycle[15433] = 1'b0;  addr_rom[15433]='h000003fc;  wr_data_rom[15433]='h00000000;
    rd_cycle[15434] = 1'b1;  wr_cycle[15434] = 1'b0;  addr_rom[15434]='h00001504;  wr_data_rom[15434]='h00000000;
    rd_cycle[15435] = 1'b0;  wr_cycle[15435] = 1'b1;  addr_rom[15435]='h00001d3c;  wr_data_rom[15435]='h00003814;
    rd_cycle[15436] = 1'b0;  wr_cycle[15436] = 1'b1;  addr_rom[15436]='h0000269c;  wr_data_rom[15436]='h000012d5;
    rd_cycle[15437] = 1'b1;  wr_cycle[15437] = 1'b0;  addr_rom[15437]='h000032e4;  wr_data_rom[15437]='h00000000;
    rd_cycle[15438] = 1'b0;  wr_cycle[15438] = 1'b1;  addr_rom[15438]='h0000015c;  wr_data_rom[15438]='h00002026;
    rd_cycle[15439] = 1'b1;  wr_cycle[15439] = 1'b0;  addr_rom[15439]='h00003538;  wr_data_rom[15439]='h00000000;
    rd_cycle[15440] = 1'b1;  wr_cycle[15440] = 1'b0;  addr_rom[15440]='h00001110;  wr_data_rom[15440]='h00000000;
    rd_cycle[15441] = 1'b1;  wr_cycle[15441] = 1'b0;  addr_rom[15441]='h00003f3c;  wr_data_rom[15441]='h00000000;
    rd_cycle[15442] = 1'b1;  wr_cycle[15442] = 1'b0;  addr_rom[15442]='h0000020c;  wr_data_rom[15442]='h00000000;
    rd_cycle[15443] = 1'b1;  wr_cycle[15443] = 1'b0;  addr_rom[15443]='h000027c0;  wr_data_rom[15443]='h00000000;
    rd_cycle[15444] = 1'b1;  wr_cycle[15444] = 1'b0;  addr_rom[15444]='h00000c08;  wr_data_rom[15444]='h00000000;
    rd_cycle[15445] = 1'b0;  wr_cycle[15445] = 1'b1;  addr_rom[15445]='h000029b4;  wr_data_rom[15445]='h00001b7c;
    rd_cycle[15446] = 1'b0;  wr_cycle[15446] = 1'b1;  addr_rom[15446]='h00000fd4;  wr_data_rom[15446]='h00003f05;
    rd_cycle[15447] = 1'b1;  wr_cycle[15447] = 1'b0;  addr_rom[15447]='h000035b4;  wr_data_rom[15447]='h00000000;
    rd_cycle[15448] = 1'b0;  wr_cycle[15448] = 1'b1;  addr_rom[15448]='h00003ffc;  wr_data_rom[15448]='h000033ed;
    rd_cycle[15449] = 1'b0;  wr_cycle[15449] = 1'b1;  addr_rom[15449]='h00003130;  wr_data_rom[15449]='h00000a83;
    rd_cycle[15450] = 1'b0;  wr_cycle[15450] = 1'b1;  addr_rom[15450]='h00002d7c;  wr_data_rom[15450]='h00002f3c;
    rd_cycle[15451] = 1'b0;  wr_cycle[15451] = 1'b1;  addr_rom[15451]='h0000254c;  wr_data_rom[15451]='h000010c7;
    rd_cycle[15452] = 1'b1;  wr_cycle[15452] = 1'b0;  addr_rom[15452]='h00002b2c;  wr_data_rom[15452]='h00000000;
    rd_cycle[15453] = 1'b1;  wr_cycle[15453] = 1'b0;  addr_rom[15453]='h00001708;  wr_data_rom[15453]='h00000000;
    rd_cycle[15454] = 1'b0;  wr_cycle[15454] = 1'b1;  addr_rom[15454]='h00002a14;  wr_data_rom[15454]='h000002c9;
    rd_cycle[15455] = 1'b1;  wr_cycle[15455] = 1'b0;  addr_rom[15455]='h000000a8;  wr_data_rom[15455]='h00000000;
    rd_cycle[15456] = 1'b1;  wr_cycle[15456] = 1'b0;  addr_rom[15456]='h00002b2c;  wr_data_rom[15456]='h00000000;
    rd_cycle[15457] = 1'b0;  wr_cycle[15457] = 1'b1;  addr_rom[15457]='h00002c60;  wr_data_rom[15457]='h000011b6;
    rd_cycle[15458] = 1'b0;  wr_cycle[15458] = 1'b1;  addr_rom[15458]='h00000e48;  wr_data_rom[15458]='h000034d0;
    rd_cycle[15459] = 1'b1;  wr_cycle[15459] = 1'b0;  addr_rom[15459]='h000022e4;  wr_data_rom[15459]='h00000000;
    rd_cycle[15460] = 1'b1;  wr_cycle[15460] = 1'b0;  addr_rom[15460]='h00003b4c;  wr_data_rom[15460]='h00000000;
    rd_cycle[15461] = 1'b0;  wr_cycle[15461] = 1'b1;  addr_rom[15461]='h000001d8;  wr_data_rom[15461]='h00001dcc;
    rd_cycle[15462] = 1'b1;  wr_cycle[15462] = 1'b0;  addr_rom[15462]='h00002b04;  wr_data_rom[15462]='h00000000;
    rd_cycle[15463] = 1'b1;  wr_cycle[15463] = 1'b0;  addr_rom[15463]='h00001c98;  wr_data_rom[15463]='h00000000;
    rd_cycle[15464] = 1'b0;  wr_cycle[15464] = 1'b1;  addr_rom[15464]='h00000124;  wr_data_rom[15464]='h00002e71;
    rd_cycle[15465] = 1'b0;  wr_cycle[15465] = 1'b1;  addr_rom[15465]='h00001820;  wr_data_rom[15465]='h00003d0c;
    rd_cycle[15466] = 1'b0;  wr_cycle[15466] = 1'b1;  addr_rom[15466]='h00001720;  wr_data_rom[15466]='h00001a53;
    rd_cycle[15467] = 1'b1;  wr_cycle[15467] = 1'b0;  addr_rom[15467]='h00002664;  wr_data_rom[15467]='h00000000;
    rd_cycle[15468] = 1'b1;  wr_cycle[15468] = 1'b0;  addr_rom[15468]='h000010a0;  wr_data_rom[15468]='h00000000;
    rd_cycle[15469] = 1'b0;  wr_cycle[15469] = 1'b1;  addr_rom[15469]='h000025ec;  wr_data_rom[15469]='h00001888;
    rd_cycle[15470] = 1'b1;  wr_cycle[15470] = 1'b0;  addr_rom[15470]='h00000700;  wr_data_rom[15470]='h00000000;
    rd_cycle[15471] = 1'b0;  wr_cycle[15471] = 1'b1;  addr_rom[15471]='h0000375c;  wr_data_rom[15471]='h00000372;
    rd_cycle[15472] = 1'b0;  wr_cycle[15472] = 1'b1;  addr_rom[15472]='h00003dbc;  wr_data_rom[15472]='h00003bf1;
    rd_cycle[15473] = 1'b1;  wr_cycle[15473] = 1'b0;  addr_rom[15473]='h00000b20;  wr_data_rom[15473]='h00000000;
    rd_cycle[15474] = 1'b1;  wr_cycle[15474] = 1'b0;  addr_rom[15474]='h000035e4;  wr_data_rom[15474]='h00000000;
    rd_cycle[15475] = 1'b0;  wr_cycle[15475] = 1'b1;  addr_rom[15475]='h00003374;  wr_data_rom[15475]='h0000256e;
    rd_cycle[15476] = 1'b1;  wr_cycle[15476] = 1'b0;  addr_rom[15476]='h00003f10;  wr_data_rom[15476]='h00000000;
    rd_cycle[15477] = 1'b0;  wr_cycle[15477] = 1'b1;  addr_rom[15477]='h00002e0c;  wr_data_rom[15477]='h00001710;
    rd_cycle[15478] = 1'b0;  wr_cycle[15478] = 1'b1;  addr_rom[15478]='h000034b8;  wr_data_rom[15478]='h00003323;
    rd_cycle[15479] = 1'b1;  wr_cycle[15479] = 1'b0;  addr_rom[15479]='h00001f40;  wr_data_rom[15479]='h00000000;
    rd_cycle[15480] = 1'b1;  wr_cycle[15480] = 1'b0;  addr_rom[15480]='h00003188;  wr_data_rom[15480]='h00000000;
    rd_cycle[15481] = 1'b1;  wr_cycle[15481] = 1'b0;  addr_rom[15481]='h00003408;  wr_data_rom[15481]='h00000000;
    rd_cycle[15482] = 1'b0;  wr_cycle[15482] = 1'b1;  addr_rom[15482]='h00002568;  wr_data_rom[15482]='h000004b5;
    rd_cycle[15483] = 1'b1;  wr_cycle[15483] = 1'b0;  addr_rom[15483]='h00003bf0;  wr_data_rom[15483]='h00000000;
    rd_cycle[15484] = 1'b0;  wr_cycle[15484] = 1'b1;  addr_rom[15484]='h000007bc;  wr_data_rom[15484]='h00003503;
    rd_cycle[15485] = 1'b0;  wr_cycle[15485] = 1'b1;  addr_rom[15485]='h00000c40;  wr_data_rom[15485]='h00003aa6;
    rd_cycle[15486] = 1'b1;  wr_cycle[15486] = 1'b0;  addr_rom[15486]='h00000f78;  wr_data_rom[15486]='h00000000;
    rd_cycle[15487] = 1'b1;  wr_cycle[15487] = 1'b0;  addr_rom[15487]='h00000898;  wr_data_rom[15487]='h00000000;
    rd_cycle[15488] = 1'b0;  wr_cycle[15488] = 1'b1;  addr_rom[15488]='h000001d0;  wr_data_rom[15488]='h00000cc4;
    rd_cycle[15489] = 1'b0;  wr_cycle[15489] = 1'b1;  addr_rom[15489]='h00002d0c;  wr_data_rom[15489]='h000020e8;
    rd_cycle[15490] = 1'b0;  wr_cycle[15490] = 1'b1;  addr_rom[15490]='h000011b4;  wr_data_rom[15490]='h0000178b;
    rd_cycle[15491] = 1'b0;  wr_cycle[15491] = 1'b1;  addr_rom[15491]='h00003a94;  wr_data_rom[15491]='h0000261a;
    rd_cycle[15492] = 1'b0;  wr_cycle[15492] = 1'b1;  addr_rom[15492]='h00000ca0;  wr_data_rom[15492]='h00003833;
    rd_cycle[15493] = 1'b1;  wr_cycle[15493] = 1'b0;  addr_rom[15493]='h000017dc;  wr_data_rom[15493]='h00000000;
    rd_cycle[15494] = 1'b1;  wr_cycle[15494] = 1'b0;  addr_rom[15494]='h00003040;  wr_data_rom[15494]='h00000000;
    rd_cycle[15495] = 1'b0;  wr_cycle[15495] = 1'b1;  addr_rom[15495]='h00000dec;  wr_data_rom[15495]='h000006d2;
    rd_cycle[15496] = 1'b1;  wr_cycle[15496] = 1'b0;  addr_rom[15496]='h00003d84;  wr_data_rom[15496]='h00000000;
    rd_cycle[15497] = 1'b0;  wr_cycle[15497] = 1'b1;  addr_rom[15497]='h00000308;  wr_data_rom[15497]='h000001e5;
    rd_cycle[15498] = 1'b1;  wr_cycle[15498] = 1'b0;  addr_rom[15498]='h00001cf0;  wr_data_rom[15498]='h00000000;
    rd_cycle[15499] = 1'b0;  wr_cycle[15499] = 1'b1;  addr_rom[15499]='h00002c24;  wr_data_rom[15499]='h00001351;
    rd_cycle[15500] = 1'b1;  wr_cycle[15500] = 1'b0;  addr_rom[15500]='h00001174;  wr_data_rom[15500]='h00000000;
    rd_cycle[15501] = 1'b1;  wr_cycle[15501] = 1'b0;  addr_rom[15501]='h00003610;  wr_data_rom[15501]='h00000000;
    rd_cycle[15502] = 1'b1;  wr_cycle[15502] = 1'b0;  addr_rom[15502]='h0000245c;  wr_data_rom[15502]='h00000000;
    rd_cycle[15503] = 1'b0;  wr_cycle[15503] = 1'b1;  addr_rom[15503]='h00000d18;  wr_data_rom[15503]='h00001d8a;
    rd_cycle[15504] = 1'b0;  wr_cycle[15504] = 1'b1;  addr_rom[15504]='h00000ac0;  wr_data_rom[15504]='h00000367;
    rd_cycle[15505] = 1'b0;  wr_cycle[15505] = 1'b1;  addr_rom[15505]='h000000cc;  wr_data_rom[15505]='h00001a35;
    rd_cycle[15506] = 1'b0;  wr_cycle[15506] = 1'b1;  addr_rom[15506]='h00003b68;  wr_data_rom[15506]='h0000113d;
    rd_cycle[15507] = 1'b0;  wr_cycle[15507] = 1'b1;  addr_rom[15507]='h000019a4;  wr_data_rom[15507]='h00003406;
    rd_cycle[15508] = 1'b0;  wr_cycle[15508] = 1'b1;  addr_rom[15508]='h00001e68;  wr_data_rom[15508]='h00003075;
    rd_cycle[15509] = 1'b0;  wr_cycle[15509] = 1'b1;  addr_rom[15509]='h000023d8;  wr_data_rom[15509]='h00001fa5;
    rd_cycle[15510] = 1'b0;  wr_cycle[15510] = 1'b1;  addr_rom[15510]='h0000143c;  wr_data_rom[15510]='h00000b54;
    rd_cycle[15511] = 1'b1;  wr_cycle[15511] = 1'b0;  addr_rom[15511]='h0000276c;  wr_data_rom[15511]='h00000000;
    rd_cycle[15512] = 1'b0;  wr_cycle[15512] = 1'b1;  addr_rom[15512]='h000032d0;  wr_data_rom[15512]='h00002a1f;
    rd_cycle[15513] = 1'b1;  wr_cycle[15513] = 1'b0;  addr_rom[15513]='h00003798;  wr_data_rom[15513]='h00000000;
    rd_cycle[15514] = 1'b0;  wr_cycle[15514] = 1'b1;  addr_rom[15514]='h00002d64;  wr_data_rom[15514]='h000039a3;
    rd_cycle[15515] = 1'b0;  wr_cycle[15515] = 1'b1;  addr_rom[15515]='h00003f80;  wr_data_rom[15515]='h00003dee;
    rd_cycle[15516] = 1'b1;  wr_cycle[15516] = 1'b0;  addr_rom[15516]='h00002400;  wr_data_rom[15516]='h00000000;
    rd_cycle[15517] = 1'b1;  wr_cycle[15517] = 1'b0;  addr_rom[15517]='h00000848;  wr_data_rom[15517]='h00000000;
    rd_cycle[15518] = 1'b1;  wr_cycle[15518] = 1'b0;  addr_rom[15518]='h00000a1c;  wr_data_rom[15518]='h00000000;
    rd_cycle[15519] = 1'b1;  wr_cycle[15519] = 1'b0;  addr_rom[15519]='h00000068;  wr_data_rom[15519]='h00000000;
    rd_cycle[15520] = 1'b1;  wr_cycle[15520] = 1'b0;  addr_rom[15520]='h0000239c;  wr_data_rom[15520]='h00000000;
    rd_cycle[15521] = 1'b0;  wr_cycle[15521] = 1'b1;  addr_rom[15521]='h00003fbc;  wr_data_rom[15521]='h00001362;
    rd_cycle[15522] = 1'b1;  wr_cycle[15522] = 1'b0;  addr_rom[15522]='h0000135c;  wr_data_rom[15522]='h00000000;
    rd_cycle[15523] = 1'b0;  wr_cycle[15523] = 1'b1;  addr_rom[15523]='h00001b84;  wr_data_rom[15523]='h0000264e;
    rd_cycle[15524] = 1'b0;  wr_cycle[15524] = 1'b1;  addr_rom[15524]='h00002cb8;  wr_data_rom[15524]='h00001d15;
    rd_cycle[15525] = 1'b0;  wr_cycle[15525] = 1'b1;  addr_rom[15525]='h000008ac;  wr_data_rom[15525]='h0000275a;
    rd_cycle[15526] = 1'b1;  wr_cycle[15526] = 1'b0;  addr_rom[15526]='h00002850;  wr_data_rom[15526]='h00000000;
    rd_cycle[15527] = 1'b1;  wr_cycle[15527] = 1'b0;  addr_rom[15527]='h00002d24;  wr_data_rom[15527]='h00000000;
    rd_cycle[15528] = 1'b0;  wr_cycle[15528] = 1'b1;  addr_rom[15528]='h000025a0;  wr_data_rom[15528]='h00001538;
    rd_cycle[15529] = 1'b1;  wr_cycle[15529] = 1'b0;  addr_rom[15529]='h00001f10;  wr_data_rom[15529]='h00000000;
    rd_cycle[15530] = 1'b0;  wr_cycle[15530] = 1'b1;  addr_rom[15530]='h00000714;  wr_data_rom[15530]='h00001846;
    rd_cycle[15531] = 1'b1;  wr_cycle[15531] = 1'b0;  addr_rom[15531]='h00001eb8;  wr_data_rom[15531]='h00000000;
    rd_cycle[15532] = 1'b1;  wr_cycle[15532] = 1'b0;  addr_rom[15532]='h00003494;  wr_data_rom[15532]='h00000000;
    rd_cycle[15533] = 1'b0;  wr_cycle[15533] = 1'b1;  addr_rom[15533]='h00002990;  wr_data_rom[15533]='h00002ffb;
    rd_cycle[15534] = 1'b1;  wr_cycle[15534] = 1'b0;  addr_rom[15534]='h00003260;  wr_data_rom[15534]='h00000000;
    rd_cycle[15535] = 1'b0;  wr_cycle[15535] = 1'b1;  addr_rom[15535]='h000032a4;  wr_data_rom[15535]='h00003d1f;
    rd_cycle[15536] = 1'b1;  wr_cycle[15536] = 1'b0;  addr_rom[15536]='h0000055c;  wr_data_rom[15536]='h00000000;
    rd_cycle[15537] = 1'b1;  wr_cycle[15537] = 1'b0;  addr_rom[15537]='h00001fd8;  wr_data_rom[15537]='h00000000;
    rd_cycle[15538] = 1'b1;  wr_cycle[15538] = 1'b0;  addr_rom[15538]='h00003a6c;  wr_data_rom[15538]='h00000000;
    rd_cycle[15539] = 1'b0;  wr_cycle[15539] = 1'b1;  addr_rom[15539]='h00000f3c;  wr_data_rom[15539]='h00000206;
    rd_cycle[15540] = 1'b1;  wr_cycle[15540] = 1'b0;  addr_rom[15540]='h00000a14;  wr_data_rom[15540]='h00000000;
    rd_cycle[15541] = 1'b0;  wr_cycle[15541] = 1'b1;  addr_rom[15541]='h00000528;  wr_data_rom[15541]='h00003e49;
    rd_cycle[15542] = 1'b0;  wr_cycle[15542] = 1'b1;  addr_rom[15542]='h00001aac;  wr_data_rom[15542]='h00002990;
    rd_cycle[15543] = 1'b1;  wr_cycle[15543] = 1'b0;  addr_rom[15543]='h00002914;  wr_data_rom[15543]='h00000000;
    rd_cycle[15544] = 1'b1;  wr_cycle[15544] = 1'b0;  addr_rom[15544]='h000002a8;  wr_data_rom[15544]='h00000000;
    rd_cycle[15545] = 1'b0;  wr_cycle[15545] = 1'b1;  addr_rom[15545]='h0000064c;  wr_data_rom[15545]='h00002a82;
    rd_cycle[15546] = 1'b0;  wr_cycle[15546] = 1'b1;  addr_rom[15546]='h00001220;  wr_data_rom[15546]='h00002135;
    rd_cycle[15547] = 1'b0;  wr_cycle[15547] = 1'b1;  addr_rom[15547]='h000012e0;  wr_data_rom[15547]='h000020cc;
    rd_cycle[15548] = 1'b1;  wr_cycle[15548] = 1'b0;  addr_rom[15548]='h00002840;  wr_data_rom[15548]='h00000000;
    rd_cycle[15549] = 1'b0;  wr_cycle[15549] = 1'b1;  addr_rom[15549]='h00002580;  wr_data_rom[15549]='h00000d02;
    rd_cycle[15550] = 1'b0;  wr_cycle[15550] = 1'b1;  addr_rom[15550]='h00002728;  wr_data_rom[15550]='h000036e6;
    rd_cycle[15551] = 1'b0;  wr_cycle[15551] = 1'b1;  addr_rom[15551]='h00001624;  wr_data_rom[15551]='h0000295b;
    rd_cycle[15552] = 1'b0;  wr_cycle[15552] = 1'b1;  addr_rom[15552]='h00002080;  wr_data_rom[15552]='h000017f7;
    rd_cycle[15553] = 1'b0;  wr_cycle[15553] = 1'b1;  addr_rom[15553]='h0000304c;  wr_data_rom[15553]='h00001070;
    rd_cycle[15554] = 1'b0;  wr_cycle[15554] = 1'b1;  addr_rom[15554]='h000009bc;  wr_data_rom[15554]='h00001e6e;
    rd_cycle[15555] = 1'b0;  wr_cycle[15555] = 1'b1;  addr_rom[15555]='h0000393c;  wr_data_rom[15555]='h0000342a;
    rd_cycle[15556] = 1'b1;  wr_cycle[15556] = 1'b0;  addr_rom[15556]='h00002408;  wr_data_rom[15556]='h00000000;
    rd_cycle[15557] = 1'b1;  wr_cycle[15557] = 1'b0;  addr_rom[15557]='h000017ec;  wr_data_rom[15557]='h00000000;
    rd_cycle[15558] = 1'b1;  wr_cycle[15558] = 1'b0;  addr_rom[15558]='h00003804;  wr_data_rom[15558]='h00000000;
    rd_cycle[15559] = 1'b0;  wr_cycle[15559] = 1'b1;  addr_rom[15559]='h00000284;  wr_data_rom[15559]='h0000038d;
    rd_cycle[15560] = 1'b1;  wr_cycle[15560] = 1'b0;  addr_rom[15560]='h000008a4;  wr_data_rom[15560]='h00000000;
    rd_cycle[15561] = 1'b1;  wr_cycle[15561] = 1'b0;  addr_rom[15561]='h00003fac;  wr_data_rom[15561]='h00000000;
    rd_cycle[15562] = 1'b1;  wr_cycle[15562] = 1'b0;  addr_rom[15562]='h000013c0;  wr_data_rom[15562]='h00000000;
    rd_cycle[15563] = 1'b0;  wr_cycle[15563] = 1'b1;  addr_rom[15563]='h000004e8;  wr_data_rom[15563]='h00003c39;
    rd_cycle[15564] = 1'b1;  wr_cycle[15564] = 1'b0;  addr_rom[15564]='h000013cc;  wr_data_rom[15564]='h00000000;
    rd_cycle[15565] = 1'b0;  wr_cycle[15565] = 1'b1;  addr_rom[15565]='h0000126c;  wr_data_rom[15565]='h00003c30;
    rd_cycle[15566] = 1'b0;  wr_cycle[15566] = 1'b1;  addr_rom[15566]='h000004a8;  wr_data_rom[15566]='h000019bf;
    rd_cycle[15567] = 1'b0;  wr_cycle[15567] = 1'b1;  addr_rom[15567]='h00001fc4;  wr_data_rom[15567]='h000038be;
    rd_cycle[15568] = 1'b0;  wr_cycle[15568] = 1'b1;  addr_rom[15568]='h00001174;  wr_data_rom[15568]='h00003e03;
    rd_cycle[15569] = 1'b1;  wr_cycle[15569] = 1'b0;  addr_rom[15569]='h00001f6c;  wr_data_rom[15569]='h00000000;
    rd_cycle[15570] = 1'b0;  wr_cycle[15570] = 1'b1;  addr_rom[15570]='h0000333c;  wr_data_rom[15570]='h000012ba;
    rd_cycle[15571] = 1'b0;  wr_cycle[15571] = 1'b1;  addr_rom[15571]='h00003514;  wr_data_rom[15571]='h000033f0;
    rd_cycle[15572] = 1'b1;  wr_cycle[15572] = 1'b0;  addr_rom[15572]='h00000104;  wr_data_rom[15572]='h00000000;
    rd_cycle[15573] = 1'b1;  wr_cycle[15573] = 1'b0;  addr_rom[15573]='h00003640;  wr_data_rom[15573]='h00000000;
    rd_cycle[15574] = 1'b1;  wr_cycle[15574] = 1'b0;  addr_rom[15574]='h00001678;  wr_data_rom[15574]='h00000000;
    rd_cycle[15575] = 1'b1;  wr_cycle[15575] = 1'b0;  addr_rom[15575]='h0000156c;  wr_data_rom[15575]='h00000000;
    rd_cycle[15576] = 1'b1;  wr_cycle[15576] = 1'b0;  addr_rom[15576]='h000025cc;  wr_data_rom[15576]='h00000000;
    rd_cycle[15577] = 1'b0;  wr_cycle[15577] = 1'b1;  addr_rom[15577]='h00001f20;  wr_data_rom[15577]='h00002cb2;
    rd_cycle[15578] = 1'b0;  wr_cycle[15578] = 1'b1;  addr_rom[15578]='h00001fd8;  wr_data_rom[15578]='h000009df;
    rd_cycle[15579] = 1'b0;  wr_cycle[15579] = 1'b1;  addr_rom[15579]='h00002fcc;  wr_data_rom[15579]='h00000d76;
    rd_cycle[15580] = 1'b1;  wr_cycle[15580] = 1'b0;  addr_rom[15580]='h00002e6c;  wr_data_rom[15580]='h00000000;
    rd_cycle[15581] = 1'b1;  wr_cycle[15581] = 1'b0;  addr_rom[15581]='h00002ae8;  wr_data_rom[15581]='h00000000;
    rd_cycle[15582] = 1'b1;  wr_cycle[15582] = 1'b0;  addr_rom[15582]='h00003474;  wr_data_rom[15582]='h00000000;
    rd_cycle[15583] = 1'b0;  wr_cycle[15583] = 1'b1;  addr_rom[15583]='h00002824;  wr_data_rom[15583]='h0000166e;
    rd_cycle[15584] = 1'b1;  wr_cycle[15584] = 1'b0;  addr_rom[15584]='h00003a9c;  wr_data_rom[15584]='h00000000;
    rd_cycle[15585] = 1'b1;  wr_cycle[15585] = 1'b0;  addr_rom[15585]='h000000c8;  wr_data_rom[15585]='h00000000;
    rd_cycle[15586] = 1'b0;  wr_cycle[15586] = 1'b1;  addr_rom[15586]='h00001e60;  wr_data_rom[15586]='h00002878;
    rd_cycle[15587] = 1'b0;  wr_cycle[15587] = 1'b1;  addr_rom[15587]='h00001dd8;  wr_data_rom[15587]='h00000cd7;
    rd_cycle[15588] = 1'b1;  wr_cycle[15588] = 1'b0;  addr_rom[15588]='h000025e4;  wr_data_rom[15588]='h00000000;
    rd_cycle[15589] = 1'b0;  wr_cycle[15589] = 1'b1;  addr_rom[15589]='h000025d4;  wr_data_rom[15589]='h00003131;
    rd_cycle[15590] = 1'b1;  wr_cycle[15590] = 1'b0;  addr_rom[15590]='h00001444;  wr_data_rom[15590]='h00000000;
    rd_cycle[15591] = 1'b0;  wr_cycle[15591] = 1'b1;  addr_rom[15591]='h00000708;  wr_data_rom[15591]='h00000b82;
    rd_cycle[15592] = 1'b1;  wr_cycle[15592] = 1'b0;  addr_rom[15592]='h000004b4;  wr_data_rom[15592]='h00000000;
    rd_cycle[15593] = 1'b0;  wr_cycle[15593] = 1'b1;  addr_rom[15593]='h00003adc;  wr_data_rom[15593]='h00000640;
    rd_cycle[15594] = 1'b1;  wr_cycle[15594] = 1'b0;  addr_rom[15594]='h00003bd4;  wr_data_rom[15594]='h00000000;
    rd_cycle[15595] = 1'b0;  wr_cycle[15595] = 1'b1;  addr_rom[15595]='h00001ef8;  wr_data_rom[15595]='h000006ff;
    rd_cycle[15596] = 1'b0;  wr_cycle[15596] = 1'b1;  addr_rom[15596]='h00001318;  wr_data_rom[15596]='h00002daf;
    rd_cycle[15597] = 1'b1;  wr_cycle[15597] = 1'b0;  addr_rom[15597]='h00001e04;  wr_data_rom[15597]='h00000000;
    rd_cycle[15598] = 1'b0;  wr_cycle[15598] = 1'b1;  addr_rom[15598]='h00003ae0;  wr_data_rom[15598]='h00003425;
    rd_cycle[15599] = 1'b0;  wr_cycle[15599] = 1'b1;  addr_rom[15599]='h000033f4;  wr_data_rom[15599]='h00002f5a;
    rd_cycle[15600] = 1'b0;  wr_cycle[15600] = 1'b1;  addr_rom[15600]='h0000321c;  wr_data_rom[15600]='h00000776;
    rd_cycle[15601] = 1'b1;  wr_cycle[15601] = 1'b0;  addr_rom[15601]='h000021d8;  wr_data_rom[15601]='h00000000;
    rd_cycle[15602] = 1'b0;  wr_cycle[15602] = 1'b1;  addr_rom[15602]='h0000309c;  wr_data_rom[15602]='h000028c1;
    rd_cycle[15603] = 1'b1;  wr_cycle[15603] = 1'b0;  addr_rom[15603]='h000009dc;  wr_data_rom[15603]='h00000000;
    rd_cycle[15604] = 1'b1;  wr_cycle[15604] = 1'b0;  addr_rom[15604]='h00002090;  wr_data_rom[15604]='h00000000;
    rd_cycle[15605] = 1'b0;  wr_cycle[15605] = 1'b1;  addr_rom[15605]='h0000277c;  wr_data_rom[15605]='h000021c7;
    rd_cycle[15606] = 1'b0;  wr_cycle[15606] = 1'b1;  addr_rom[15606]='h00003c7c;  wr_data_rom[15606]='h00000893;
    rd_cycle[15607] = 1'b1;  wr_cycle[15607] = 1'b0;  addr_rom[15607]='h00002aa4;  wr_data_rom[15607]='h00000000;
    rd_cycle[15608] = 1'b0;  wr_cycle[15608] = 1'b1;  addr_rom[15608]='h000030e8;  wr_data_rom[15608]='h00000d4e;
    rd_cycle[15609] = 1'b0;  wr_cycle[15609] = 1'b1;  addr_rom[15609]='h00001ea4;  wr_data_rom[15609]='h00003b64;
    rd_cycle[15610] = 1'b1;  wr_cycle[15610] = 1'b0;  addr_rom[15610]='h00003874;  wr_data_rom[15610]='h00000000;
    rd_cycle[15611] = 1'b1;  wr_cycle[15611] = 1'b0;  addr_rom[15611]='h000030f4;  wr_data_rom[15611]='h00000000;
    rd_cycle[15612] = 1'b1;  wr_cycle[15612] = 1'b0;  addr_rom[15612]='h00002758;  wr_data_rom[15612]='h00000000;
    rd_cycle[15613] = 1'b1;  wr_cycle[15613] = 1'b0;  addr_rom[15613]='h000004c8;  wr_data_rom[15613]='h00000000;
    rd_cycle[15614] = 1'b0;  wr_cycle[15614] = 1'b1;  addr_rom[15614]='h000038e4;  wr_data_rom[15614]='h0000246c;
    rd_cycle[15615] = 1'b1;  wr_cycle[15615] = 1'b0;  addr_rom[15615]='h0000284c;  wr_data_rom[15615]='h00000000;
    rd_cycle[15616] = 1'b0;  wr_cycle[15616] = 1'b1;  addr_rom[15616]='h00001660;  wr_data_rom[15616]='h00003e22;
    rd_cycle[15617] = 1'b1;  wr_cycle[15617] = 1'b0;  addr_rom[15617]='h00002360;  wr_data_rom[15617]='h00000000;
    rd_cycle[15618] = 1'b1;  wr_cycle[15618] = 1'b0;  addr_rom[15618]='h000027ac;  wr_data_rom[15618]='h00000000;
    rd_cycle[15619] = 1'b0;  wr_cycle[15619] = 1'b1;  addr_rom[15619]='h00003714;  wr_data_rom[15619]='h00000218;
    rd_cycle[15620] = 1'b0;  wr_cycle[15620] = 1'b1;  addr_rom[15620]='h00003094;  wr_data_rom[15620]='h000019a0;
    rd_cycle[15621] = 1'b0;  wr_cycle[15621] = 1'b1;  addr_rom[15621]='h000033b8;  wr_data_rom[15621]='h00000081;
    rd_cycle[15622] = 1'b0;  wr_cycle[15622] = 1'b1;  addr_rom[15622]='h00003acc;  wr_data_rom[15622]='h00002035;
    rd_cycle[15623] = 1'b0;  wr_cycle[15623] = 1'b1;  addr_rom[15623]='h000006f4;  wr_data_rom[15623]='h00002a9e;
    rd_cycle[15624] = 1'b0;  wr_cycle[15624] = 1'b1;  addr_rom[15624]='h00002e08;  wr_data_rom[15624]='h00002bc6;
    rd_cycle[15625] = 1'b0;  wr_cycle[15625] = 1'b1;  addr_rom[15625]='h00002818;  wr_data_rom[15625]='h000011f0;
    rd_cycle[15626] = 1'b1;  wr_cycle[15626] = 1'b0;  addr_rom[15626]='h0000009c;  wr_data_rom[15626]='h00000000;
    rd_cycle[15627] = 1'b1;  wr_cycle[15627] = 1'b0;  addr_rom[15627]='h00001c38;  wr_data_rom[15627]='h00000000;
    rd_cycle[15628] = 1'b1;  wr_cycle[15628] = 1'b0;  addr_rom[15628]='h00000dc8;  wr_data_rom[15628]='h00000000;
    rd_cycle[15629] = 1'b0;  wr_cycle[15629] = 1'b1;  addr_rom[15629]='h000038fc;  wr_data_rom[15629]='h00000656;
    rd_cycle[15630] = 1'b0;  wr_cycle[15630] = 1'b1;  addr_rom[15630]='h00001b14;  wr_data_rom[15630]='h00003fcf;
    rd_cycle[15631] = 1'b1;  wr_cycle[15631] = 1'b0;  addr_rom[15631]='h00003e1c;  wr_data_rom[15631]='h00000000;
    rd_cycle[15632] = 1'b0;  wr_cycle[15632] = 1'b1;  addr_rom[15632]='h00001248;  wr_data_rom[15632]='h00003ecb;
    rd_cycle[15633] = 1'b0;  wr_cycle[15633] = 1'b1;  addr_rom[15633]='h00000bec;  wr_data_rom[15633]='h00002a1b;
    rd_cycle[15634] = 1'b1;  wr_cycle[15634] = 1'b0;  addr_rom[15634]='h00001ef8;  wr_data_rom[15634]='h00000000;
    rd_cycle[15635] = 1'b0;  wr_cycle[15635] = 1'b1;  addr_rom[15635]='h00001a7c;  wr_data_rom[15635]='h00001e53;
    rd_cycle[15636] = 1'b0;  wr_cycle[15636] = 1'b1;  addr_rom[15636]='h00000e6c;  wr_data_rom[15636]='h0000073a;
    rd_cycle[15637] = 1'b1;  wr_cycle[15637] = 1'b0;  addr_rom[15637]='h000025f8;  wr_data_rom[15637]='h00000000;
    rd_cycle[15638] = 1'b1;  wr_cycle[15638] = 1'b0;  addr_rom[15638]='h0000279c;  wr_data_rom[15638]='h00000000;
    rd_cycle[15639] = 1'b1;  wr_cycle[15639] = 1'b0;  addr_rom[15639]='h00002e9c;  wr_data_rom[15639]='h00000000;
    rd_cycle[15640] = 1'b0;  wr_cycle[15640] = 1'b1;  addr_rom[15640]='h00002388;  wr_data_rom[15640]='h0000268d;
    rd_cycle[15641] = 1'b0;  wr_cycle[15641] = 1'b1;  addr_rom[15641]='h00000030;  wr_data_rom[15641]='h00003f11;
    rd_cycle[15642] = 1'b0;  wr_cycle[15642] = 1'b1;  addr_rom[15642]='h00003bd4;  wr_data_rom[15642]='h00003fb6;
    rd_cycle[15643] = 1'b1;  wr_cycle[15643] = 1'b0;  addr_rom[15643]='h000029ac;  wr_data_rom[15643]='h00000000;
    rd_cycle[15644] = 1'b1;  wr_cycle[15644] = 1'b0;  addr_rom[15644]='h00000008;  wr_data_rom[15644]='h00000000;
    rd_cycle[15645] = 1'b0;  wr_cycle[15645] = 1'b1;  addr_rom[15645]='h000009b8;  wr_data_rom[15645]='h00000a3e;
    rd_cycle[15646] = 1'b0;  wr_cycle[15646] = 1'b1;  addr_rom[15646]='h00002ca0;  wr_data_rom[15646]='h0000395f;
    rd_cycle[15647] = 1'b0;  wr_cycle[15647] = 1'b1;  addr_rom[15647]='h00001e3c;  wr_data_rom[15647]='h00001ab8;
    rd_cycle[15648] = 1'b0;  wr_cycle[15648] = 1'b1;  addr_rom[15648]='h000008c4;  wr_data_rom[15648]='h00001d1f;
    rd_cycle[15649] = 1'b0;  wr_cycle[15649] = 1'b1;  addr_rom[15649]='h000009d8;  wr_data_rom[15649]='h00000b8d;
    rd_cycle[15650] = 1'b0;  wr_cycle[15650] = 1'b1;  addr_rom[15650]='h00003144;  wr_data_rom[15650]='h000028e8;
    rd_cycle[15651] = 1'b1;  wr_cycle[15651] = 1'b0;  addr_rom[15651]='h0000163c;  wr_data_rom[15651]='h00000000;
    rd_cycle[15652] = 1'b0;  wr_cycle[15652] = 1'b1;  addr_rom[15652]='h00002290;  wr_data_rom[15652]='h00000bd9;
    rd_cycle[15653] = 1'b0;  wr_cycle[15653] = 1'b1;  addr_rom[15653]='h00001580;  wr_data_rom[15653]='h000036f0;
    rd_cycle[15654] = 1'b0;  wr_cycle[15654] = 1'b1;  addr_rom[15654]='h00002668;  wr_data_rom[15654]='h0000047c;
    rd_cycle[15655] = 1'b1;  wr_cycle[15655] = 1'b0;  addr_rom[15655]='h00000bcc;  wr_data_rom[15655]='h00000000;
    rd_cycle[15656] = 1'b0;  wr_cycle[15656] = 1'b1;  addr_rom[15656]='h00001828;  wr_data_rom[15656]='h00002f9a;
    rd_cycle[15657] = 1'b1;  wr_cycle[15657] = 1'b0;  addr_rom[15657]='h00000b34;  wr_data_rom[15657]='h00000000;
    rd_cycle[15658] = 1'b0;  wr_cycle[15658] = 1'b1;  addr_rom[15658]='h00000d98;  wr_data_rom[15658]='h00003995;
    rd_cycle[15659] = 1'b0;  wr_cycle[15659] = 1'b1;  addr_rom[15659]='h00000550;  wr_data_rom[15659]='h00000dfa;
    rd_cycle[15660] = 1'b0;  wr_cycle[15660] = 1'b1;  addr_rom[15660]='h00000154;  wr_data_rom[15660]='h000039e6;
    rd_cycle[15661] = 1'b1;  wr_cycle[15661] = 1'b0;  addr_rom[15661]='h000030f4;  wr_data_rom[15661]='h00000000;
    rd_cycle[15662] = 1'b1;  wr_cycle[15662] = 1'b0;  addr_rom[15662]='h00002d54;  wr_data_rom[15662]='h00000000;
    rd_cycle[15663] = 1'b0;  wr_cycle[15663] = 1'b1;  addr_rom[15663]='h00003d28;  wr_data_rom[15663]='h000025e5;
    rd_cycle[15664] = 1'b0;  wr_cycle[15664] = 1'b1;  addr_rom[15664]='h00003d50;  wr_data_rom[15664]='h00002947;
    rd_cycle[15665] = 1'b1;  wr_cycle[15665] = 1'b0;  addr_rom[15665]='h0000184c;  wr_data_rom[15665]='h00000000;
    rd_cycle[15666] = 1'b1;  wr_cycle[15666] = 1'b0;  addr_rom[15666]='h00003c34;  wr_data_rom[15666]='h00000000;
    rd_cycle[15667] = 1'b0;  wr_cycle[15667] = 1'b1;  addr_rom[15667]='h00003f4c;  wr_data_rom[15667]='h00003dd5;
    rd_cycle[15668] = 1'b0;  wr_cycle[15668] = 1'b1;  addr_rom[15668]='h00002b20;  wr_data_rom[15668]='h00002595;
    rd_cycle[15669] = 1'b1;  wr_cycle[15669] = 1'b0;  addr_rom[15669]='h00003cd4;  wr_data_rom[15669]='h00000000;
    rd_cycle[15670] = 1'b0;  wr_cycle[15670] = 1'b1;  addr_rom[15670]='h000001fc;  wr_data_rom[15670]='h00003d50;
    rd_cycle[15671] = 1'b1;  wr_cycle[15671] = 1'b0;  addr_rom[15671]='h00003568;  wr_data_rom[15671]='h00000000;
    rd_cycle[15672] = 1'b1;  wr_cycle[15672] = 1'b0;  addr_rom[15672]='h00003380;  wr_data_rom[15672]='h00000000;
    rd_cycle[15673] = 1'b0;  wr_cycle[15673] = 1'b1;  addr_rom[15673]='h0000231c;  wr_data_rom[15673]='h00001251;
    rd_cycle[15674] = 1'b0;  wr_cycle[15674] = 1'b1;  addr_rom[15674]='h00000aac;  wr_data_rom[15674]='h00003e94;
    rd_cycle[15675] = 1'b1;  wr_cycle[15675] = 1'b0;  addr_rom[15675]='h000015b8;  wr_data_rom[15675]='h00000000;
    rd_cycle[15676] = 1'b0;  wr_cycle[15676] = 1'b1;  addr_rom[15676]='h000035f4;  wr_data_rom[15676]='h00002ad8;
    rd_cycle[15677] = 1'b1;  wr_cycle[15677] = 1'b0;  addr_rom[15677]='h00001da0;  wr_data_rom[15677]='h00000000;
    rd_cycle[15678] = 1'b1;  wr_cycle[15678] = 1'b0;  addr_rom[15678]='h00000ab8;  wr_data_rom[15678]='h00000000;
    rd_cycle[15679] = 1'b1;  wr_cycle[15679] = 1'b0;  addr_rom[15679]='h000024fc;  wr_data_rom[15679]='h00000000;
    rd_cycle[15680] = 1'b0;  wr_cycle[15680] = 1'b1;  addr_rom[15680]='h00001a70;  wr_data_rom[15680]='h0000078f;
    rd_cycle[15681] = 1'b1;  wr_cycle[15681] = 1'b0;  addr_rom[15681]='h00003430;  wr_data_rom[15681]='h00000000;
    rd_cycle[15682] = 1'b0;  wr_cycle[15682] = 1'b1;  addr_rom[15682]='h00000244;  wr_data_rom[15682]='h0000221f;
    rd_cycle[15683] = 1'b1;  wr_cycle[15683] = 1'b0;  addr_rom[15683]='h00003a6c;  wr_data_rom[15683]='h00000000;
    rd_cycle[15684] = 1'b1;  wr_cycle[15684] = 1'b0;  addr_rom[15684]='h00000250;  wr_data_rom[15684]='h00000000;
    rd_cycle[15685] = 1'b1;  wr_cycle[15685] = 1'b0;  addr_rom[15685]='h000024d0;  wr_data_rom[15685]='h00000000;
    rd_cycle[15686] = 1'b0;  wr_cycle[15686] = 1'b1;  addr_rom[15686]='h000035b4;  wr_data_rom[15686]='h000022b4;
    rd_cycle[15687] = 1'b0;  wr_cycle[15687] = 1'b1;  addr_rom[15687]='h00003f5c;  wr_data_rom[15687]='h000038b5;
    rd_cycle[15688] = 1'b0;  wr_cycle[15688] = 1'b1;  addr_rom[15688]='h00000b20;  wr_data_rom[15688]='h000006c7;
    rd_cycle[15689] = 1'b0;  wr_cycle[15689] = 1'b1;  addr_rom[15689]='h00002774;  wr_data_rom[15689]='h000039fe;
    rd_cycle[15690] = 1'b0;  wr_cycle[15690] = 1'b1;  addr_rom[15690]='h00003f20;  wr_data_rom[15690]='h00003d4b;
    rd_cycle[15691] = 1'b0;  wr_cycle[15691] = 1'b1;  addr_rom[15691]='h000018e8;  wr_data_rom[15691]='h00000be7;
    rd_cycle[15692] = 1'b0;  wr_cycle[15692] = 1'b1;  addr_rom[15692]='h00002810;  wr_data_rom[15692]='h00001097;
    rd_cycle[15693] = 1'b0;  wr_cycle[15693] = 1'b1;  addr_rom[15693]='h000017c4;  wr_data_rom[15693]='h0000054d;
    rd_cycle[15694] = 1'b0;  wr_cycle[15694] = 1'b1;  addr_rom[15694]='h00000ec4;  wr_data_rom[15694]='h000010a5;
    rd_cycle[15695] = 1'b0;  wr_cycle[15695] = 1'b1;  addr_rom[15695]='h0000241c;  wr_data_rom[15695]='h0000129f;
    rd_cycle[15696] = 1'b0;  wr_cycle[15696] = 1'b1;  addr_rom[15696]='h00003734;  wr_data_rom[15696]='h00003772;
    rd_cycle[15697] = 1'b1;  wr_cycle[15697] = 1'b0;  addr_rom[15697]='h000014e8;  wr_data_rom[15697]='h00000000;
    rd_cycle[15698] = 1'b1;  wr_cycle[15698] = 1'b0;  addr_rom[15698]='h00003140;  wr_data_rom[15698]='h00000000;
    rd_cycle[15699] = 1'b1;  wr_cycle[15699] = 1'b0;  addr_rom[15699]='h00003144;  wr_data_rom[15699]='h00000000;
    rd_cycle[15700] = 1'b1;  wr_cycle[15700] = 1'b0;  addr_rom[15700]='h00001614;  wr_data_rom[15700]='h00000000;
    rd_cycle[15701] = 1'b0;  wr_cycle[15701] = 1'b1;  addr_rom[15701]='h00003994;  wr_data_rom[15701]='h00000be2;
    rd_cycle[15702] = 1'b1;  wr_cycle[15702] = 1'b0;  addr_rom[15702]='h00000828;  wr_data_rom[15702]='h00000000;
    rd_cycle[15703] = 1'b1;  wr_cycle[15703] = 1'b0;  addr_rom[15703]='h000003bc;  wr_data_rom[15703]='h00000000;
    rd_cycle[15704] = 1'b0;  wr_cycle[15704] = 1'b1;  addr_rom[15704]='h00000208;  wr_data_rom[15704]='h0000095d;
    rd_cycle[15705] = 1'b0;  wr_cycle[15705] = 1'b1;  addr_rom[15705]='h0000043c;  wr_data_rom[15705]='h00003553;
    rd_cycle[15706] = 1'b0;  wr_cycle[15706] = 1'b1;  addr_rom[15706]='h000027e4;  wr_data_rom[15706]='h00002967;
    rd_cycle[15707] = 1'b1;  wr_cycle[15707] = 1'b0;  addr_rom[15707]='h00003ae4;  wr_data_rom[15707]='h00000000;
    rd_cycle[15708] = 1'b0;  wr_cycle[15708] = 1'b1;  addr_rom[15708]='h000016e8;  wr_data_rom[15708]='h00001f26;
    rd_cycle[15709] = 1'b1;  wr_cycle[15709] = 1'b0;  addr_rom[15709]='h0000111c;  wr_data_rom[15709]='h00000000;
    rd_cycle[15710] = 1'b0;  wr_cycle[15710] = 1'b1;  addr_rom[15710]='h000005b8;  wr_data_rom[15710]='h000011d3;
    rd_cycle[15711] = 1'b1;  wr_cycle[15711] = 1'b0;  addr_rom[15711]='h00001158;  wr_data_rom[15711]='h00000000;
    rd_cycle[15712] = 1'b0;  wr_cycle[15712] = 1'b1;  addr_rom[15712]='h000008b4;  wr_data_rom[15712]='h00000613;
    rd_cycle[15713] = 1'b1;  wr_cycle[15713] = 1'b0;  addr_rom[15713]='h00000060;  wr_data_rom[15713]='h00000000;
    rd_cycle[15714] = 1'b0;  wr_cycle[15714] = 1'b1;  addr_rom[15714]='h00003510;  wr_data_rom[15714]='h00003740;
    rd_cycle[15715] = 1'b0;  wr_cycle[15715] = 1'b1;  addr_rom[15715]='h00000e18;  wr_data_rom[15715]='h00001840;
    rd_cycle[15716] = 1'b1;  wr_cycle[15716] = 1'b0;  addr_rom[15716]='h00001324;  wr_data_rom[15716]='h00000000;
    rd_cycle[15717] = 1'b0;  wr_cycle[15717] = 1'b1;  addr_rom[15717]='h00000978;  wr_data_rom[15717]='h000007b4;
    rd_cycle[15718] = 1'b0;  wr_cycle[15718] = 1'b1;  addr_rom[15718]='h00001860;  wr_data_rom[15718]='h00003f18;
    rd_cycle[15719] = 1'b1;  wr_cycle[15719] = 1'b0;  addr_rom[15719]='h000036c0;  wr_data_rom[15719]='h00000000;
    rd_cycle[15720] = 1'b0;  wr_cycle[15720] = 1'b1;  addr_rom[15720]='h00000078;  wr_data_rom[15720]='h000011ae;
    rd_cycle[15721] = 1'b1;  wr_cycle[15721] = 1'b0;  addr_rom[15721]='h00001928;  wr_data_rom[15721]='h00000000;
    rd_cycle[15722] = 1'b1;  wr_cycle[15722] = 1'b0;  addr_rom[15722]='h00000d0c;  wr_data_rom[15722]='h00000000;
    rd_cycle[15723] = 1'b1;  wr_cycle[15723] = 1'b0;  addr_rom[15723]='h000012b8;  wr_data_rom[15723]='h00000000;
    rd_cycle[15724] = 1'b1;  wr_cycle[15724] = 1'b0;  addr_rom[15724]='h00001ec0;  wr_data_rom[15724]='h00000000;
    rd_cycle[15725] = 1'b0;  wr_cycle[15725] = 1'b1;  addr_rom[15725]='h00000d0c;  wr_data_rom[15725]='h00000ec1;
    rd_cycle[15726] = 1'b1;  wr_cycle[15726] = 1'b0;  addr_rom[15726]='h00003244;  wr_data_rom[15726]='h00000000;
    rd_cycle[15727] = 1'b0;  wr_cycle[15727] = 1'b1;  addr_rom[15727]='h00003bf8;  wr_data_rom[15727]='h00001be8;
    rd_cycle[15728] = 1'b1;  wr_cycle[15728] = 1'b0;  addr_rom[15728]='h00001128;  wr_data_rom[15728]='h00000000;
    rd_cycle[15729] = 1'b1;  wr_cycle[15729] = 1'b0;  addr_rom[15729]='h000014ac;  wr_data_rom[15729]='h00000000;
    rd_cycle[15730] = 1'b1;  wr_cycle[15730] = 1'b0;  addr_rom[15730]='h000025ac;  wr_data_rom[15730]='h00000000;
    rd_cycle[15731] = 1'b0;  wr_cycle[15731] = 1'b1;  addr_rom[15731]='h00003efc;  wr_data_rom[15731]='h00003022;
    rd_cycle[15732] = 1'b1;  wr_cycle[15732] = 1'b0;  addr_rom[15732]='h00001ff0;  wr_data_rom[15732]='h00000000;
    rd_cycle[15733] = 1'b1;  wr_cycle[15733] = 1'b0;  addr_rom[15733]='h0000087c;  wr_data_rom[15733]='h00000000;
    rd_cycle[15734] = 1'b0;  wr_cycle[15734] = 1'b1;  addr_rom[15734]='h000037c4;  wr_data_rom[15734]='h000015b5;
    rd_cycle[15735] = 1'b1;  wr_cycle[15735] = 1'b0;  addr_rom[15735]='h00001d9c;  wr_data_rom[15735]='h00000000;
    rd_cycle[15736] = 1'b1;  wr_cycle[15736] = 1'b0;  addr_rom[15736]='h000027f0;  wr_data_rom[15736]='h00000000;
    rd_cycle[15737] = 1'b0;  wr_cycle[15737] = 1'b1;  addr_rom[15737]='h00003d44;  wr_data_rom[15737]='h000010cf;
    rd_cycle[15738] = 1'b1;  wr_cycle[15738] = 1'b0;  addr_rom[15738]='h00003498;  wr_data_rom[15738]='h00000000;
    rd_cycle[15739] = 1'b1;  wr_cycle[15739] = 1'b0;  addr_rom[15739]='h0000141c;  wr_data_rom[15739]='h00000000;
    rd_cycle[15740] = 1'b0;  wr_cycle[15740] = 1'b1;  addr_rom[15740]='h000016c0;  wr_data_rom[15740]='h00000a5c;
    rd_cycle[15741] = 1'b0;  wr_cycle[15741] = 1'b1;  addr_rom[15741]='h00001fbc;  wr_data_rom[15741]='h00001411;
    rd_cycle[15742] = 1'b1;  wr_cycle[15742] = 1'b0;  addr_rom[15742]='h00001b68;  wr_data_rom[15742]='h00000000;
    rd_cycle[15743] = 1'b1;  wr_cycle[15743] = 1'b0;  addr_rom[15743]='h000032b8;  wr_data_rom[15743]='h00000000;
    rd_cycle[15744] = 1'b1;  wr_cycle[15744] = 1'b0;  addr_rom[15744]='h00003f10;  wr_data_rom[15744]='h00000000;
    rd_cycle[15745] = 1'b0;  wr_cycle[15745] = 1'b1;  addr_rom[15745]='h00003b00;  wr_data_rom[15745]='h00000029;
    rd_cycle[15746] = 1'b0;  wr_cycle[15746] = 1'b1;  addr_rom[15746]='h00003500;  wr_data_rom[15746]='h0000274c;
    rd_cycle[15747] = 1'b0;  wr_cycle[15747] = 1'b1;  addr_rom[15747]='h00001cdc;  wr_data_rom[15747]='h00002244;
    rd_cycle[15748] = 1'b1;  wr_cycle[15748] = 1'b0;  addr_rom[15748]='h00003708;  wr_data_rom[15748]='h00000000;
    rd_cycle[15749] = 1'b1;  wr_cycle[15749] = 1'b0;  addr_rom[15749]='h000019ec;  wr_data_rom[15749]='h00000000;
    rd_cycle[15750] = 1'b1;  wr_cycle[15750] = 1'b0;  addr_rom[15750]='h0000084c;  wr_data_rom[15750]='h00000000;
    rd_cycle[15751] = 1'b0;  wr_cycle[15751] = 1'b1;  addr_rom[15751]='h00002f1c;  wr_data_rom[15751]='h000020d7;
    rd_cycle[15752] = 1'b0;  wr_cycle[15752] = 1'b1;  addr_rom[15752]='h0000098c;  wr_data_rom[15752]='h0000392a;
    rd_cycle[15753] = 1'b0;  wr_cycle[15753] = 1'b1;  addr_rom[15753]='h0000155c;  wr_data_rom[15753]='h00000387;
    rd_cycle[15754] = 1'b0;  wr_cycle[15754] = 1'b1;  addr_rom[15754]='h00001c90;  wr_data_rom[15754]='h000015f7;
    rd_cycle[15755] = 1'b0;  wr_cycle[15755] = 1'b1;  addr_rom[15755]='h000031f4;  wr_data_rom[15755]='h00002c0e;
    rd_cycle[15756] = 1'b1;  wr_cycle[15756] = 1'b0;  addr_rom[15756]='h000037a0;  wr_data_rom[15756]='h00000000;
    rd_cycle[15757] = 1'b1;  wr_cycle[15757] = 1'b0;  addr_rom[15757]='h00000f40;  wr_data_rom[15757]='h00000000;
    rd_cycle[15758] = 1'b1;  wr_cycle[15758] = 1'b0;  addr_rom[15758]='h00003ac0;  wr_data_rom[15758]='h00000000;
    rd_cycle[15759] = 1'b1;  wr_cycle[15759] = 1'b0;  addr_rom[15759]='h000015b4;  wr_data_rom[15759]='h00000000;
    rd_cycle[15760] = 1'b0;  wr_cycle[15760] = 1'b1;  addr_rom[15760]='h000038d4;  wr_data_rom[15760]='h00000e93;
    rd_cycle[15761] = 1'b0;  wr_cycle[15761] = 1'b1;  addr_rom[15761]='h00000094;  wr_data_rom[15761]='h00002797;
    rd_cycle[15762] = 1'b1;  wr_cycle[15762] = 1'b0;  addr_rom[15762]='h000030a0;  wr_data_rom[15762]='h00000000;
    rd_cycle[15763] = 1'b1;  wr_cycle[15763] = 1'b0;  addr_rom[15763]='h00000164;  wr_data_rom[15763]='h00000000;
    rd_cycle[15764] = 1'b1;  wr_cycle[15764] = 1'b0;  addr_rom[15764]='h000018e0;  wr_data_rom[15764]='h00000000;
    rd_cycle[15765] = 1'b0;  wr_cycle[15765] = 1'b1;  addr_rom[15765]='h00003368;  wr_data_rom[15765]='h00001303;
    rd_cycle[15766] = 1'b1;  wr_cycle[15766] = 1'b0;  addr_rom[15766]='h00001160;  wr_data_rom[15766]='h00000000;
    rd_cycle[15767] = 1'b1;  wr_cycle[15767] = 1'b0;  addr_rom[15767]='h00002144;  wr_data_rom[15767]='h00000000;
    rd_cycle[15768] = 1'b1;  wr_cycle[15768] = 1'b0;  addr_rom[15768]='h00003ea0;  wr_data_rom[15768]='h00000000;
    rd_cycle[15769] = 1'b0;  wr_cycle[15769] = 1'b1;  addr_rom[15769]='h0000017c;  wr_data_rom[15769]='h000010e9;
    rd_cycle[15770] = 1'b0;  wr_cycle[15770] = 1'b1;  addr_rom[15770]='h00003e7c;  wr_data_rom[15770]='h00000cb5;
    rd_cycle[15771] = 1'b0;  wr_cycle[15771] = 1'b1;  addr_rom[15771]='h00002494;  wr_data_rom[15771]='h000029ad;
    rd_cycle[15772] = 1'b0;  wr_cycle[15772] = 1'b1;  addr_rom[15772]='h000005d4;  wr_data_rom[15772]='h00001a83;
    rd_cycle[15773] = 1'b0;  wr_cycle[15773] = 1'b1;  addr_rom[15773]='h00001324;  wr_data_rom[15773]='h00003361;
    rd_cycle[15774] = 1'b0;  wr_cycle[15774] = 1'b1;  addr_rom[15774]='h00003040;  wr_data_rom[15774]='h0000226d;
    rd_cycle[15775] = 1'b1;  wr_cycle[15775] = 1'b0;  addr_rom[15775]='h0000021c;  wr_data_rom[15775]='h00000000;
    rd_cycle[15776] = 1'b0;  wr_cycle[15776] = 1'b1;  addr_rom[15776]='h00001700;  wr_data_rom[15776]='h00000add;
    rd_cycle[15777] = 1'b1;  wr_cycle[15777] = 1'b0;  addr_rom[15777]='h00000718;  wr_data_rom[15777]='h00000000;
    rd_cycle[15778] = 1'b1;  wr_cycle[15778] = 1'b0;  addr_rom[15778]='h00002228;  wr_data_rom[15778]='h00000000;
    rd_cycle[15779] = 1'b0;  wr_cycle[15779] = 1'b1;  addr_rom[15779]='h000004e4;  wr_data_rom[15779]='h00001ca4;
    rd_cycle[15780] = 1'b0;  wr_cycle[15780] = 1'b1;  addr_rom[15780]='h000023d0;  wr_data_rom[15780]='h00003b0e;
    rd_cycle[15781] = 1'b1;  wr_cycle[15781] = 1'b0;  addr_rom[15781]='h00002080;  wr_data_rom[15781]='h00000000;
    rd_cycle[15782] = 1'b0;  wr_cycle[15782] = 1'b1;  addr_rom[15782]='h000030a8;  wr_data_rom[15782]='h0000362d;
    rd_cycle[15783] = 1'b1;  wr_cycle[15783] = 1'b0;  addr_rom[15783]='h00001c3c;  wr_data_rom[15783]='h00000000;
    rd_cycle[15784] = 1'b1;  wr_cycle[15784] = 1'b0;  addr_rom[15784]='h00003f74;  wr_data_rom[15784]='h00000000;
    rd_cycle[15785] = 1'b0;  wr_cycle[15785] = 1'b1;  addr_rom[15785]='h0000166c;  wr_data_rom[15785]='h00001af7;
    rd_cycle[15786] = 1'b1;  wr_cycle[15786] = 1'b0;  addr_rom[15786]='h00003b7c;  wr_data_rom[15786]='h00000000;
    rd_cycle[15787] = 1'b1;  wr_cycle[15787] = 1'b0;  addr_rom[15787]='h00003730;  wr_data_rom[15787]='h00000000;
    rd_cycle[15788] = 1'b1;  wr_cycle[15788] = 1'b0;  addr_rom[15788]='h00003168;  wr_data_rom[15788]='h00000000;
    rd_cycle[15789] = 1'b1;  wr_cycle[15789] = 1'b0;  addr_rom[15789]='h00000710;  wr_data_rom[15789]='h00000000;
    rd_cycle[15790] = 1'b0;  wr_cycle[15790] = 1'b1;  addr_rom[15790]='h00003b98;  wr_data_rom[15790]='h00000d55;
    rd_cycle[15791] = 1'b1;  wr_cycle[15791] = 1'b0;  addr_rom[15791]='h00001c30;  wr_data_rom[15791]='h00000000;
    rd_cycle[15792] = 1'b1;  wr_cycle[15792] = 1'b0;  addr_rom[15792]='h00000b88;  wr_data_rom[15792]='h00000000;
    rd_cycle[15793] = 1'b1;  wr_cycle[15793] = 1'b0;  addr_rom[15793]='h00003b44;  wr_data_rom[15793]='h00000000;
    rd_cycle[15794] = 1'b0;  wr_cycle[15794] = 1'b1;  addr_rom[15794]='h000029e0;  wr_data_rom[15794]='h00002158;
    rd_cycle[15795] = 1'b1;  wr_cycle[15795] = 1'b0;  addr_rom[15795]='h000019c4;  wr_data_rom[15795]='h00000000;
    rd_cycle[15796] = 1'b0;  wr_cycle[15796] = 1'b1;  addr_rom[15796]='h000002c8;  wr_data_rom[15796]='h0000221e;
    rd_cycle[15797] = 1'b1;  wr_cycle[15797] = 1'b0;  addr_rom[15797]='h000001a4;  wr_data_rom[15797]='h00000000;
    rd_cycle[15798] = 1'b1;  wr_cycle[15798] = 1'b0;  addr_rom[15798]='h00003144;  wr_data_rom[15798]='h00000000;
    rd_cycle[15799] = 1'b0;  wr_cycle[15799] = 1'b1;  addr_rom[15799]='h000028c4;  wr_data_rom[15799]='h000024f0;
    rd_cycle[15800] = 1'b0;  wr_cycle[15800] = 1'b1;  addr_rom[15800]='h00001dc4;  wr_data_rom[15800]='h00002ff9;
    rd_cycle[15801] = 1'b0;  wr_cycle[15801] = 1'b1;  addr_rom[15801]='h00003670;  wr_data_rom[15801]='h0000071d;
    rd_cycle[15802] = 1'b0;  wr_cycle[15802] = 1'b1;  addr_rom[15802]='h00002aec;  wr_data_rom[15802]='h00000c36;
    rd_cycle[15803] = 1'b0;  wr_cycle[15803] = 1'b1;  addr_rom[15803]='h000025c4;  wr_data_rom[15803]='h00003c0c;
    rd_cycle[15804] = 1'b1;  wr_cycle[15804] = 1'b0;  addr_rom[15804]='h00000b48;  wr_data_rom[15804]='h00000000;
    rd_cycle[15805] = 1'b0;  wr_cycle[15805] = 1'b1;  addr_rom[15805]='h00000c1c;  wr_data_rom[15805]='h00002649;
    rd_cycle[15806] = 1'b1;  wr_cycle[15806] = 1'b0;  addr_rom[15806]='h00003a50;  wr_data_rom[15806]='h00000000;
    rd_cycle[15807] = 1'b1;  wr_cycle[15807] = 1'b0;  addr_rom[15807]='h000038d4;  wr_data_rom[15807]='h00000000;
    rd_cycle[15808] = 1'b0;  wr_cycle[15808] = 1'b1;  addr_rom[15808]='h00001b74;  wr_data_rom[15808]='h000002ac;
    rd_cycle[15809] = 1'b1;  wr_cycle[15809] = 1'b0;  addr_rom[15809]='h00000e24;  wr_data_rom[15809]='h00000000;
    rd_cycle[15810] = 1'b1;  wr_cycle[15810] = 1'b0;  addr_rom[15810]='h0000154c;  wr_data_rom[15810]='h00000000;
    rd_cycle[15811] = 1'b1;  wr_cycle[15811] = 1'b0;  addr_rom[15811]='h0000151c;  wr_data_rom[15811]='h00000000;
    rd_cycle[15812] = 1'b1;  wr_cycle[15812] = 1'b0;  addr_rom[15812]='h00002978;  wr_data_rom[15812]='h00000000;
    rd_cycle[15813] = 1'b0;  wr_cycle[15813] = 1'b1;  addr_rom[15813]='h00002b04;  wr_data_rom[15813]='h00000cca;
    rd_cycle[15814] = 1'b1;  wr_cycle[15814] = 1'b0;  addr_rom[15814]='h00003050;  wr_data_rom[15814]='h00000000;
    rd_cycle[15815] = 1'b1;  wr_cycle[15815] = 1'b0;  addr_rom[15815]='h00002c1c;  wr_data_rom[15815]='h00000000;
    rd_cycle[15816] = 1'b1;  wr_cycle[15816] = 1'b0;  addr_rom[15816]='h0000359c;  wr_data_rom[15816]='h00000000;
    rd_cycle[15817] = 1'b1;  wr_cycle[15817] = 1'b0;  addr_rom[15817]='h000025ec;  wr_data_rom[15817]='h00000000;
    rd_cycle[15818] = 1'b1;  wr_cycle[15818] = 1'b0;  addr_rom[15818]='h00003adc;  wr_data_rom[15818]='h00000000;
    rd_cycle[15819] = 1'b0;  wr_cycle[15819] = 1'b1;  addr_rom[15819]='h00001040;  wr_data_rom[15819]='h000007db;
    rd_cycle[15820] = 1'b1;  wr_cycle[15820] = 1'b0;  addr_rom[15820]='h00001220;  wr_data_rom[15820]='h00000000;
    rd_cycle[15821] = 1'b1;  wr_cycle[15821] = 1'b0;  addr_rom[15821]='h0000074c;  wr_data_rom[15821]='h00000000;
    rd_cycle[15822] = 1'b0;  wr_cycle[15822] = 1'b1;  addr_rom[15822]='h000012b8;  wr_data_rom[15822]='h000027e0;
    rd_cycle[15823] = 1'b1;  wr_cycle[15823] = 1'b0;  addr_rom[15823]='h00000980;  wr_data_rom[15823]='h00000000;
    rd_cycle[15824] = 1'b0;  wr_cycle[15824] = 1'b1;  addr_rom[15824]='h000004cc;  wr_data_rom[15824]='h00002191;
    rd_cycle[15825] = 1'b1;  wr_cycle[15825] = 1'b0;  addr_rom[15825]='h00000050;  wr_data_rom[15825]='h00000000;
    rd_cycle[15826] = 1'b0;  wr_cycle[15826] = 1'b1;  addr_rom[15826]='h000013a0;  wr_data_rom[15826]='h0000257c;
    rd_cycle[15827] = 1'b1;  wr_cycle[15827] = 1'b0;  addr_rom[15827]='h00003e40;  wr_data_rom[15827]='h00000000;
    rd_cycle[15828] = 1'b0;  wr_cycle[15828] = 1'b1;  addr_rom[15828]='h00001c80;  wr_data_rom[15828]='h00002d9d;
    rd_cycle[15829] = 1'b0;  wr_cycle[15829] = 1'b1;  addr_rom[15829]='h0000046c;  wr_data_rom[15829]='h0000352f;
    rd_cycle[15830] = 1'b1;  wr_cycle[15830] = 1'b0;  addr_rom[15830]='h00001440;  wr_data_rom[15830]='h00000000;
    rd_cycle[15831] = 1'b0;  wr_cycle[15831] = 1'b1;  addr_rom[15831]='h000019d8;  wr_data_rom[15831]='h00000972;
    rd_cycle[15832] = 1'b0;  wr_cycle[15832] = 1'b1;  addr_rom[15832]='h00001ac0;  wr_data_rom[15832]='h000034d5;
    rd_cycle[15833] = 1'b0;  wr_cycle[15833] = 1'b1;  addr_rom[15833]='h00003a80;  wr_data_rom[15833]='h00001394;
    rd_cycle[15834] = 1'b1;  wr_cycle[15834] = 1'b0;  addr_rom[15834]='h00003a38;  wr_data_rom[15834]='h00000000;
    rd_cycle[15835] = 1'b1;  wr_cycle[15835] = 1'b0;  addr_rom[15835]='h000014d0;  wr_data_rom[15835]='h00000000;
    rd_cycle[15836] = 1'b0;  wr_cycle[15836] = 1'b1;  addr_rom[15836]='h00000124;  wr_data_rom[15836]='h000025f9;
    rd_cycle[15837] = 1'b1;  wr_cycle[15837] = 1'b0;  addr_rom[15837]='h000032d0;  wr_data_rom[15837]='h00000000;
    rd_cycle[15838] = 1'b0;  wr_cycle[15838] = 1'b1;  addr_rom[15838]='h000023fc;  wr_data_rom[15838]='h00001228;
    rd_cycle[15839] = 1'b1;  wr_cycle[15839] = 1'b0;  addr_rom[15839]='h000001ec;  wr_data_rom[15839]='h00000000;
    rd_cycle[15840] = 1'b0;  wr_cycle[15840] = 1'b1;  addr_rom[15840]='h000024b8;  wr_data_rom[15840]='h00000188;
    rd_cycle[15841] = 1'b0;  wr_cycle[15841] = 1'b1;  addr_rom[15841]='h00003048;  wr_data_rom[15841]='h000038a7;
    rd_cycle[15842] = 1'b1;  wr_cycle[15842] = 1'b0;  addr_rom[15842]='h000007cc;  wr_data_rom[15842]='h00000000;
    rd_cycle[15843] = 1'b1;  wr_cycle[15843] = 1'b0;  addr_rom[15843]='h000009c4;  wr_data_rom[15843]='h00000000;
    rd_cycle[15844] = 1'b1;  wr_cycle[15844] = 1'b0;  addr_rom[15844]='h00001c20;  wr_data_rom[15844]='h00000000;
    rd_cycle[15845] = 1'b0;  wr_cycle[15845] = 1'b1;  addr_rom[15845]='h000002bc;  wr_data_rom[15845]='h00000c3f;
    rd_cycle[15846] = 1'b0;  wr_cycle[15846] = 1'b1;  addr_rom[15846]='h00001f00;  wr_data_rom[15846]='h0000212c;
    rd_cycle[15847] = 1'b1;  wr_cycle[15847] = 1'b0;  addr_rom[15847]='h00002264;  wr_data_rom[15847]='h00000000;
    rd_cycle[15848] = 1'b0;  wr_cycle[15848] = 1'b1;  addr_rom[15848]='h00001a20;  wr_data_rom[15848]='h000002f1;
    rd_cycle[15849] = 1'b1;  wr_cycle[15849] = 1'b0;  addr_rom[15849]='h000009f0;  wr_data_rom[15849]='h00000000;
    rd_cycle[15850] = 1'b0;  wr_cycle[15850] = 1'b1;  addr_rom[15850]='h00000fc4;  wr_data_rom[15850]='h00003584;
    rd_cycle[15851] = 1'b0;  wr_cycle[15851] = 1'b1;  addr_rom[15851]='h00003dc0;  wr_data_rom[15851]='h0000147c;
    rd_cycle[15852] = 1'b0;  wr_cycle[15852] = 1'b1;  addr_rom[15852]='h00003414;  wr_data_rom[15852]='h000007d9;
    rd_cycle[15853] = 1'b0;  wr_cycle[15853] = 1'b1;  addr_rom[15853]='h00000208;  wr_data_rom[15853]='h00003359;
    rd_cycle[15854] = 1'b0;  wr_cycle[15854] = 1'b1;  addr_rom[15854]='h000034e4;  wr_data_rom[15854]='h00002bf3;
    rd_cycle[15855] = 1'b1;  wr_cycle[15855] = 1'b0;  addr_rom[15855]='h000006a0;  wr_data_rom[15855]='h00000000;
    rd_cycle[15856] = 1'b0;  wr_cycle[15856] = 1'b1;  addr_rom[15856]='h00001c08;  wr_data_rom[15856]='h00000def;
    rd_cycle[15857] = 1'b1;  wr_cycle[15857] = 1'b0;  addr_rom[15857]='h00002dd0;  wr_data_rom[15857]='h00000000;
    rd_cycle[15858] = 1'b0;  wr_cycle[15858] = 1'b1;  addr_rom[15858]='h00000bb8;  wr_data_rom[15858]='h00002c6d;
    rd_cycle[15859] = 1'b1;  wr_cycle[15859] = 1'b0;  addr_rom[15859]='h000001dc;  wr_data_rom[15859]='h00000000;
    rd_cycle[15860] = 1'b1;  wr_cycle[15860] = 1'b0;  addr_rom[15860]='h00003094;  wr_data_rom[15860]='h00000000;
    rd_cycle[15861] = 1'b0;  wr_cycle[15861] = 1'b1;  addr_rom[15861]='h00003df0;  wr_data_rom[15861]='h0000059e;
    rd_cycle[15862] = 1'b0;  wr_cycle[15862] = 1'b1;  addr_rom[15862]='h000000a4;  wr_data_rom[15862]='h00003bf8;
    rd_cycle[15863] = 1'b1;  wr_cycle[15863] = 1'b0;  addr_rom[15863]='h000000a8;  wr_data_rom[15863]='h00000000;
    rd_cycle[15864] = 1'b1;  wr_cycle[15864] = 1'b0;  addr_rom[15864]='h0000004c;  wr_data_rom[15864]='h00000000;
    rd_cycle[15865] = 1'b1;  wr_cycle[15865] = 1'b0;  addr_rom[15865]='h0000248c;  wr_data_rom[15865]='h00000000;
    rd_cycle[15866] = 1'b0;  wr_cycle[15866] = 1'b1;  addr_rom[15866]='h000038ac;  wr_data_rom[15866]='h00000237;
    rd_cycle[15867] = 1'b1;  wr_cycle[15867] = 1'b0;  addr_rom[15867]='h00003c40;  wr_data_rom[15867]='h00000000;
    rd_cycle[15868] = 1'b0;  wr_cycle[15868] = 1'b1;  addr_rom[15868]='h0000331c;  wr_data_rom[15868]='h00002dd5;
    rd_cycle[15869] = 1'b1;  wr_cycle[15869] = 1'b0;  addr_rom[15869]='h000031b8;  wr_data_rom[15869]='h00000000;
    rd_cycle[15870] = 1'b0;  wr_cycle[15870] = 1'b1;  addr_rom[15870]='h00003cac;  wr_data_rom[15870]='h0000176f;
    rd_cycle[15871] = 1'b1;  wr_cycle[15871] = 1'b0;  addr_rom[15871]='h000036dc;  wr_data_rom[15871]='h00000000;
    rd_cycle[15872] = 1'b0;  wr_cycle[15872] = 1'b1;  addr_rom[15872]='h0000031c;  wr_data_rom[15872]='h0000252d;
    rd_cycle[15873] = 1'b1;  wr_cycle[15873] = 1'b0;  addr_rom[15873]='h000037e8;  wr_data_rom[15873]='h00000000;
    rd_cycle[15874] = 1'b1;  wr_cycle[15874] = 1'b0;  addr_rom[15874]='h00003f70;  wr_data_rom[15874]='h00000000;
    rd_cycle[15875] = 1'b0;  wr_cycle[15875] = 1'b1;  addr_rom[15875]='h00002ed8;  wr_data_rom[15875]='h00002219;
    rd_cycle[15876] = 1'b0;  wr_cycle[15876] = 1'b1;  addr_rom[15876]='h00001f3c;  wr_data_rom[15876]='h00003296;
    rd_cycle[15877] = 1'b0;  wr_cycle[15877] = 1'b1;  addr_rom[15877]='h000016ac;  wr_data_rom[15877]='h00002144;
    rd_cycle[15878] = 1'b0;  wr_cycle[15878] = 1'b1;  addr_rom[15878]='h00001d74;  wr_data_rom[15878]='h000022bc;
    rd_cycle[15879] = 1'b0;  wr_cycle[15879] = 1'b1;  addr_rom[15879]='h000034e8;  wr_data_rom[15879]='h00001216;
    rd_cycle[15880] = 1'b0;  wr_cycle[15880] = 1'b1;  addr_rom[15880]='h0000193c;  wr_data_rom[15880]='h00003989;
    rd_cycle[15881] = 1'b0;  wr_cycle[15881] = 1'b1;  addr_rom[15881]='h00000750;  wr_data_rom[15881]='h00001ae0;
    rd_cycle[15882] = 1'b1;  wr_cycle[15882] = 1'b0;  addr_rom[15882]='h00002260;  wr_data_rom[15882]='h00000000;
    rd_cycle[15883] = 1'b1;  wr_cycle[15883] = 1'b0;  addr_rom[15883]='h00001f98;  wr_data_rom[15883]='h00000000;
    rd_cycle[15884] = 1'b1;  wr_cycle[15884] = 1'b0;  addr_rom[15884]='h00000bec;  wr_data_rom[15884]='h00000000;
    rd_cycle[15885] = 1'b1;  wr_cycle[15885] = 1'b0;  addr_rom[15885]='h00003ae8;  wr_data_rom[15885]='h00000000;
    rd_cycle[15886] = 1'b1;  wr_cycle[15886] = 1'b0;  addr_rom[15886]='h00001f90;  wr_data_rom[15886]='h00000000;
    rd_cycle[15887] = 1'b0;  wr_cycle[15887] = 1'b1;  addr_rom[15887]='h00003b94;  wr_data_rom[15887]='h00003c86;
    rd_cycle[15888] = 1'b1;  wr_cycle[15888] = 1'b0;  addr_rom[15888]='h000025e0;  wr_data_rom[15888]='h00000000;
    rd_cycle[15889] = 1'b1;  wr_cycle[15889] = 1'b0;  addr_rom[15889]='h000009c8;  wr_data_rom[15889]='h00000000;
    rd_cycle[15890] = 1'b0;  wr_cycle[15890] = 1'b1;  addr_rom[15890]='h0000248c;  wr_data_rom[15890]='h00002e2f;
    rd_cycle[15891] = 1'b0;  wr_cycle[15891] = 1'b1;  addr_rom[15891]='h00001488;  wr_data_rom[15891]='h00003d52;
    rd_cycle[15892] = 1'b0;  wr_cycle[15892] = 1'b1;  addr_rom[15892]='h00001b14;  wr_data_rom[15892]='h0000324d;
    rd_cycle[15893] = 1'b1;  wr_cycle[15893] = 1'b0;  addr_rom[15893]='h000002b4;  wr_data_rom[15893]='h00000000;
    rd_cycle[15894] = 1'b0;  wr_cycle[15894] = 1'b1;  addr_rom[15894]='h00000a1c;  wr_data_rom[15894]='h00001f58;
    rd_cycle[15895] = 1'b1;  wr_cycle[15895] = 1'b0;  addr_rom[15895]='h00001d94;  wr_data_rom[15895]='h00000000;
    rd_cycle[15896] = 1'b1;  wr_cycle[15896] = 1'b0;  addr_rom[15896]='h0000130c;  wr_data_rom[15896]='h00000000;
    rd_cycle[15897] = 1'b1;  wr_cycle[15897] = 1'b0;  addr_rom[15897]='h00002f1c;  wr_data_rom[15897]='h00000000;
    rd_cycle[15898] = 1'b1;  wr_cycle[15898] = 1'b0;  addr_rom[15898]='h0000190c;  wr_data_rom[15898]='h00000000;
    rd_cycle[15899] = 1'b0;  wr_cycle[15899] = 1'b1;  addr_rom[15899]='h00000640;  wr_data_rom[15899]='h00002149;
    rd_cycle[15900] = 1'b0;  wr_cycle[15900] = 1'b1;  addr_rom[15900]='h000026e0;  wr_data_rom[15900]='h000010d4;
    rd_cycle[15901] = 1'b0;  wr_cycle[15901] = 1'b1;  addr_rom[15901]='h00002e54;  wr_data_rom[15901]='h00002f50;
    rd_cycle[15902] = 1'b1;  wr_cycle[15902] = 1'b0;  addr_rom[15902]='h000010c8;  wr_data_rom[15902]='h00000000;
    rd_cycle[15903] = 1'b1;  wr_cycle[15903] = 1'b0;  addr_rom[15903]='h000014dc;  wr_data_rom[15903]='h00000000;
    rd_cycle[15904] = 1'b0;  wr_cycle[15904] = 1'b1;  addr_rom[15904]='h000022f4;  wr_data_rom[15904]='h00000597;
    rd_cycle[15905] = 1'b1;  wr_cycle[15905] = 1'b0;  addr_rom[15905]='h000031d4;  wr_data_rom[15905]='h00000000;
    rd_cycle[15906] = 1'b0;  wr_cycle[15906] = 1'b1;  addr_rom[15906]='h0000024c;  wr_data_rom[15906]='h00003f82;
    rd_cycle[15907] = 1'b1;  wr_cycle[15907] = 1'b0;  addr_rom[15907]='h00001360;  wr_data_rom[15907]='h00000000;
    rd_cycle[15908] = 1'b1;  wr_cycle[15908] = 1'b0;  addr_rom[15908]='h00000f58;  wr_data_rom[15908]='h00000000;
    rd_cycle[15909] = 1'b1;  wr_cycle[15909] = 1'b0;  addr_rom[15909]='h00000cdc;  wr_data_rom[15909]='h00000000;
    rd_cycle[15910] = 1'b1;  wr_cycle[15910] = 1'b0;  addr_rom[15910]='h00003474;  wr_data_rom[15910]='h00000000;
    rd_cycle[15911] = 1'b0;  wr_cycle[15911] = 1'b1;  addr_rom[15911]='h00001650;  wr_data_rom[15911]='h00002b0e;
    rd_cycle[15912] = 1'b0;  wr_cycle[15912] = 1'b1;  addr_rom[15912]='h00000f68;  wr_data_rom[15912]='h00003a2d;
    rd_cycle[15913] = 1'b1;  wr_cycle[15913] = 1'b0;  addr_rom[15913]='h00002914;  wr_data_rom[15913]='h00000000;
    rd_cycle[15914] = 1'b0;  wr_cycle[15914] = 1'b1;  addr_rom[15914]='h00001714;  wr_data_rom[15914]='h00002abc;
    rd_cycle[15915] = 1'b0;  wr_cycle[15915] = 1'b1;  addr_rom[15915]='h0000033c;  wr_data_rom[15915]='h00002d5d;
    rd_cycle[15916] = 1'b0;  wr_cycle[15916] = 1'b1;  addr_rom[15916]='h00002c80;  wr_data_rom[15916]='h00000196;
    rd_cycle[15917] = 1'b1;  wr_cycle[15917] = 1'b0;  addr_rom[15917]='h00001a74;  wr_data_rom[15917]='h00000000;
    rd_cycle[15918] = 1'b0;  wr_cycle[15918] = 1'b1;  addr_rom[15918]='h000000dc;  wr_data_rom[15918]='h00000ee1;
    rd_cycle[15919] = 1'b1;  wr_cycle[15919] = 1'b0;  addr_rom[15919]='h000026f4;  wr_data_rom[15919]='h00000000;
    rd_cycle[15920] = 1'b1;  wr_cycle[15920] = 1'b0;  addr_rom[15920]='h00000a70;  wr_data_rom[15920]='h00000000;
    rd_cycle[15921] = 1'b0;  wr_cycle[15921] = 1'b1;  addr_rom[15921]='h000005f8;  wr_data_rom[15921]='h00001785;
    rd_cycle[15922] = 1'b0;  wr_cycle[15922] = 1'b1;  addr_rom[15922]='h00003a10;  wr_data_rom[15922]='h000031d0;
    rd_cycle[15923] = 1'b0;  wr_cycle[15923] = 1'b1;  addr_rom[15923]='h00003ad0;  wr_data_rom[15923]='h00002196;
    rd_cycle[15924] = 1'b0;  wr_cycle[15924] = 1'b1;  addr_rom[15924]='h00003a24;  wr_data_rom[15924]='h00002480;
    rd_cycle[15925] = 1'b1;  wr_cycle[15925] = 1'b0;  addr_rom[15925]='h000001a8;  wr_data_rom[15925]='h00000000;
    rd_cycle[15926] = 1'b0;  wr_cycle[15926] = 1'b1;  addr_rom[15926]='h00003b68;  wr_data_rom[15926]='h0000165d;
    rd_cycle[15927] = 1'b1;  wr_cycle[15927] = 1'b0;  addr_rom[15927]='h00002930;  wr_data_rom[15927]='h00000000;
    rd_cycle[15928] = 1'b0;  wr_cycle[15928] = 1'b1;  addr_rom[15928]='h00001474;  wr_data_rom[15928]='h00002f15;
    rd_cycle[15929] = 1'b0;  wr_cycle[15929] = 1'b1;  addr_rom[15929]='h00002104;  wr_data_rom[15929]='h000013be;
    rd_cycle[15930] = 1'b1;  wr_cycle[15930] = 1'b0;  addr_rom[15930]='h00001414;  wr_data_rom[15930]='h00000000;
    rd_cycle[15931] = 1'b1;  wr_cycle[15931] = 1'b0;  addr_rom[15931]='h00001f80;  wr_data_rom[15931]='h00000000;
    rd_cycle[15932] = 1'b0;  wr_cycle[15932] = 1'b1;  addr_rom[15932]='h000020d8;  wr_data_rom[15932]='h00000ec1;
    rd_cycle[15933] = 1'b0;  wr_cycle[15933] = 1'b1;  addr_rom[15933]='h00003c2c;  wr_data_rom[15933]='h00002912;
    rd_cycle[15934] = 1'b0;  wr_cycle[15934] = 1'b1;  addr_rom[15934]='h00003ac8;  wr_data_rom[15934]='h000016d3;
    rd_cycle[15935] = 1'b0;  wr_cycle[15935] = 1'b1;  addr_rom[15935]='h000018d4;  wr_data_rom[15935]='h000020f1;
    rd_cycle[15936] = 1'b0;  wr_cycle[15936] = 1'b1;  addr_rom[15936]='h00002ba4;  wr_data_rom[15936]='h00001383;
    rd_cycle[15937] = 1'b0;  wr_cycle[15937] = 1'b1;  addr_rom[15937]='h00001504;  wr_data_rom[15937]='h00003bcf;
    rd_cycle[15938] = 1'b0;  wr_cycle[15938] = 1'b1;  addr_rom[15938]='h00001be8;  wr_data_rom[15938]='h00000625;
    rd_cycle[15939] = 1'b1;  wr_cycle[15939] = 1'b0;  addr_rom[15939]='h0000322c;  wr_data_rom[15939]='h00000000;
    rd_cycle[15940] = 1'b1;  wr_cycle[15940] = 1'b0;  addr_rom[15940]='h00003380;  wr_data_rom[15940]='h00000000;
    rd_cycle[15941] = 1'b1;  wr_cycle[15941] = 1'b0;  addr_rom[15941]='h00002224;  wr_data_rom[15941]='h00000000;
    rd_cycle[15942] = 1'b0;  wr_cycle[15942] = 1'b1;  addr_rom[15942]='h00002ae0;  wr_data_rom[15942]='h00001ab8;
    rd_cycle[15943] = 1'b1;  wr_cycle[15943] = 1'b0;  addr_rom[15943]='h00000b68;  wr_data_rom[15943]='h00000000;
    rd_cycle[15944] = 1'b1;  wr_cycle[15944] = 1'b0;  addr_rom[15944]='h00000b40;  wr_data_rom[15944]='h00000000;
    rd_cycle[15945] = 1'b1;  wr_cycle[15945] = 1'b0;  addr_rom[15945]='h000015ec;  wr_data_rom[15945]='h00000000;
    rd_cycle[15946] = 1'b1;  wr_cycle[15946] = 1'b0;  addr_rom[15946]='h00001358;  wr_data_rom[15946]='h00000000;
    rd_cycle[15947] = 1'b1;  wr_cycle[15947] = 1'b0;  addr_rom[15947]='h00001a30;  wr_data_rom[15947]='h00000000;
    rd_cycle[15948] = 1'b1;  wr_cycle[15948] = 1'b0;  addr_rom[15948]='h00000b08;  wr_data_rom[15948]='h00000000;
    rd_cycle[15949] = 1'b0;  wr_cycle[15949] = 1'b1;  addr_rom[15949]='h0000334c;  wr_data_rom[15949]='h000037de;
    rd_cycle[15950] = 1'b0;  wr_cycle[15950] = 1'b1;  addr_rom[15950]='h00001a2c;  wr_data_rom[15950]='h00001724;
    rd_cycle[15951] = 1'b1;  wr_cycle[15951] = 1'b0;  addr_rom[15951]='h00002e70;  wr_data_rom[15951]='h00000000;
    rd_cycle[15952] = 1'b0;  wr_cycle[15952] = 1'b1;  addr_rom[15952]='h00001c64;  wr_data_rom[15952]='h0000367c;
    rd_cycle[15953] = 1'b0;  wr_cycle[15953] = 1'b1;  addr_rom[15953]='h000038ec;  wr_data_rom[15953]='h00002d00;
    rd_cycle[15954] = 1'b0;  wr_cycle[15954] = 1'b1;  addr_rom[15954]='h00002fe4;  wr_data_rom[15954]='h0000221e;
    rd_cycle[15955] = 1'b0;  wr_cycle[15955] = 1'b1;  addr_rom[15955]='h000017cc;  wr_data_rom[15955]='h00001cae;
    rd_cycle[15956] = 1'b0;  wr_cycle[15956] = 1'b1;  addr_rom[15956]='h000031a8;  wr_data_rom[15956]='h000039c8;
    rd_cycle[15957] = 1'b1;  wr_cycle[15957] = 1'b0;  addr_rom[15957]='h000015c4;  wr_data_rom[15957]='h00000000;
    rd_cycle[15958] = 1'b0;  wr_cycle[15958] = 1'b1;  addr_rom[15958]='h00003b58;  wr_data_rom[15958]='h00001e12;
    rd_cycle[15959] = 1'b0;  wr_cycle[15959] = 1'b1;  addr_rom[15959]='h00000068;  wr_data_rom[15959]='h00001ae3;
    rd_cycle[15960] = 1'b1;  wr_cycle[15960] = 1'b0;  addr_rom[15960]='h0000186c;  wr_data_rom[15960]='h00000000;
    rd_cycle[15961] = 1'b0;  wr_cycle[15961] = 1'b1;  addr_rom[15961]='h0000070c;  wr_data_rom[15961]='h000008a3;
    rd_cycle[15962] = 1'b0;  wr_cycle[15962] = 1'b1;  addr_rom[15962]='h00003d4c;  wr_data_rom[15962]='h00001d52;
    rd_cycle[15963] = 1'b0;  wr_cycle[15963] = 1'b1;  addr_rom[15963]='h00001d14;  wr_data_rom[15963]='h00003678;
    rd_cycle[15964] = 1'b1;  wr_cycle[15964] = 1'b0;  addr_rom[15964]='h00002d7c;  wr_data_rom[15964]='h00000000;
    rd_cycle[15965] = 1'b0;  wr_cycle[15965] = 1'b1;  addr_rom[15965]='h00000864;  wr_data_rom[15965]='h000000bb;
    rd_cycle[15966] = 1'b0;  wr_cycle[15966] = 1'b1;  addr_rom[15966]='h00001d3c;  wr_data_rom[15966]='h00002912;
    rd_cycle[15967] = 1'b0;  wr_cycle[15967] = 1'b1;  addr_rom[15967]='h00000330;  wr_data_rom[15967]='h0000373b;
    rd_cycle[15968] = 1'b1;  wr_cycle[15968] = 1'b0;  addr_rom[15968]='h00000214;  wr_data_rom[15968]='h00000000;
    rd_cycle[15969] = 1'b1;  wr_cycle[15969] = 1'b0;  addr_rom[15969]='h000024c0;  wr_data_rom[15969]='h00000000;
    rd_cycle[15970] = 1'b0;  wr_cycle[15970] = 1'b1;  addr_rom[15970]='h00002784;  wr_data_rom[15970]='h000022d0;
    rd_cycle[15971] = 1'b1;  wr_cycle[15971] = 1'b0;  addr_rom[15971]='h000028ec;  wr_data_rom[15971]='h00000000;
    rd_cycle[15972] = 1'b1;  wr_cycle[15972] = 1'b0;  addr_rom[15972]='h00001d50;  wr_data_rom[15972]='h00000000;
    rd_cycle[15973] = 1'b0;  wr_cycle[15973] = 1'b1;  addr_rom[15973]='h00000ac4;  wr_data_rom[15973]='h0000292b;
    rd_cycle[15974] = 1'b0;  wr_cycle[15974] = 1'b1;  addr_rom[15974]='h000022ac;  wr_data_rom[15974]='h00003fd4;
    rd_cycle[15975] = 1'b1;  wr_cycle[15975] = 1'b0;  addr_rom[15975]='h0000244c;  wr_data_rom[15975]='h00000000;
    rd_cycle[15976] = 1'b0;  wr_cycle[15976] = 1'b1;  addr_rom[15976]='h000038b4;  wr_data_rom[15976]='h00000f45;
    rd_cycle[15977] = 1'b0;  wr_cycle[15977] = 1'b1;  addr_rom[15977]='h00003b70;  wr_data_rom[15977]='h00000a58;
    rd_cycle[15978] = 1'b1;  wr_cycle[15978] = 1'b0;  addr_rom[15978]='h00003f3c;  wr_data_rom[15978]='h00000000;
    rd_cycle[15979] = 1'b0;  wr_cycle[15979] = 1'b1;  addr_rom[15979]='h00000084;  wr_data_rom[15979]='h00002cb6;
    rd_cycle[15980] = 1'b0;  wr_cycle[15980] = 1'b1;  addr_rom[15980]='h00002984;  wr_data_rom[15980]='h0000384f;
    rd_cycle[15981] = 1'b1;  wr_cycle[15981] = 1'b0;  addr_rom[15981]='h00000448;  wr_data_rom[15981]='h00000000;
    rd_cycle[15982] = 1'b0;  wr_cycle[15982] = 1'b1;  addr_rom[15982]='h00002db4;  wr_data_rom[15982]='h00002bc6;
    rd_cycle[15983] = 1'b0;  wr_cycle[15983] = 1'b1;  addr_rom[15983]='h00000c40;  wr_data_rom[15983]='h000013f2;
    rd_cycle[15984] = 1'b1;  wr_cycle[15984] = 1'b0;  addr_rom[15984]='h00003ee4;  wr_data_rom[15984]='h00000000;
    rd_cycle[15985] = 1'b1;  wr_cycle[15985] = 1'b0;  addr_rom[15985]='h00001504;  wr_data_rom[15985]='h00000000;
    rd_cycle[15986] = 1'b1;  wr_cycle[15986] = 1'b0;  addr_rom[15986]='h00001678;  wr_data_rom[15986]='h00000000;
    rd_cycle[15987] = 1'b1;  wr_cycle[15987] = 1'b0;  addr_rom[15987]='h00002f58;  wr_data_rom[15987]='h00000000;
    rd_cycle[15988] = 1'b1;  wr_cycle[15988] = 1'b0;  addr_rom[15988]='h000019a8;  wr_data_rom[15988]='h00000000;
    rd_cycle[15989] = 1'b1;  wr_cycle[15989] = 1'b0;  addr_rom[15989]='h000010b8;  wr_data_rom[15989]='h00000000;
    rd_cycle[15990] = 1'b1;  wr_cycle[15990] = 1'b0;  addr_rom[15990]='h00002ae0;  wr_data_rom[15990]='h00000000;
    rd_cycle[15991] = 1'b1;  wr_cycle[15991] = 1'b0;  addr_rom[15991]='h000002a0;  wr_data_rom[15991]='h00000000;
    rd_cycle[15992] = 1'b1;  wr_cycle[15992] = 1'b0;  addr_rom[15992]='h000036b0;  wr_data_rom[15992]='h00000000;
    rd_cycle[15993] = 1'b1;  wr_cycle[15993] = 1'b0;  addr_rom[15993]='h00003edc;  wr_data_rom[15993]='h00000000;
    rd_cycle[15994] = 1'b0;  wr_cycle[15994] = 1'b1;  addr_rom[15994]='h00000284;  wr_data_rom[15994]='h00001485;
    rd_cycle[15995] = 1'b1;  wr_cycle[15995] = 1'b0;  addr_rom[15995]='h00002a18;  wr_data_rom[15995]='h00000000;
    rd_cycle[15996] = 1'b1;  wr_cycle[15996] = 1'b0;  addr_rom[15996]='h0000155c;  wr_data_rom[15996]='h00000000;
    rd_cycle[15997] = 1'b0;  wr_cycle[15997] = 1'b1;  addr_rom[15997]='h000010b4;  wr_data_rom[15997]='h00001c21;
    rd_cycle[15998] = 1'b0;  wr_cycle[15998] = 1'b1;  addr_rom[15998]='h00003380;  wr_data_rom[15998]='h000037b9;
    rd_cycle[15999] = 1'b1;  wr_cycle[15999] = 1'b0;  addr_rom[15999]='h00003974;  wr_data_rom[15999]='h00000000;
    rd_cycle[16000] = 1'b1;  wr_cycle[16000] = 1'b0;  addr_rom[16000]='h000014bc;  wr_data_rom[16000]='h00000000;
    rd_cycle[16001] = 1'b1;  wr_cycle[16001] = 1'b0;  addr_rom[16001]='h00002bc0;  wr_data_rom[16001]='h00000000;
    rd_cycle[16002] = 1'b0;  wr_cycle[16002] = 1'b1;  addr_rom[16002]='h00002b0c;  wr_data_rom[16002]='h00001e55;
    rd_cycle[16003] = 1'b0;  wr_cycle[16003] = 1'b1;  addr_rom[16003]='h00002758;  wr_data_rom[16003]='h000022ee;
    rd_cycle[16004] = 1'b0;  wr_cycle[16004] = 1'b1;  addr_rom[16004]='h0000080c;  wr_data_rom[16004]='h000032f8;
    rd_cycle[16005] = 1'b1;  wr_cycle[16005] = 1'b0;  addr_rom[16005]='h00003e44;  wr_data_rom[16005]='h00000000;
    rd_cycle[16006] = 1'b1;  wr_cycle[16006] = 1'b0;  addr_rom[16006]='h000031c0;  wr_data_rom[16006]='h00000000;
    rd_cycle[16007] = 1'b0;  wr_cycle[16007] = 1'b1;  addr_rom[16007]='h00000008;  wr_data_rom[16007]='h000020d5;
    rd_cycle[16008] = 1'b0;  wr_cycle[16008] = 1'b1;  addr_rom[16008]='h00001eb4;  wr_data_rom[16008]='h00002f1c;
    rd_cycle[16009] = 1'b1;  wr_cycle[16009] = 1'b0;  addr_rom[16009]='h00001264;  wr_data_rom[16009]='h00000000;
    rd_cycle[16010] = 1'b0;  wr_cycle[16010] = 1'b1;  addr_rom[16010]='h00001e74;  wr_data_rom[16010]='h00001f55;
    rd_cycle[16011] = 1'b0;  wr_cycle[16011] = 1'b1;  addr_rom[16011]='h00000a84;  wr_data_rom[16011]='h0000193c;
    rd_cycle[16012] = 1'b0;  wr_cycle[16012] = 1'b1;  addr_rom[16012]='h00003128;  wr_data_rom[16012]='h00003aae;
    rd_cycle[16013] = 1'b0;  wr_cycle[16013] = 1'b1;  addr_rom[16013]='h0000024c;  wr_data_rom[16013]='h000000e3;
    rd_cycle[16014] = 1'b1;  wr_cycle[16014] = 1'b0;  addr_rom[16014]='h00000658;  wr_data_rom[16014]='h00000000;
    rd_cycle[16015] = 1'b0;  wr_cycle[16015] = 1'b1;  addr_rom[16015]='h00001350;  wr_data_rom[16015]='h00000aba;
    rd_cycle[16016] = 1'b1;  wr_cycle[16016] = 1'b0;  addr_rom[16016]='h00001b88;  wr_data_rom[16016]='h00000000;
    rd_cycle[16017] = 1'b1;  wr_cycle[16017] = 1'b0;  addr_rom[16017]='h00001b00;  wr_data_rom[16017]='h00000000;
    rd_cycle[16018] = 1'b0;  wr_cycle[16018] = 1'b1;  addr_rom[16018]='h00002610;  wr_data_rom[16018]='h000038f3;
    rd_cycle[16019] = 1'b1;  wr_cycle[16019] = 1'b0;  addr_rom[16019]='h00000190;  wr_data_rom[16019]='h00000000;
    rd_cycle[16020] = 1'b0;  wr_cycle[16020] = 1'b1;  addr_rom[16020]='h00002fa0;  wr_data_rom[16020]='h000012d4;
    rd_cycle[16021] = 1'b0;  wr_cycle[16021] = 1'b1;  addr_rom[16021]='h00000670;  wr_data_rom[16021]='h00000ea1;
    rd_cycle[16022] = 1'b1;  wr_cycle[16022] = 1'b0;  addr_rom[16022]='h0000129c;  wr_data_rom[16022]='h00000000;
    rd_cycle[16023] = 1'b1;  wr_cycle[16023] = 1'b0;  addr_rom[16023]='h00003798;  wr_data_rom[16023]='h00000000;
    rd_cycle[16024] = 1'b1;  wr_cycle[16024] = 1'b0;  addr_rom[16024]='h00002614;  wr_data_rom[16024]='h00000000;
    rd_cycle[16025] = 1'b0;  wr_cycle[16025] = 1'b1;  addr_rom[16025]='h000001e8;  wr_data_rom[16025]='h00000cf7;
    rd_cycle[16026] = 1'b0;  wr_cycle[16026] = 1'b1;  addr_rom[16026]='h00003a20;  wr_data_rom[16026]='h00002714;
    rd_cycle[16027] = 1'b0;  wr_cycle[16027] = 1'b1;  addr_rom[16027]='h00002f8c;  wr_data_rom[16027]='h00001707;
    rd_cycle[16028] = 1'b1;  wr_cycle[16028] = 1'b0;  addr_rom[16028]='h00003c64;  wr_data_rom[16028]='h00000000;
    rd_cycle[16029] = 1'b1;  wr_cycle[16029] = 1'b0;  addr_rom[16029]='h00001a34;  wr_data_rom[16029]='h00000000;
    rd_cycle[16030] = 1'b0;  wr_cycle[16030] = 1'b1;  addr_rom[16030]='h000027ac;  wr_data_rom[16030]='h000000f8;
    rd_cycle[16031] = 1'b0;  wr_cycle[16031] = 1'b1;  addr_rom[16031]='h00000050;  wr_data_rom[16031]='h00000e19;
    rd_cycle[16032] = 1'b1;  wr_cycle[16032] = 1'b0;  addr_rom[16032]='h00000dd4;  wr_data_rom[16032]='h00000000;
    rd_cycle[16033] = 1'b1;  wr_cycle[16033] = 1'b0;  addr_rom[16033]='h00000c90;  wr_data_rom[16033]='h00000000;
    rd_cycle[16034] = 1'b0;  wr_cycle[16034] = 1'b1;  addr_rom[16034]='h00001f1c;  wr_data_rom[16034]='h00000faa;
    rd_cycle[16035] = 1'b1;  wr_cycle[16035] = 1'b0;  addr_rom[16035]='h0000146c;  wr_data_rom[16035]='h00000000;
    rd_cycle[16036] = 1'b0;  wr_cycle[16036] = 1'b1;  addr_rom[16036]='h0000142c;  wr_data_rom[16036]='h00001c5a;
    rd_cycle[16037] = 1'b1;  wr_cycle[16037] = 1'b0;  addr_rom[16037]='h000014e8;  wr_data_rom[16037]='h00000000;
    rd_cycle[16038] = 1'b1;  wr_cycle[16038] = 1'b0;  addr_rom[16038]='h000010cc;  wr_data_rom[16038]='h00000000;
    rd_cycle[16039] = 1'b0;  wr_cycle[16039] = 1'b1;  addr_rom[16039]='h00000580;  wr_data_rom[16039]='h00001aa8;
    rd_cycle[16040] = 1'b0;  wr_cycle[16040] = 1'b1;  addr_rom[16040]='h000032a4;  wr_data_rom[16040]='h00002178;
    rd_cycle[16041] = 1'b0;  wr_cycle[16041] = 1'b1;  addr_rom[16041]='h000002a4;  wr_data_rom[16041]='h000006fd;
    rd_cycle[16042] = 1'b0;  wr_cycle[16042] = 1'b1;  addr_rom[16042]='h000029e0;  wr_data_rom[16042]='h0000024a;
    rd_cycle[16043] = 1'b1;  wr_cycle[16043] = 1'b0;  addr_rom[16043]='h000007bc;  wr_data_rom[16043]='h00000000;
    rd_cycle[16044] = 1'b0;  wr_cycle[16044] = 1'b1;  addr_rom[16044]='h00001390;  wr_data_rom[16044]='h000036dc;
    rd_cycle[16045] = 1'b1;  wr_cycle[16045] = 1'b0;  addr_rom[16045]='h00002da8;  wr_data_rom[16045]='h00000000;
    rd_cycle[16046] = 1'b0;  wr_cycle[16046] = 1'b1;  addr_rom[16046]='h00000ff0;  wr_data_rom[16046]='h00002b25;
    rd_cycle[16047] = 1'b1;  wr_cycle[16047] = 1'b0;  addr_rom[16047]='h00002e18;  wr_data_rom[16047]='h00000000;
    rd_cycle[16048] = 1'b0;  wr_cycle[16048] = 1'b1;  addr_rom[16048]='h00002940;  wr_data_rom[16048]='h00003250;
    rd_cycle[16049] = 1'b0;  wr_cycle[16049] = 1'b1;  addr_rom[16049]='h000039d0;  wr_data_rom[16049]='h00002813;
    rd_cycle[16050] = 1'b0;  wr_cycle[16050] = 1'b1;  addr_rom[16050]='h00001d4c;  wr_data_rom[16050]='h0000347e;
    rd_cycle[16051] = 1'b1;  wr_cycle[16051] = 1'b0;  addr_rom[16051]='h0000151c;  wr_data_rom[16051]='h00000000;
    rd_cycle[16052] = 1'b1;  wr_cycle[16052] = 1'b0;  addr_rom[16052]='h00003f50;  wr_data_rom[16052]='h00000000;
    rd_cycle[16053] = 1'b1;  wr_cycle[16053] = 1'b0;  addr_rom[16053]='h00000b80;  wr_data_rom[16053]='h00000000;
    rd_cycle[16054] = 1'b1;  wr_cycle[16054] = 1'b0;  addr_rom[16054]='h000005d0;  wr_data_rom[16054]='h00000000;
    rd_cycle[16055] = 1'b0;  wr_cycle[16055] = 1'b1;  addr_rom[16055]='h00002358;  wr_data_rom[16055]='h0000327a;
    rd_cycle[16056] = 1'b0;  wr_cycle[16056] = 1'b1;  addr_rom[16056]='h00000030;  wr_data_rom[16056]='h00001fc2;
    rd_cycle[16057] = 1'b0;  wr_cycle[16057] = 1'b1;  addr_rom[16057]='h000012e4;  wr_data_rom[16057]='h00003cd9;
    rd_cycle[16058] = 1'b0;  wr_cycle[16058] = 1'b1;  addr_rom[16058]='h00000f38;  wr_data_rom[16058]='h00003772;
    rd_cycle[16059] = 1'b0;  wr_cycle[16059] = 1'b1;  addr_rom[16059]='h00001310;  wr_data_rom[16059]='h00000552;
    rd_cycle[16060] = 1'b0;  wr_cycle[16060] = 1'b1;  addr_rom[16060]='h00002c24;  wr_data_rom[16060]='h00001a96;
    rd_cycle[16061] = 1'b1;  wr_cycle[16061] = 1'b0;  addr_rom[16061]='h00001ce4;  wr_data_rom[16061]='h00000000;
    rd_cycle[16062] = 1'b1;  wr_cycle[16062] = 1'b0;  addr_rom[16062]='h000031f0;  wr_data_rom[16062]='h00000000;
    rd_cycle[16063] = 1'b0;  wr_cycle[16063] = 1'b1;  addr_rom[16063]='h00002698;  wr_data_rom[16063]='h000002cf;
    rd_cycle[16064] = 1'b0;  wr_cycle[16064] = 1'b1;  addr_rom[16064]='h00000168;  wr_data_rom[16064]='h00000c7a;
    rd_cycle[16065] = 1'b0;  wr_cycle[16065] = 1'b1;  addr_rom[16065]='h00001774;  wr_data_rom[16065]='h00001bec;
    rd_cycle[16066] = 1'b0;  wr_cycle[16066] = 1'b1;  addr_rom[16066]='h00003ed4;  wr_data_rom[16066]='h00002651;
    rd_cycle[16067] = 1'b0;  wr_cycle[16067] = 1'b1;  addr_rom[16067]='h00003df8;  wr_data_rom[16067]='h00000a9c;
    rd_cycle[16068] = 1'b1;  wr_cycle[16068] = 1'b0;  addr_rom[16068]='h00001860;  wr_data_rom[16068]='h00000000;
    rd_cycle[16069] = 1'b0;  wr_cycle[16069] = 1'b1;  addr_rom[16069]='h0000112c;  wr_data_rom[16069]='h0000170c;
    rd_cycle[16070] = 1'b1;  wr_cycle[16070] = 1'b0;  addr_rom[16070]='h000011c4;  wr_data_rom[16070]='h00000000;
    rd_cycle[16071] = 1'b1;  wr_cycle[16071] = 1'b0;  addr_rom[16071]='h0000105c;  wr_data_rom[16071]='h00000000;
    rd_cycle[16072] = 1'b0;  wr_cycle[16072] = 1'b1;  addr_rom[16072]='h00001a24;  wr_data_rom[16072]='h000017a3;
    rd_cycle[16073] = 1'b0;  wr_cycle[16073] = 1'b1;  addr_rom[16073]='h00001eb4;  wr_data_rom[16073]='h00000eec;
    rd_cycle[16074] = 1'b1;  wr_cycle[16074] = 1'b0;  addr_rom[16074]='h00003ce0;  wr_data_rom[16074]='h00000000;
    rd_cycle[16075] = 1'b0;  wr_cycle[16075] = 1'b1;  addr_rom[16075]='h00000c60;  wr_data_rom[16075]='h00002daa;
    rd_cycle[16076] = 1'b0;  wr_cycle[16076] = 1'b1;  addr_rom[16076]='h00003890;  wr_data_rom[16076]='h0000232d;
    rd_cycle[16077] = 1'b0;  wr_cycle[16077] = 1'b1;  addr_rom[16077]='h0000234c;  wr_data_rom[16077]='h00003059;
    rd_cycle[16078] = 1'b1;  wr_cycle[16078] = 1'b0;  addr_rom[16078]='h000022bc;  wr_data_rom[16078]='h00000000;
    rd_cycle[16079] = 1'b1;  wr_cycle[16079] = 1'b0;  addr_rom[16079]='h00003260;  wr_data_rom[16079]='h00000000;
    rd_cycle[16080] = 1'b1;  wr_cycle[16080] = 1'b0;  addr_rom[16080]='h00000c6c;  wr_data_rom[16080]='h00000000;
    rd_cycle[16081] = 1'b1;  wr_cycle[16081] = 1'b0;  addr_rom[16081]='h000007e8;  wr_data_rom[16081]='h00000000;
    rd_cycle[16082] = 1'b1;  wr_cycle[16082] = 1'b0;  addr_rom[16082]='h0000188c;  wr_data_rom[16082]='h00000000;
    rd_cycle[16083] = 1'b1;  wr_cycle[16083] = 1'b0;  addr_rom[16083]='h0000062c;  wr_data_rom[16083]='h00000000;
    rd_cycle[16084] = 1'b0;  wr_cycle[16084] = 1'b1;  addr_rom[16084]='h00002bdc;  wr_data_rom[16084]='h0000187e;
    rd_cycle[16085] = 1'b0;  wr_cycle[16085] = 1'b1;  addr_rom[16085]='h00000b90;  wr_data_rom[16085]='h00001f69;
    rd_cycle[16086] = 1'b1;  wr_cycle[16086] = 1'b0;  addr_rom[16086]='h000013dc;  wr_data_rom[16086]='h00000000;
    rd_cycle[16087] = 1'b1;  wr_cycle[16087] = 1'b0;  addr_rom[16087]='h000004f4;  wr_data_rom[16087]='h00000000;
    rd_cycle[16088] = 1'b1;  wr_cycle[16088] = 1'b0;  addr_rom[16088]='h00002a90;  wr_data_rom[16088]='h00000000;
    rd_cycle[16089] = 1'b1;  wr_cycle[16089] = 1'b0;  addr_rom[16089]='h00000dd0;  wr_data_rom[16089]='h00000000;
    rd_cycle[16090] = 1'b0;  wr_cycle[16090] = 1'b1;  addr_rom[16090]='h000025d4;  wr_data_rom[16090]='h00000418;
    rd_cycle[16091] = 1'b0;  wr_cycle[16091] = 1'b1;  addr_rom[16091]='h00001e00;  wr_data_rom[16091]='h00002963;
    rd_cycle[16092] = 1'b0;  wr_cycle[16092] = 1'b1;  addr_rom[16092]='h00002450;  wr_data_rom[16092]='h000031ba;
    rd_cycle[16093] = 1'b0;  wr_cycle[16093] = 1'b1;  addr_rom[16093]='h00003bb4;  wr_data_rom[16093]='h00001f35;
    rd_cycle[16094] = 1'b0;  wr_cycle[16094] = 1'b1;  addr_rom[16094]='h000016ec;  wr_data_rom[16094]='h00001e30;
    rd_cycle[16095] = 1'b1;  wr_cycle[16095] = 1'b0;  addr_rom[16095]='h00003bb4;  wr_data_rom[16095]='h00000000;
    rd_cycle[16096] = 1'b0;  wr_cycle[16096] = 1'b1;  addr_rom[16096]='h00001ae4;  wr_data_rom[16096]='h00000a70;
    rd_cycle[16097] = 1'b0;  wr_cycle[16097] = 1'b1;  addr_rom[16097]='h00001200;  wr_data_rom[16097]='h00000dc5;
    rd_cycle[16098] = 1'b0;  wr_cycle[16098] = 1'b1;  addr_rom[16098]='h00002804;  wr_data_rom[16098]='h000013e9;
    rd_cycle[16099] = 1'b1;  wr_cycle[16099] = 1'b0;  addr_rom[16099]='h00000410;  wr_data_rom[16099]='h00000000;
    rd_cycle[16100] = 1'b0;  wr_cycle[16100] = 1'b1;  addr_rom[16100]='h00002d70;  wr_data_rom[16100]='h00003066;
    rd_cycle[16101] = 1'b0;  wr_cycle[16101] = 1'b1;  addr_rom[16101]='h00003ea8;  wr_data_rom[16101]='h000023de;
    rd_cycle[16102] = 1'b1;  wr_cycle[16102] = 1'b0;  addr_rom[16102]='h0000333c;  wr_data_rom[16102]='h00000000;
    rd_cycle[16103] = 1'b1;  wr_cycle[16103] = 1'b0;  addr_rom[16103]='h000023a4;  wr_data_rom[16103]='h00000000;
    rd_cycle[16104] = 1'b1;  wr_cycle[16104] = 1'b0;  addr_rom[16104]='h00000b78;  wr_data_rom[16104]='h00000000;
    rd_cycle[16105] = 1'b0;  wr_cycle[16105] = 1'b1;  addr_rom[16105]='h00003918;  wr_data_rom[16105]='h00003f5f;
    rd_cycle[16106] = 1'b0;  wr_cycle[16106] = 1'b1;  addr_rom[16106]='h00001ce4;  wr_data_rom[16106]='h00003544;
    rd_cycle[16107] = 1'b0;  wr_cycle[16107] = 1'b1;  addr_rom[16107]='h00003c40;  wr_data_rom[16107]='h00001177;
    rd_cycle[16108] = 1'b0;  wr_cycle[16108] = 1'b1;  addr_rom[16108]='h000039c0;  wr_data_rom[16108]='h0000130a;
    rd_cycle[16109] = 1'b0;  wr_cycle[16109] = 1'b1;  addr_rom[16109]='h00001030;  wr_data_rom[16109]='h0000268b;
    rd_cycle[16110] = 1'b1;  wr_cycle[16110] = 1'b0;  addr_rom[16110]='h00003ff8;  wr_data_rom[16110]='h00000000;
    rd_cycle[16111] = 1'b1;  wr_cycle[16111] = 1'b0;  addr_rom[16111]='h000009cc;  wr_data_rom[16111]='h00000000;
    rd_cycle[16112] = 1'b1;  wr_cycle[16112] = 1'b0;  addr_rom[16112]='h000028d4;  wr_data_rom[16112]='h00000000;
    rd_cycle[16113] = 1'b0;  wr_cycle[16113] = 1'b1;  addr_rom[16113]='h0000349c;  wr_data_rom[16113]='h000027da;
    rd_cycle[16114] = 1'b0;  wr_cycle[16114] = 1'b1;  addr_rom[16114]='h000013a0;  wr_data_rom[16114]='h0000346a;
    rd_cycle[16115] = 1'b0;  wr_cycle[16115] = 1'b1;  addr_rom[16115]='h00001d80;  wr_data_rom[16115]='h000032d0;
    rd_cycle[16116] = 1'b1;  wr_cycle[16116] = 1'b0;  addr_rom[16116]='h000016e0;  wr_data_rom[16116]='h00000000;
    rd_cycle[16117] = 1'b1;  wr_cycle[16117] = 1'b0;  addr_rom[16117]='h00002f2c;  wr_data_rom[16117]='h00000000;
    rd_cycle[16118] = 1'b1;  wr_cycle[16118] = 1'b0;  addr_rom[16118]='h00003c10;  wr_data_rom[16118]='h00000000;
    rd_cycle[16119] = 1'b1;  wr_cycle[16119] = 1'b0;  addr_rom[16119]='h00003834;  wr_data_rom[16119]='h00000000;
    rd_cycle[16120] = 1'b0;  wr_cycle[16120] = 1'b1;  addr_rom[16120]='h00000f38;  wr_data_rom[16120]='h00003686;
    rd_cycle[16121] = 1'b0;  wr_cycle[16121] = 1'b1;  addr_rom[16121]='h00003b28;  wr_data_rom[16121]='h00002fce;
    rd_cycle[16122] = 1'b1;  wr_cycle[16122] = 1'b0;  addr_rom[16122]='h0000227c;  wr_data_rom[16122]='h00000000;
    rd_cycle[16123] = 1'b1;  wr_cycle[16123] = 1'b0;  addr_rom[16123]='h00001bb0;  wr_data_rom[16123]='h00000000;
    rd_cycle[16124] = 1'b0;  wr_cycle[16124] = 1'b1;  addr_rom[16124]='h00000188;  wr_data_rom[16124]='h000038d0;
    rd_cycle[16125] = 1'b0;  wr_cycle[16125] = 1'b1;  addr_rom[16125]='h00002da8;  wr_data_rom[16125]='h0000358b;
    rd_cycle[16126] = 1'b1;  wr_cycle[16126] = 1'b0;  addr_rom[16126]='h0000221c;  wr_data_rom[16126]='h00000000;
    rd_cycle[16127] = 1'b1;  wr_cycle[16127] = 1'b0;  addr_rom[16127]='h00001a80;  wr_data_rom[16127]='h00000000;
    rd_cycle[16128] = 1'b1;  wr_cycle[16128] = 1'b0;  addr_rom[16128]='h000037f0;  wr_data_rom[16128]='h00000000;
    rd_cycle[16129] = 1'b1;  wr_cycle[16129] = 1'b0;  addr_rom[16129]='h00003580;  wr_data_rom[16129]='h00000000;
    rd_cycle[16130] = 1'b1;  wr_cycle[16130] = 1'b0;  addr_rom[16130]='h00002620;  wr_data_rom[16130]='h00000000;
    rd_cycle[16131] = 1'b0;  wr_cycle[16131] = 1'b1;  addr_rom[16131]='h00003f40;  wr_data_rom[16131]='h0000075c;
    rd_cycle[16132] = 1'b1;  wr_cycle[16132] = 1'b0;  addr_rom[16132]='h00003d88;  wr_data_rom[16132]='h00000000;
    rd_cycle[16133] = 1'b0;  wr_cycle[16133] = 1'b1;  addr_rom[16133]='h000022bc;  wr_data_rom[16133]='h000021ec;
    rd_cycle[16134] = 1'b0;  wr_cycle[16134] = 1'b1;  addr_rom[16134]='h00003c90;  wr_data_rom[16134]='h0000076a;
    rd_cycle[16135] = 1'b1;  wr_cycle[16135] = 1'b0;  addr_rom[16135]='h00000f48;  wr_data_rom[16135]='h00000000;
    rd_cycle[16136] = 1'b1;  wr_cycle[16136] = 1'b0;  addr_rom[16136]='h00000a08;  wr_data_rom[16136]='h00000000;
    rd_cycle[16137] = 1'b0;  wr_cycle[16137] = 1'b1;  addr_rom[16137]='h00002ddc;  wr_data_rom[16137]='h00003c5e;
    rd_cycle[16138] = 1'b0;  wr_cycle[16138] = 1'b1;  addr_rom[16138]='h00001470;  wr_data_rom[16138]='h000037c2;
    rd_cycle[16139] = 1'b0;  wr_cycle[16139] = 1'b1;  addr_rom[16139]='h00002d00;  wr_data_rom[16139]='h0000363f;
    rd_cycle[16140] = 1'b1;  wr_cycle[16140] = 1'b0;  addr_rom[16140]='h00002594;  wr_data_rom[16140]='h00000000;
    rd_cycle[16141] = 1'b1;  wr_cycle[16141] = 1'b0;  addr_rom[16141]='h00000ee4;  wr_data_rom[16141]='h00000000;
    rd_cycle[16142] = 1'b0;  wr_cycle[16142] = 1'b1;  addr_rom[16142]='h00003030;  wr_data_rom[16142]='h00001349;
    rd_cycle[16143] = 1'b0;  wr_cycle[16143] = 1'b1;  addr_rom[16143]='h000011cc;  wr_data_rom[16143]='h00003ee7;
    rd_cycle[16144] = 1'b1;  wr_cycle[16144] = 1'b0;  addr_rom[16144]='h00001448;  wr_data_rom[16144]='h00000000;
    rd_cycle[16145] = 1'b1;  wr_cycle[16145] = 1'b0;  addr_rom[16145]='h00000c1c;  wr_data_rom[16145]='h00000000;
    rd_cycle[16146] = 1'b1;  wr_cycle[16146] = 1'b0;  addr_rom[16146]='h000039cc;  wr_data_rom[16146]='h00000000;
    rd_cycle[16147] = 1'b0;  wr_cycle[16147] = 1'b1;  addr_rom[16147]='h000019f4;  wr_data_rom[16147]='h000015f6;
    rd_cycle[16148] = 1'b1;  wr_cycle[16148] = 1'b0;  addr_rom[16148]='h00002fd4;  wr_data_rom[16148]='h00000000;
    rd_cycle[16149] = 1'b1;  wr_cycle[16149] = 1'b0;  addr_rom[16149]='h00002388;  wr_data_rom[16149]='h00000000;
    rd_cycle[16150] = 1'b0;  wr_cycle[16150] = 1'b1;  addr_rom[16150]='h0000266c;  wr_data_rom[16150]='h000012e3;
    rd_cycle[16151] = 1'b1;  wr_cycle[16151] = 1'b0;  addr_rom[16151]='h00000284;  wr_data_rom[16151]='h00000000;
    rd_cycle[16152] = 1'b0;  wr_cycle[16152] = 1'b1;  addr_rom[16152]='h000021c4;  wr_data_rom[16152]='h00003b22;
    rd_cycle[16153] = 1'b1;  wr_cycle[16153] = 1'b0;  addr_rom[16153]='h0000394c;  wr_data_rom[16153]='h00000000;
    rd_cycle[16154] = 1'b1;  wr_cycle[16154] = 1'b0;  addr_rom[16154]='h00000624;  wr_data_rom[16154]='h00000000;
    rd_cycle[16155] = 1'b1;  wr_cycle[16155] = 1'b0;  addr_rom[16155]='h00000f80;  wr_data_rom[16155]='h00000000;
    rd_cycle[16156] = 1'b1;  wr_cycle[16156] = 1'b0;  addr_rom[16156]='h00000b60;  wr_data_rom[16156]='h00000000;
    rd_cycle[16157] = 1'b1;  wr_cycle[16157] = 1'b0;  addr_rom[16157]='h00000b50;  wr_data_rom[16157]='h00000000;
    rd_cycle[16158] = 1'b1;  wr_cycle[16158] = 1'b0;  addr_rom[16158]='h00002c30;  wr_data_rom[16158]='h00000000;
    rd_cycle[16159] = 1'b1;  wr_cycle[16159] = 1'b0;  addr_rom[16159]='h00003580;  wr_data_rom[16159]='h00000000;
    rd_cycle[16160] = 1'b0;  wr_cycle[16160] = 1'b1;  addr_rom[16160]='h00000754;  wr_data_rom[16160]='h00002766;
    rd_cycle[16161] = 1'b0;  wr_cycle[16161] = 1'b1;  addr_rom[16161]='h00000520;  wr_data_rom[16161]='h00001053;
    rd_cycle[16162] = 1'b0;  wr_cycle[16162] = 1'b1;  addr_rom[16162]='h00002540;  wr_data_rom[16162]='h00001c82;
    rd_cycle[16163] = 1'b0;  wr_cycle[16163] = 1'b1;  addr_rom[16163]='h0000036c;  wr_data_rom[16163]='h0000024a;
    rd_cycle[16164] = 1'b1;  wr_cycle[16164] = 1'b0;  addr_rom[16164]='h000018b8;  wr_data_rom[16164]='h00000000;
    rd_cycle[16165] = 1'b0;  wr_cycle[16165] = 1'b1;  addr_rom[16165]='h00002af4;  wr_data_rom[16165]='h000012e5;
    rd_cycle[16166] = 1'b1;  wr_cycle[16166] = 1'b0;  addr_rom[16166]='h00002e60;  wr_data_rom[16166]='h00000000;
    rd_cycle[16167] = 1'b1;  wr_cycle[16167] = 1'b0;  addr_rom[16167]='h000007a4;  wr_data_rom[16167]='h00000000;
    rd_cycle[16168] = 1'b1;  wr_cycle[16168] = 1'b0;  addr_rom[16168]='h000026f8;  wr_data_rom[16168]='h00000000;
    rd_cycle[16169] = 1'b1;  wr_cycle[16169] = 1'b0;  addr_rom[16169]='h000000fc;  wr_data_rom[16169]='h00000000;
    rd_cycle[16170] = 1'b1;  wr_cycle[16170] = 1'b0;  addr_rom[16170]='h000012fc;  wr_data_rom[16170]='h00000000;
    rd_cycle[16171] = 1'b0;  wr_cycle[16171] = 1'b1;  addr_rom[16171]='h000007e4;  wr_data_rom[16171]='h000025e3;
    rd_cycle[16172] = 1'b0;  wr_cycle[16172] = 1'b1;  addr_rom[16172]='h000024e4;  wr_data_rom[16172]='h000020d6;
    rd_cycle[16173] = 1'b1;  wr_cycle[16173] = 1'b0;  addr_rom[16173]='h00002364;  wr_data_rom[16173]='h00000000;
    rd_cycle[16174] = 1'b1;  wr_cycle[16174] = 1'b0;  addr_rom[16174]='h00001774;  wr_data_rom[16174]='h00000000;
    rd_cycle[16175] = 1'b0;  wr_cycle[16175] = 1'b1;  addr_rom[16175]='h00000ef8;  wr_data_rom[16175]='h00000c5b;
    rd_cycle[16176] = 1'b0;  wr_cycle[16176] = 1'b1;  addr_rom[16176]='h00003cc8;  wr_data_rom[16176]='h0000351c;
    rd_cycle[16177] = 1'b1;  wr_cycle[16177] = 1'b0;  addr_rom[16177]='h00001638;  wr_data_rom[16177]='h00000000;
    rd_cycle[16178] = 1'b0;  wr_cycle[16178] = 1'b1;  addr_rom[16178]='h0000224c;  wr_data_rom[16178]='h00003a48;
    rd_cycle[16179] = 1'b1;  wr_cycle[16179] = 1'b0;  addr_rom[16179]='h00001ab8;  wr_data_rom[16179]='h00000000;
    rd_cycle[16180] = 1'b1;  wr_cycle[16180] = 1'b0;  addr_rom[16180]='h000039f4;  wr_data_rom[16180]='h00000000;
    rd_cycle[16181] = 1'b0;  wr_cycle[16181] = 1'b1;  addr_rom[16181]='h00000188;  wr_data_rom[16181]='h00001176;
    rd_cycle[16182] = 1'b0;  wr_cycle[16182] = 1'b1;  addr_rom[16182]='h00000b68;  wr_data_rom[16182]='h0000306c;
    rd_cycle[16183] = 1'b0;  wr_cycle[16183] = 1'b1;  addr_rom[16183]='h00003d78;  wr_data_rom[16183]='h000025be;
    rd_cycle[16184] = 1'b1;  wr_cycle[16184] = 1'b0;  addr_rom[16184]='h00001048;  wr_data_rom[16184]='h00000000;
    rd_cycle[16185] = 1'b0;  wr_cycle[16185] = 1'b1;  addr_rom[16185]='h00002568;  wr_data_rom[16185]='h00003272;
    rd_cycle[16186] = 1'b1;  wr_cycle[16186] = 1'b0;  addr_rom[16186]='h00000a74;  wr_data_rom[16186]='h00000000;
    rd_cycle[16187] = 1'b1;  wr_cycle[16187] = 1'b0;  addr_rom[16187]='h00001f04;  wr_data_rom[16187]='h00000000;
    rd_cycle[16188] = 1'b0;  wr_cycle[16188] = 1'b1;  addr_rom[16188]='h00001ac4;  wr_data_rom[16188]='h00003276;
    rd_cycle[16189] = 1'b1;  wr_cycle[16189] = 1'b0;  addr_rom[16189]='h00001f6c;  wr_data_rom[16189]='h00000000;
    rd_cycle[16190] = 1'b1;  wr_cycle[16190] = 1'b0;  addr_rom[16190]='h00000cd0;  wr_data_rom[16190]='h00000000;
    rd_cycle[16191] = 1'b1;  wr_cycle[16191] = 1'b0;  addr_rom[16191]='h00001424;  wr_data_rom[16191]='h00000000;
    rd_cycle[16192] = 1'b1;  wr_cycle[16192] = 1'b0;  addr_rom[16192]='h00002328;  wr_data_rom[16192]='h00000000;
    rd_cycle[16193] = 1'b1;  wr_cycle[16193] = 1'b0;  addr_rom[16193]='h00001a74;  wr_data_rom[16193]='h00000000;
    rd_cycle[16194] = 1'b0;  wr_cycle[16194] = 1'b1;  addr_rom[16194]='h00003f0c;  wr_data_rom[16194]='h0000220a;
    rd_cycle[16195] = 1'b1;  wr_cycle[16195] = 1'b0;  addr_rom[16195]='h00000f88;  wr_data_rom[16195]='h00000000;
    rd_cycle[16196] = 1'b0;  wr_cycle[16196] = 1'b1;  addr_rom[16196]='h00002944;  wr_data_rom[16196]='h0000362f;
    rd_cycle[16197] = 1'b1;  wr_cycle[16197] = 1'b0;  addr_rom[16197]='h000020fc;  wr_data_rom[16197]='h00000000;
    rd_cycle[16198] = 1'b0;  wr_cycle[16198] = 1'b1;  addr_rom[16198]='h00001c74;  wr_data_rom[16198]='h00000dda;
    rd_cycle[16199] = 1'b0;  wr_cycle[16199] = 1'b1;  addr_rom[16199]='h000017f4;  wr_data_rom[16199]='h00003926;
    rd_cycle[16200] = 1'b1;  wr_cycle[16200] = 1'b0;  addr_rom[16200]='h00002dac;  wr_data_rom[16200]='h00000000;
    rd_cycle[16201] = 1'b0;  wr_cycle[16201] = 1'b1;  addr_rom[16201]='h00003c0c;  wr_data_rom[16201]='h0000090a;
    rd_cycle[16202] = 1'b1;  wr_cycle[16202] = 1'b0;  addr_rom[16202]='h00003740;  wr_data_rom[16202]='h00000000;
    rd_cycle[16203] = 1'b0;  wr_cycle[16203] = 1'b1;  addr_rom[16203]='h00002204;  wr_data_rom[16203]='h00000827;
    rd_cycle[16204] = 1'b0;  wr_cycle[16204] = 1'b1;  addr_rom[16204]='h00002a20;  wr_data_rom[16204]='h00002ac6;
    rd_cycle[16205] = 1'b1;  wr_cycle[16205] = 1'b0;  addr_rom[16205]='h000020a4;  wr_data_rom[16205]='h00000000;
    rd_cycle[16206] = 1'b1;  wr_cycle[16206] = 1'b0;  addr_rom[16206]='h000012c0;  wr_data_rom[16206]='h00000000;
    rd_cycle[16207] = 1'b1;  wr_cycle[16207] = 1'b0;  addr_rom[16207]='h00000d90;  wr_data_rom[16207]='h00000000;
    rd_cycle[16208] = 1'b0;  wr_cycle[16208] = 1'b1;  addr_rom[16208]='h00001d24;  wr_data_rom[16208]='h000029e7;
    rd_cycle[16209] = 1'b1;  wr_cycle[16209] = 1'b0;  addr_rom[16209]='h00000b48;  wr_data_rom[16209]='h00000000;
    rd_cycle[16210] = 1'b1;  wr_cycle[16210] = 1'b0;  addr_rom[16210]='h000022f0;  wr_data_rom[16210]='h00000000;
    rd_cycle[16211] = 1'b0;  wr_cycle[16211] = 1'b1;  addr_rom[16211]='h0000142c;  wr_data_rom[16211]='h00003a77;
    rd_cycle[16212] = 1'b0;  wr_cycle[16212] = 1'b1;  addr_rom[16212]='h00000b84;  wr_data_rom[16212]='h0000169d;
    rd_cycle[16213] = 1'b0;  wr_cycle[16213] = 1'b1;  addr_rom[16213]='h000006a8;  wr_data_rom[16213]='h000009df;
    rd_cycle[16214] = 1'b0;  wr_cycle[16214] = 1'b1;  addr_rom[16214]='h00000658;  wr_data_rom[16214]='h00002977;
    rd_cycle[16215] = 1'b1;  wr_cycle[16215] = 1'b0;  addr_rom[16215]='h00002c24;  wr_data_rom[16215]='h00000000;
    rd_cycle[16216] = 1'b1;  wr_cycle[16216] = 1'b0;  addr_rom[16216]='h000015ec;  wr_data_rom[16216]='h00000000;
    rd_cycle[16217] = 1'b1;  wr_cycle[16217] = 1'b0;  addr_rom[16217]='h000001d0;  wr_data_rom[16217]='h00000000;
    rd_cycle[16218] = 1'b1;  wr_cycle[16218] = 1'b0;  addr_rom[16218]='h00000bd8;  wr_data_rom[16218]='h00000000;
    rd_cycle[16219] = 1'b1;  wr_cycle[16219] = 1'b0;  addr_rom[16219]='h000034b0;  wr_data_rom[16219]='h00000000;
    rd_cycle[16220] = 1'b1;  wr_cycle[16220] = 1'b0;  addr_rom[16220]='h000021f8;  wr_data_rom[16220]='h00000000;
    rd_cycle[16221] = 1'b1;  wr_cycle[16221] = 1'b0;  addr_rom[16221]='h00001eb8;  wr_data_rom[16221]='h00000000;
    rd_cycle[16222] = 1'b1;  wr_cycle[16222] = 1'b0;  addr_rom[16222]='h000020b8;  wr_data_rom[16222]='h00000000;
    rd_cycle[16223] = 1'b0;  wr_cycle[16223] = 1'b1;  addr_rom[16223]='h00000594;  wr_data_rom[16223]='h00001911;
    rd_cycle[16224] = 1'b1;  wr_cycle[16224] = 1'b0;  addr_rom[16224]='h00003c98;  wr_data_rom[16224]='h00000000;
    rd_cycle[16225] = 1'b1;  wr_cycle[16225] = 1'b0;  addr_rom[16225]='h00002e88;  wr_data_rom[16225]='h00000000;
    rd_cycle[16226] = 1'b0;  wr_cycle[16226] = 1'b1;  addr_rom[16226]='h00001e60;  wr_data_rom[16226]='h00003882;
    rd_cycle[16227] = 1'b0;  wr_cycle[16227] = 1'b1;  addr_rom[16227]='h00003a74;  wr_data_rom[16227]='h00000b77;
    rd_cycle[16228] = 1'b0;  wr_cycle[16228] = 1'b1;  addr_rom[16228]='h00003638;  wr_data_rom[16228]='h00002f45;
    rd_cycle[16229] = 1'b0;  wr_cycle[16229] = 1'b1;  addr_rom[16229]='h00000b38;  wr_data_rom[16229]='h00003861;
    rd_cycle[16230] = 1'b1;  wr_cycle[16230] = 1'b0;  addr_rom[16230]='h00000888;  wr_data_rom[16230]='h00000000;
    rd_cycle[16231] = 1'b0;  wr_cycle[16231] = 1'b1;  addr_rom[16231]='h00003d04;  wr_data_rom[16231]='h00000fb6;
    rd_cycle[16232] = 1'b1;  wr_cycle[16232] = 1'b0;  addr_rom[16232]='h00003798;  wr_data_rom[16232]='h00000000;
    rd_cycle[16233] = 1'b1;  wr_cycle[16233] = 1'b0;  addr_rom[16233]='h00000a08;  wr_data_rom[16233]='h00000000;
    rd_cycle[16234] = 1'b1;  wr_cycle[16234] = 1'b0;  addr_rom[16234]='h000001dc;  wr_data_rom[16234]='h00000000;
    rd_cycle[16235] = 1'b0;  wr_cycle[16235] = 1'b1;  addr_rom[16235]='h000004d4;  wr_data_rom[16235]='h000003c3;
    rd_cycle[16236] = 1'b1;  wr_cycle[16236] = 1'b0;  addr_rom[16236]='h00000948;  wr_data_rom[16236]='h00000000;
    rd_cycle[16237] = 1'b0;  wr_cycle[16237] = 1'b1;  addr_rom[16237]='h00000af8;  wr_data_rom[16237]='h0000094f;
    rd_cycle[16238] = 1'b0;  wr_cycle[16238] = 1'b1;  addr_rom[16238]='h00001754;  wr_data_rom[16238]='h00000b72;
    rd_cycle[16239] = 1'b1;  wr_cycle[16239] = 1'b0;  addr_rom[16239]='h000010f8;  wr_data_rom[16239]='h00000000;
    rd_cycle[16240] = 1'b0;  wr_cycle[16240] = 1'b1;  addr_rom[16240]='h00003ba0;  wr_data_rom[16240]='h00002af2;
    rd_cycle[16241] = 1'b1;  wr_cycle[16241] = 1'b0;  addr_rom[16241]='h00002624;  wr_data_rom[16241]='h00000000;
    rd_cycle[16242] = 1'b1;  wr_cycle[16242] = 1'b0;  addr_rom[16242]='h00003c14;  wr_data_rom[16242]='h00000000;
    rd_cycle[16243] = 1'b0;  wr_cycle[16243] = 1'b1;  addr_rom[16243]='h00001c88;  wr_data_rom[16243]='h00000b6c;
    rd_cycle[16244] = 1'b0;  wr_cycle[16244] = 1'b1;  addr_rom[16244]='h000000fc;  wr_data_rom[16244]='h00002e09;
    rd_cycle[16245] = 1'b1;  wr_cycle[16245] = 1'b0;  addr_rom[16245]='h00001ff8;  wr_data_rom[16245]='h00000000;
    rd_cycle[16246] = 1'b0;  wr_cycle[16246] = 1'b1;  addr_rom[16246]='h00002bc0;  wr_data_rom[16246]='h00003ef1;
    rd_cycle[16247] = 1'b1;  wr_cycle[16247] = 1'b0;  addr_rom[16247]='h000005f8;  wr_data_rom[16247]='h00000000;
    rd_cycle[16248] = 1'b1;  wr_cycle[16248] = 1'b0;  addr_rom[16248]='h0000204c;  wr_data_rom[16248]='h00000000;
    rd_cycle[16249] = 1'b0;  wr_cycle[16249] = 1'b1;  addr_rom[16249]='h00000930;  wr_data_rom[16249]='h00003baa;
    rd_cycle[16250] = 1'b0;  wr_cycle[16250] = 1'b1;  addr_rom[16250]='h00000da8;  wr_data_rom[16250]='h00002e13;
    rd_cycle[16251] = 1'b0;  wr_cycle[16251] = 1'b1;  addr_rom[16251]='h00003ab4;  wr_data_rom[16251]='h00002c1b;
    rd_cycle[16252] = 1'b1;  wr_cycle[16252] = 1'b0;  addr_rom[16252]='h000026a0;  wr_data_rom[16252]='h00000000;
    rd_cycle[16253] = 1'b1;  wr_cycle[16253] = 1'b0;  addr_rom[16253]='h00001f74;  wr_data_rom[16253]='h00000000;
    rd_cycle[16254] = 1'b0;  wr_cycle[16254] = 1'b1;  addr_rom[16254]='h00002b70;  wr_data_rom[16254]='h00001ad0;
    rd_cycle[16255] = 1'b0;  wr_cycle[16255] = 1'b1;  addr_rom[16255]='h00002b94;  wr_data_rom[16255]='h00002580;
    rd_cycle[16256] = 1'b0;  wr_cycle[16256] = 1'b1;  addr_rom[16256]='h000011d4;  wr_data_rom[16256]='h00002115;
    rd_cycle[16257] = 1'b1;  wr_cycle[16257] = 1'b0;  addr_rom[16257]='h00001e4c;  wr_data_rom[16257]='h00000000;
    rd_cycle[16258] = 1'b0;  wr_cycle[16258] = 1'b1;  addr_rom[16258]='h00001afc;  wr_data_rom[16258]='h00000067;
    rd_cycle[16259] = 1'b1;  wr_cycle[16259] = 1'b0;  addr_rom[16259]='h000017c8;  wr_data_rom[16259]='h00000000;
    rd_cycle[16260] = 1'b1;  wr_cycle[16260] = 1'b0;  addr_rom[16260]='h00003fd8;  wr_data_rom[16260]='h00000000;
    rd_cycle[16261] = 1'b0;  wr_cycle[16261] = 1'b1;  addr_rom[16261]='h00003c84;  wr_data_rom[16261]='h0000050c;
    rd_cycle[16262] = 1'b1;  wr_cycle[16262] = 1'b0;  addr_rom[16262]='h000033ac;  wr_data_rom[16262]='h00000000;
    rd_cycle[16263] = 1'b0;  wr_cycle[16263] = 1'b1;  addr_rom[16263]='h00003a7c;  wr_data_rom[16263]='h00003185;
    rd_cycle[16264] = 1'b0;  wr_cycle[16264] = 1'b1;  addr_rom[16264]='h00000650;  wr_data_rom[16264]='h00001574;
    rd_cycle[16265] = 1'b1;  wr_cycle[16265] = 1'b0;  addr_rom[16265]='h00003fcc;  wr_data_rom[16265]='h00000000;
    rd_cycle[16266] = 1'b0;  wr_cycle[16266] = 1'b1;  addr_rom[16266]='h00003b64;  wr_data_rom[16266]='h00000928;
    rd_cycle[16267] = 1'b1;  wr_cycle[16267] = 1'b0;  addr_rom[16267]='h00001214;  wr_data_rom[16267]='h00000000;
    rd_cycle[16268] = 1'b1;  wr_cycle[16268] = 1'b0;  addr_rom[16268]='h00000cdc;  wr_data_rom[16268]='h00000000;
    rd_cycle[16269] = 1'b1;  wr_cycle[16269] = 1'b0;  addr_rom[16269]='h00000e78;  wr_data_rom[16269]='h00000000;
    rd_cycle[16270] = 1'b1;  wr_cycle[16270] = 1'b0;  addr_rom[16270]='h00003fb8;  wr_data_rom[16270]='h00000000;
    rd_cycle[16271] = 1'b0;  wr_cycle[16271] = 1'b1;  addr_rom[16271]='h000006ec;  wr_data_rom[16271]='h000010a3;
    rd_cycle[16272] = 1'b0;  wr_cycle[16272] = 1'b1;  addr_rom[16272]='h00002830;  wr_data_rom[16272]='h00000ce1;
    rd_cycle[16273] = 1'b1;  wr_cycle[16273] = 1'b0;  addr_rom[16273]='h000030b0;  wr_data_rom[16273]='h00000000;
    rd_cycle[16274] = 1'b0;  wr_cycle[16274] = 1'b1;  addr_rom[16274]='h00002298;  wr_data_rom[16274]='h00001e16;
    rd_cycle[16275] = 1'b1;  wr_cycle[16275] = 1'b0;  addr_rom[16275]='h00000d48;  wr_data_rom[16275]='h00000000;
    rd_cycle[16276] = 1'b0;  wr_cycle[16276] = 1'b1;  addr_rom[16276]='h0000187c;  wr_data_rom[16276]='h0000081c;
    rd_cycle[16277] = 1'b0;  wr_cycle[16277] = 1'b1;  addr_rom[16277]='h00001a0c;  wr_data_rom[16277]='h00000dde;
    rd_cycle[16278] = 1'b1;  wr_cycle[16278] = 1'b0;  addr_rom[16278]='h00000578;  wr_data_rom[16278]='h00000000;
    rd_cycle[16279] = 1'b0;  wr_cycle[16279] = 1'b1;  addr_rom[16279]='h000015a8;  wr_data_rom[16279]='h000009c0;
    rd_cycle[16280] = 1'b1;  wr_cycle[16280] = 1'b0;  addr_rom[16280]='h000018b0;  wr_data_rom[16280]='h00000000;
    rd_cycle[16281] = 1'b1;  wr_cycle[16281] = 1'b0;  addr_rom[16281]='h00003948;  wr_data_rom[16281]='h00000000;
    rd_cycle[16282] = 1'b1;  wr_cycle[16282] = 1'b0;  addr_rom[16282]='h00003fec;  wr_data_rom[16282]='h00000000;
    rd_cycle[16283] = 1'b1;  wr_cycle[16283] = 1'b0;  addr_rom[16283]='h000023f8;  wr_data_rom[16283]='h00000000;
    rd_cycle[16284] = 1'b1;  wr_cycle[16284] = 1'b0;  addr_rom[16284]='h00001de4;  wr_data_rom[16284]='h00000000;
    rd_cycle[16285] = 1'b0;  wr_cycle[16285] = 1'b1;  addr_rom[16285]='h000039b8;  wr_data_rom[16285]='h000004b7;
    rd_cycle[16286] = 1'b1;  wr_cycle[16286] = 1'b0;  addr_rom[16286]='h00003c9c;  wr_data_rom[16286]='h00000000;
    rd_cycle[16287] = 1'b0;  wr_cycle[16287] = 1'b1;  addr_rom[16287]='h000001c4;  wr_data_rom[16287]='h00000706;
    rd_cycle[16288] = 1'b1;  wr_cycle[16288] = 1'b0;  addr_rom[16288]='h00003f20;  wr_data_rom[16288]='h00000000;
    rd_cycle[16289] = 1'b0;  wr_cycle[16289] = 1'b1;  addr_rom[16289]='h00001c94;  wr_data_rom[16289]='h00001d23;
    rd_cycle[16290] = 1'b1;  wr_cycle[16290] = 1'b0;  addr_rom[16290]='h000019dc;  wr_data_rom[16290]='h00000000;
    rd_cycle[16291] = 1'b1;  wr_cycle[16291] = 1'b0;  addr_rom[16291]='h0000155c;  wr_data_rom[16291]='h00000000;
    rd_cycle[16292] = 1'b0;  wr_cycle[16292] = 1'b1;  addr_rom[16292]='h00001700;  wr_data_rom[16292]='h00002421;
    rd_cycle[16293] = 1'b1;  wr_cycle[16293] = 1'b0;  addr_rom[16293]='h00001aa8;  wr_data_rom[16293]='h00000000;
    rd_cycle[16294] = 1'b1;  wr_cycle[16294] = 1'b0;  addr_rom[16294]='h0000001c;  wr_data_rom[16294]='h00000000;
    rd_cycle[16295] = 1'b0;  wr_cycle[16295] = 1'b1;  addr_rom[16295]='h00001d70;  wr_data_rom[16295]='h000020b8;
    rd_cycle[16296] = 1'b0;  wr_cycle[16296] = 1'b1;  addr_rom[16296]='h00003448;  wr_data_rom[16296]='h00002f21;
    rd_cycle[16297] = 1'b1;  wr_cycle[16297] = 1'b0;  addr_rom[16297]='h00003970;  wr_data_rom[16297]='h00000000;
    rd_cycle[16298] = 1'b1;  wr_cycle[16298] = 1'b0;  addr_rom[16298]='h0000158c;  wr_data_rom[16298]='h00000000;
    rd_cycle[16299] = 1'b1;  wr_cycle[16299] = 1'b0;  addr_rom[16299]='h00001200;  wr_data_rom[16299]='h00000000;
    rd_cycle[16300] = 1'b1;  wr_cycle[16300] = 1'b0;  addr_rom[16300]='h00000210;  wr_data_rom[16300]='h00000000;
    rd_cycle[16301] = 1'b1;  wr_cycle[16301] = 1'b0;  addr_rom[16301]='h00000624;  wr_data_rom[16301]='h00000000;
    rd_cycle[16302] = 1'b1;  wr_cycle[16302] = 1'b0;  addr_rom[16302]='h000020c8;  wr_data_rom[16302]='h00000000;
    rd_cycle[16303] = 1'b0;  wr_cycle[16303] = 1'b1;  addr_rom[16303]='h000021c8;  wr_data_rom[16303]='h0000291d;
    rd_cycle[16304] = 1'b1;  wr_cycle[16304] = 1'b0;  addr_rom[16304]='h000020b8;  wr_data_rom[16304]='h00000000;
    rd_cycle[16305] = 1'b0;  wr_cycle[16305] = 1'b1;  addr_rom[16305]='h00002cac;  wr_data_rom[16305]='h00002eaf;
    rd_cycle[16306] = 1'b1;  wr_cycle[16306] = 1'b0;  addr_rom[16306]='h000012e8;  wr_data_rom[16306]='h00000000;
    rd_cycle[16307] = 1'b0;  wr_cycle[16307] = 1'b1;  addr_rom[16307]='h0000146c;  wr_data_rom[16307]='h00000951;
    rd_cycle[16308] = 1'b0;  wr_cycle[16308] = 1'b1;  addr_rom[16308]='h00000e30;  wr_data_rom[16308]='h00003c06;
    rd_cycle[16309] = 1'b1;  wr_cycle[16309] = 1'b0;  addr_rom[16309]='h00003830;  wr_data_rom[16309]='h00000000;
    rd_cycle[16310] = 1'b0;  wr_cycle[16310] = 1'b1;  addr_rom[16310]='h00002104;  wr_data_rom[16310]='h00001616;
    rd_cycle[16311] = 1'b0;  wr_cycle[16311] = 1'b1;  addr_rom[16311]='h00002a24;  wr_data_rom[16311]='h000020f7;
    rd_cycle[16312] = 1'b1;  wr_cycle[16312] = 1'b0;  addr_rom[16312]='h0000190c;  wr_data_rom[16312]='h00000000;
    rd_cycle[16313] = 1'b0;  wr_cycle[16313] = 1'b1;  addr_rom[16313]='h00001f40;  wr_data_rom[16313]='h000035cb;
    rd_cycle[16314] = 1'b0;  wr_cycle[16314] = 1'b1;  addr_rom[16314]='h000019dc;  wr_data_rom[16314]='h0000095f;
    rd_cycle[16315] = 1'b0;  wr_cycle[16315] = 1'b1;  addr_rom[16315]='h00002fc0;  wr_data_rom[16315]='h000001b2;
    rd_cycle[16316] = 1'b0;  wr_cycle[16316] = 1'b1;  addr_rom[16316]='h000039a8;  wr_data_rom[16316]='h00000621;
    rd_cycle[16317] = 1'b0;  wr_cycle[16317] = 1'b1;  addr_rom[16317]='h00001068;  wr_data_rom[16317]='h00001a5c;
    rd_cycle[16318] = 1'b0;  wr_cycle[16318] = 1'b1;  addr_rom[16318]='h00002534;  wr_data_rom[16318]='h00000aa8;
    rd_cycle[16319] = 1'b0;  wr_cycle[16319] = 1'b1;  addr_rom[16319]='h00003168;  wr_data_rom[16319]='h000006f2;
    rd_cycle[16320] = 1'b1;  wr_cycle[16320] = 1'b0;  addr_rom[16320]='h00001914;  wr_data_rom[16320]='h00000000;
    rd_cycle[16321] = 1'b0;  wr_cycle[16321] = 1'b1;  addr_rom[16321]='h000034f4;  wr_data_rom[16321]='h00001dec;
    rd_cycle[16322] = 1'b1;  wr_cycle[16322] = 1'b0;  addr_rom[16322]='h0000257c;  wr_data_rom[16322]='h00000000;
    rd_cycle[16323] = 1'b0;  wr_cycle[16323] = 1'b1;  addr_rom[16323]='h00001aa4;  wr_data_rom[16323]='h00001db5;
    rd_cycle[16324] = 1'b0;  wr_cycle[16324] = 1'b1;  addr_rom[16324]='h000007bc;  wr_data_rom[16324]='h000010b7;
    rd_cycle[16325] = 1'b0;  wr_cycle[16325] = 1'b1;  addr_rom[16325]='h00000dd4;  wr_data_rom[16325]='h00002cad;
    rd_cycle[16326] = 1'b0;  wr_cycle[16326] = 1'b1;  addr_rom[16326]='h000019e8;  wr_data_rom[16326]='h00002526;
    rd_cycle[16327] = 1'b1;  wr_cycle[16327] = 1'b0;  addr_rom[16327]='h0000136c;  wr_data_rom[16327]='h00000000;
    rd_cycle[16328] = 1'b0;  wr_cycle[16328] = 1'b1;  addr_rom[16328]='h00003ac0;  wr_data_rom[16328]='h000020df;
    rd_cycle[16329] = 1'b1;  wr_cycle[16329] = 1'b0;  addr_rom[16329]='h00000510;  wr_data_rom[16329]='h00000000;
    rd_cycle[16330] = 1'b0;  wr_cycle[16330] = 1'b1;  addr_rom[16330]='h00000a68;  wr_data_rom[16330]='h00000942;
    rd_cycle[16331] = 1'b1;  wr_cycle[16331] = 1'b0;  addr_rom[16331]='h00000fac;  wr_data_rom[16331]='h00000000;
    rd_cycle[16332] = 1'b1;  wr_cycle[16332] = 1'b0;  addr_rom[16332]='h0000271c;  wr_data_rom[16332]='h00000000;
    rd_cycle[16333] = 1'b1;  wr_cycle[16333] = 1'b0;  addr_rom[16333]='h000010b0;  wr_data_rom[16333]='h00000000;
    rd_cycle[16334] = 1'b0;  wr_cycle[16334] = 1'b1;  addr_rom[16334]='h00001b88;  wr_data_rom[16334]='h00002e88;
    rd_cycle[16335] = 1'b1;  wr_cycle[16335] = 1'b0;  addr_rom[16335]='h000003e4;  wr_data_rom[16335]='h00000000;
    rd_cycle[16336] = 1'b1;  wr_cycle[16336] = 1'b0;  addr_rom[16336]='h00002744;  wr_data_rom[16336]='h00000000;
    rd_cycle[16337] = 1'b0;  wr_cycle[16337] = 1'b1;  addr_rom[16337]='h00000440;  wr_data_rom[16337]='h000021c4;
    rd_cycle[16338] = 1'b1;  wr_cycle[16338] = 1'b0;  addr_rom[16338]='h00001134;  wr_data_rom[16338]='h00000000;
    rd_cycle[16339] = 1'b0;  wr_cycle[16339] = 1'b1;  addr_rom[16339]='h00002268;  wr_data_rom[16339]='h0000335d;
    rd_cycle[16340] = 1'b0;  wr_cycle[16340] = 1'b1;  addr_rom[16340]='h00001330;  wr_data_rom[16340]='h000005a8;
    rd_cycle[16341] = 1'b0;  wr_cycle[16341] = 1'b1;  addr_rom[16341]='h00000a2c;  wr_data_rom[16341]='h00002124;
    rd_cycle[16342] = 1'b1;  wr_cycle[16342] = 1'b0;  addr_rom[16342]='h00000690;  wr_data_rom[16342]='h00000000;
    rd_cycle[16343] = 1'b1;  wr_cycle[16343] = 1'b0;  addr_rom[16343]='h00002728;  wr_data_rom[16343]='h00000000;
    rd_cycle[16344] = 1'b0;  wr_cycle[16344] = 1'b1;  addr_rom[16344]='h00002430;  wr_data_rom[16344]='h000035d3;
    rd_cycle[16345] = 1'b0;  wr_cycle[16345] = 1'b1;  addr_rom[16345]='h00003150;  wr_data_rom[16345]='h00002996;
    rd_cycle[16346] = 1'b1;  wr_cycle[16346] = 1'b0;  addr_rom[16346]='h00000e58;  wr_data_rom[16346]='h00000000;
    rd_cycle[16347] = 1'b0;  wr_cycle[16347] = 1'b1;  addr_rom[16347]='h00003d38;  wr_data_rom[16347]='h00000273;
    rd_cycle[16348] = 1'b1;  wr_cycle[16348] = 1'b0;  addr_rom[16348]='h00000808;  wr_data_rom[16348]='h00000000;
    rd_cycle[16349] = 1'b1;  wr_cycle[16349] = 1'b0;  addr_rom[16349]='h00001940;  wr_data_rom[16349]='h00000000;
    rd_cycle[16350] = 1'b0;  wr_cycle[16350] = 1'b1;  addr_rom[16350]='h00002404;  wr_data_rom[16350]='h0000282c;
    rd_cycle[16351] = 1'b1;  wr_cycle[16351] = 1'b0;  addr_rom[16351]='h0000376c;  wr_data_rom[16351]='h00000000;
    rd_cycle[16352] = 1'b0;  wr_cycle[16352] = 1'b1;  addr_rom[16352]='h00001328;  wr_data_rom[16352]='h0000296b;
    rd_cycle[16353] = 1'b1;  wr_cycle[16353] = 1'b0;  addr_rom[16353]='h000021cc;  wr_data_rom[16353]='h00000000;
    rd_cycle[16354] = 1'b1;  wr_cycle[16354] = 1'b0;  addr_rom[16354]='h00000dc0;  wr_data_rom[16354]='h00000000;
    rd_cycle[16355] = 1'b1;  wr_cycle[16355] = 1'b0;  addr_rom[16355]='h00002624;  wr_data_rom[16355]='h00000000;
    rd_cycle[16356] = 1'b0;  wr_cycle[16356] = 1'b1;  addr_rom[16356]='h00000584;  wr_data_rom[16356]='h00000931;
    rd_cycle[16357] = 1'b1;  wr_cycle[16357] = 1'b0;  addr_rom[16357]='h000016f0;  wr_data_rom[16357]='h00000000;
    rd_cycle[16358] = 1'b1;  wr_cycle[16358] = 1'b0;  addr_rom[16358]='h00001cfc;  wr_data_rom[16358]='h00000000;
    rd_cycle[16359] = 1'b1;  wr_cycle[16359] = 1'b0;  addr_rom[16359]='h00001644;  wr_data_rom[16359]='h00000000;
    rd_cycle[16360] = 1'b1;  wr_cycle[16360] = 1'b0;  addr_rom[16360]='h00000464;  wr_data_rom[16360]='h00000000;
    rd_cycle[16361] = 1'b0;  wr_cycle[16361] = 1'b1;  addr_rom[16361]='h00002958;  wr_data_rom[16361]='h00002bcd;
    rd_cycle[16362] = 1'b1;  wr_cycle[16362] = 1'b0;  addr_rom[16362]='h0000223c;  wr_data_rom[16362]='h00000000;
    rd_cycle[16363] = 1'b1;  wr_cycle[16363] = 1'b0;  addr_rom[16363]='h000008fc;  wr_data_rom[16363]='h00000000;
    rd_cycle[16364] = 1'b0;  wr_cycle[16364] = 1'b1;  addr_rom[16364]='h00001acc;  wr_data_rom[16364]='h0000232e;
    rd_cycle[16365] = 1'b1;  wr_cycle[16365] = 1'b0;  addr_rom[16365]='h00001be4;  wr_data_rom[16365]='h00000000;
    rd_cycle[16366] = 1'b0;  wr_cycle[16366] = 1'b1;  addr_rom[16366]='h00001014;  wr_data_rom[16366]='h00001b8d;
    rd_cycle[16367] = 1'b0;  wr_cycle[16367] = 1'b1;  addr_rom[16367]='h00000010;  wr_data_rom[16367]='h00002082;
    rd_cycle[16368] = 1'b1;  wr_cycle[16368] = 1'b0;  addr_rom[16368]='h00002a2c;  wr_data_rom[16368]='h00000000;
    rd_cycle[16369] = 1'b1;  wr_cycle[16369] = 1'b0;  addr_rom[16369]='h00001fb0;  wr_data_rom[16369]='h00000000;
    rd_cycle[16370] = 1'b1;  wr_cycle[16370] = 1'b0;  addr_rom[16370]='h000028dc;  wr_data_rom[16370]='h00000000;
    rd_cycle[16371] = 1'b0;  wr_cycle[16371] = 1'b1;  addr_rom[16371]='h00001700;  wr_data_rom[16371]='h000030e1;
    rd_cycle[16372] = 1'b0;  wr_cycle[16372] = 1'b1;  addr_rom[16372]='h000029d4;  wr_data_rom[16372]='h00002fef;
    rd_cycle[16373] = 1'b1;  wr_cycle[16373] = 1'b0;  addr_rom[16373]='h00000200;  wr_data_rom[16373]='h00000000;
    rd_cycle[16374] = 1'b0;  wr_cycle[16374] = 1'b1;  addr_rom[16374]='h00002b9c;  wr_data_rom[16374]='h000021a5;
    rd_cycle[16375] = 1'b0;  wr_cycle[16375] = 1'b1;  addr_rom[16375]='h00000840;  wr_data_rom[16375]='h0000298b;
    rd_cycle[16376] = 1'b0;  wr_cycle[16376] = 1'b1;  addr_rom[16376]='h000019b4;  wr_data_rom[16376]='h00002840;
    rd_cycle[16377] = 1'b0;  wr_cycle[16377] = 1'b1;  addr_rom[16377]='h00003e48;  wr_data_rom[16377]='h00001e1b;
    rd_cycle[16378] = 1'b0;  wr_cycle[16378] = 1'b1;  addr_rom[16378]='h000008e0;  wr_data_rom[16378]='h000032d4;
    rd_cycle[16379] = 1'b0;  wr_cycle[16379] = 1'b1;  addr_rom[16379]='h00001f5c;  wr_data_rom[16379]='h00001236;
    rd_cycle[16380] = 1'b0;  wr_cycle[16380] = 1'b1;  addr_rom[16380]='h00001a10;  wr_data_rom[16380]='h00001d05;
    rd_cycle[16381] = 1'b0;  wr_cycle[16381] = 1'b1;  addr_rom[16381]='h0000069c;  wr_data_rom[16381]='h00003257;
    rd_cycle[16382] = 1'b0;  wr_cycle[16382] = 1'b1;  addr_rom[16382]='h00003180;  wr_data_rom[16382]='h00001370;
    rd_cycle[16383] = 1'b0;  wr_cycle[16383] = 1'b1;  addr_rom[16383]='h00003268;  wr_data_rom[16383]='h000001ec;
    // 4096 silence cycles
    rd_cycle[16384] = 1'b0;  wr_cycle[16384] = 1'b0;  addr_rom[16384]='h00000000;  wr_data_rom[16384]='h00000000;
    rd_cycle[16385] = 1'b0;  wr_cycle[16385] = 1'b0;  addr_rom[16385]='h00000000;  wr_data_rom[16385]='h00000000;
    rd_cycle[16386] = 1'b0;  wr_cycle[16386] = 1'b0;  addr_rom[16386]='h00000000;  wr_data_rom[16386]='h00000000;
    rd_cycle[16387] = 1'b0;  wr_cycle[16387] = 1'b0;  addr_rom[16387]='h00000000;  wr_data_rom[16387]='h00000000;
    rd_cycle[16388] = 1'b0;  wr_cycle[16388] = 1'b0;  addr_rom[16388]='h00000000;  wr_data_rom[16388]='h00000000;
    rd_cycle[16389] = 1'b0;  wr_cycle[16389] = 1'b0;  addr_rom[16389]='h00000000;  wr_data_rom[16389]='h00000000;
    rd_cycle[16390] = 1'b0;  wr_cycle[16390] = 1'b0;  addr_rom[16390]='h00000000;  wr_data_rom[16390]='h00000000;
    rd_cycle[16391] = 1'b0;  wr_cycle[16391] = 1'b0;  addr_rom[16391]='h00000000;  wr_data_rom[16391]='h00000000;
    rd_cycle[16392] = 1'b0;  wr_cycle[16392] = 1'b0;  addr_rom[16392]='h00000000;  wr_data_rom[16392]='h00000000;
    rd_cycle[16393] = 1'b0;  wr_cycle[16393] = 1'b0;  addr_rom[16393]='h00000000;  wr_data_rom[16393]='h00000000;
    rd_cycle[16394] = 1'b0;  wr_cycle[16394] = 1'b0;  addr_rom[16394]='h00000000;  wr_data_rom[16394]='h00000000;
    rd_cycle[16395] = 1'b0;  wr_cycle[16395] = 1'b0;  addr_rom[16395]='h00000000;  wr_data_rom[16395]='h00000000;
    rd_cycle[16396] = 1'b0;  wr_cycle[16396] = 1'b0;  addr_rom[16396]='h00000000;  wr_data_rom[16396]='h00000000;
    rd_cycle[16397] = 1'b0;  wr_cycle[16397] = 1'b0;  addr_rom[16397]='h00000000;  wr_data_rom[16397]='h00000000;
    rd_cycle[16398] = 1'b0;  wr_cycle[16398] = 1'b0;  addr_rom[16398]='h00000000;  wr_data_rom[16398]='h00000000;
    rd_cycle[16399] = 1'b0;  wr_cycle[16399] = 1'b0;  addr_rom[16399]='h00000000;  wr_data_rom[16399]='h00000000;
    rd_cycle[16400] = 1'b0;  wr_cycle[16400] = 1'b0;  addr_rom[16400]='h00000000;  wr_data_rom[16400]='h00000000;
    rd_cycle[16401] = 1'b0;  wr_cycle[16401] = 1'b0;  addr_rom[16401]='h00000000;  wr_data_rom[16401]='h00000000;
    rd_cycle[16402] = 1'b0;  wr_cycle[16402] = 1'b0;  addr_rom[16402]='h00000000;  wr_data_rom[16402]='h00000000;
    rd_cycle[16403] = 1'b0;  wr_cycle[16403] = 1'b0;  addr_rom[16403]='h00000000;  wr_data_rom[16403]='h00000000;
    rd_cycle[16404] = 1'b0;  wr_cycle[16404] = 1'b0;  addr_rom[16404]='h00000000;  wr_data_rom[16404]='h00000000;
    rd_cycle[16405] = 1'b0;  wr_cycle[16405] = 1'b0;  addr_rom[16405]='h00000000;  wr_data_rom[16405]='h00000000;
    rd_cycle[16406] = 1'b0;  wr_cycle[16406] = 1'b0;  addr_rom[16406]='h00000000;  wr_data_rom[16406]='h00000000;
    rd_cycle[16407] = 1'b0;  wr_cycle[16407] = 1'b0;  addr_rom[16407]='h00000000;  wr_data_rom[16407]='h00000000;
    rd_cycle[16408] = 1'b0;  wr_cycle[16408] = 1'b0;  addr_rom[16408]='h00000000;  wr_data_rom[16408]='h00000000;
    rd_cycle[16409] = 1'b0;  wr_cycle[16409] = 1'b0;  addr_rom[16409]='h00000000;  wr_data_rom[16409]='h00000000;
    rd_cycle[16410] = 1'b0;  wr_cycle[16410] = 1'b0;  addr_rom[16410]='h00000000;  wr_data_rom[16410]='h00000000;
    rd_cycle[16411] = 1'b0;  wr_cycle[16411] = 1'b0;  addr_rom[16411]='h00000000;  wr_data_rom[16411]='h00000000;
    rd_cycle[16412] = 1'b0;  wr_cycle[16412] = 1'b0;  addr_rom[16412]='h00000000;  wr_data_rom[16412]='h00000000;
    rd_cycle[16413] = 1'b0;  wr_cycle[16413] = 1'b0;  addr_rom[16413]='h00000000;  wr_data_rom[16413]='h00000000;
    rd_cycle[16414] = 1'b0;  wr_cycle[16414] = 1'b0;  addr_rom[16414]='h00000000;  wr_data_rom[16414]='h00000000;
    rd_cycle[16415] = 1'b0;  wr_cycle[16415] = 1'b0;  addr_rom[16415]='h00000000;  wr_data_rom[16415]='h00000000;
    rd_cycle[16416] = 1'b0;  wr_cycle[16416] = 1'b0;  addr_rom[16416]='h00000000;  wr_data_rom[16416]='h00000000;
    rd_cycle[16417] = 1'b0;  wr_cycle[16417] = 1'b0;  addr_rom[16417]='h00000000;  wr_data_rom[16417]='h00000000;
    rd_cycle[16418] = 1'b0;  wr_cycle[16418] = 1'b0;  addr_rom[16418]='h00000000;  wr_data_rom[16418]='h00000000;
    rd_cycle[16419] = 1'b0;  wr_cycle[16419] = 1'b0;  addr_rom[16419]='h00000000;  wr_data_rom[16419]='h00000000;
    rd_cycle[16420] = 1'b0;  wr_cycle[16420] = 1'b0;  addr_rom[16420]='h00000000;  wr_data_rom[16420]='h00000000;
    rd_cycle[16421] = 1'b0;  wr_cycle[16421] = 1'b0;  addr_rom[16421]='h00000000;  wr_data_rom[16421]='h00000000;
    rd_cycle[16422] = 1'b0;  wr_cycle[16422] = 1'b0;  addr_rom[16422]='h00000000;  wr_data_rom[16422]='h00000000;
    rd_cycle[16423] = 1'b0;  wr_cycle[16423] = 1'b0;  addr_rom[16423]='h00000000;  wr_data_rom[16423]='h00000000;
    rd_cycle[16424] = 1'b0;  wr_cycle[16424] = 1'b0;  addr_rom[16424]='h00000000;  wr_data_rom[16424]='h00000000;
    rd_cycle[16425] = 1'b0;  wr_cycle[16425] = 1'b0;  addr_rom[16425]='h00000000;  wr_data_rom[16425]='h00000000;
    rd_cycle[16426] = 1'b0;  wr_cycle[16426] = 1'b0;  addr_rom[16426]='h00000000;  wr_data_rom[16426]='h00000000;
    rd_cycle[16427] = 1'b0;  wr_cycle[16427] = 1'b0;  addr_rom[16427]='h00000000;  wr_data_rom[16427]='h00000000;
    rd_cycle[16428] = 1'b0;  wr_cycle[16428] = 1'b0;  addr_rom[16428]='h00000000;  wr_data_rom[16428]='h00000000;
    rd_cycle[16429] = 1'b0;  wr_cycle[16429] = 1'b0;  addr_rom[16429]='h00000000;  wr_data_rom[16429]='h00000000;
    rd_cycle[16430] = 1'b0;  wr_cycle[16430] = 1'b0;  addr_rom[16430]='h00000000;  wr_data_rom[16430]='h00000000;
    rd_cycle[16431] = 1'b0;  wr_cycle[16431] = 1'b0;  addr_rom[16431]='h00000000;  wr_data_rom[16431]='h00000000;
    rd_cycle[16432] = 1'b0;  wr_cycle[16432] = 1'b0;  addr_rom[16432]='h00000000;  wr_data_rom[16432]='h00000000;
    rd_cycle[16433] = 1'b0;  wr_cycle[16433] = 1'b0;  addr_rom[16433]='h00000000;  wr_data_rom[16433]='h00000000;
    rd_cycle[16434] = 1'b0;  wr_cycle[16434] = 1'b0;  addr_rom[16434]='h00000000;  wr_data_rom[16434]='h00000000;
    rd_cycle[16435] = 1'b0;  wr_cycle[16435] = 1'b0;  addr_rom[16435]='h00000000;  wr_data_rom[16435]='h00000000;
    rd_cycle[16436] = 1'b0;  wr_cycle[16436] = 1'b0;  addr_rom[16436]='h00000000;  wr_data_rom[16436]='h00000000;
    rd_cycle[16437] = 1'b0;  wr_cycle[16437] = 1'b0;  addr_rom[16437]='h00000000;  wr_data_rom[16437]='h00000000;
    rd_cycle[16438] = 1'b0;  wr_cycle[16438] = 1'b0;  addr_rom[16438]='h00000000;  wr_data_rom[16438]='h00000000;
    rd_cycle[16439] = 1'b0;  wr_cycle[16439] = 1'b0;  addr_rom[16439]='h00000000;  wr_data_rom[16439]='h00000000;
    rd_cycle[16440] = 1'b0;  wr_cycle[16440] = 1'b0;  addr_rom[16440]='h00000000;  wr_data_rom[16440]='h00000000;
    rd_cycle[16441] = 1'b0;  wr_cycle[16441] = 1'b0;  addr_rom[16441]='h00000000;  wr_data_rom[16441]='h00000000;
    rd_cycle[16442] = 1'b0;  wr_cycle[16442] = 1'b0;  addr_rom[16442]='h00000000;  wr_data_rom[16442]='h00000000;
    rd_cycle[16443] = 1'b0;  wr_cycle[16443] = 1'b0;  addr_rom[16443]='h00000000;  wr_data_rom[16443]='h00000000;
    rd_cycle[16444] = 1'b0;  wr_cycle[16444] = 1'b0;  addr_rom[16444]='h00000000;  wr_data_rom[16444]='h00000000;
    rd_cycle[16445] = 1'b0;  wr_cycle[16445] = 1'b0;  addr_rom[16445]='h00000000;  wr_data_rom[16445]='h00000000;
    rd_cycle[16446] = 1'b0;  wr_cycle[16446] = 1'b0;  addr_rom[16446]='h00000000;  wr_data_rom[16446]='h00000000;
    rd_cycle[16447] = 1'b0;  wr_cycle[16447] = 1'b0;  addr_rom[16447]='h00000000;  wr_data_rom[16447]='h00000000;
    rd_cycle[16448] = 1'b0;  wr_cycle[16448] = 1'b0;  addr_rom[16448]='h00000000;  wr_data_rom[16448]='h00000000;
    rd_cycle[16449] = 1'b0;  wr_cycle[16449] = 1'b0;  addr_rom[16449]='h00000000;  wr_data_rom[16449]='h00000000;
    rd_cycle[16450] = 1'b0;  wr_cycle[16450] = 1'b0;  addr_rom[16450]='h00000000;  wr_data_rom[16450]='h00000000;
    rd_cycle[16451] = 1'b0;  wr_cycle[16451] = 1'b0;  addr_rom[16451]='h00000000;  wr_data_rom[16451]='h00000000;
    rd_cycle[16452] = 1'b0;  wr_cycle[16452] = 1'b0;  addr_rom[16452]='h00000000;  wr_data_rom[16452]='h00000000;
    rd_cycle[16453] = 1'b0;  wr_cycle[16453] = 1'b0;  addr_rom[16453]='h00000000;  wr_data_rom[16453]='h00000000;
    rd_cycle[16454] = 1'b0;  wr_cycle[16454] = 1'b0;  addr_rom[16454]='h00000000;  wr_data_rom[16454]='h00000000;
    rd_cycle[16455] = 1'b0;  wr_cycle[16455] = 1'b0;  addr_rom[16455]='h00000000;  wr_data_rom[16455]='h00000000;
    rd_cycle[16456] = 1'b0;  wr_cycle[16456] = 1'b0;  addr_rom[16456]='h00000000;  wr_data_rom[16456]='h00000000;
    rd_cycle[16457] = 1'b0;  wr_cycle[16457] = 1'b0;  addr_rom[16457]='h00000000;  wr_data_rom[16457]='h00000000;
    rd_cycle[16458] = 1'b0;  wr_cycle[16458] = 1'b0;  addr_rom[16458]='h00000000;  wr_data_rom[16458]='h00000000;
    rd_cycle[16459] = 1'b0;  wr_cycle[16459] = 1'b0;  addr_rom[16459]='h00000000;  wr_data_rom[16459]='h00000000;
    rd_cycle[16460] = 1'b0;  wr_cycle[16460] = 1'b0;  addr_rom[16460]='h00000000;  wr_data_rom[16460]='h00000000;
    rd_cycle[16461] = 1'b0;  wr_cycle[16461] = 1'b0;  addr_rom[16461]='h00000000;  wr_data_rom[16461]='h00000000;
    rd_cycle[16462] = 1'b0;  wr_cycle[16462] = 1'b0;  addr_rom[16462]='h00000000;  wr_data_rom[16462]='h00000000;
    rd_cycle[16463] = 1'b0;  wr_cycle[16463] = 1'b0;  addr_rom[16463]='h00000000;  wr_data_rom[16463]='h00000000;
    rd_cycle[16464] = 1'b0;  wr_cycle[16464] = 1'b0;  addr_rom[16464]='h00000000;  wr_data_rom[16464]='h00000000;
    rd_cycle[16465] = 1'b0;  wr_cycle[16465] = 1'b0;  addr_rom[16465]='h00000000;  wr_data_rom[16465]='h00000000;
    rd_cycle[16466] = 1'b0;  wr_cycle[16466] = 1'b0;  addr_rom[16466]='h00000000;  wr_data_rom[16466]='h00000000;
    rd_cycle[16467] = 1'b0;  wr_cycle[16467] = 1'b0;  addr_rom[16467]='h00000000;  wr_data_rom[16467]='h00000000;
    rd_cycle[16468] = 1'b0;  wr_cycle[16468] = 1'b0;  addr_rom[16468]='h00000000;  wr_data_rom[16468]='h00000000;
    rd_cycle[16469] = 1'b0;  wr_cycle[16469] = 1'b0;  addr_rom[16469]='h00000000;  wr_data_rom[16469]='h00000000;
    rd_cycle[16470] = 1'b0;  wr_cycle[16470] = 1'b0;  addr_rom[16470]='h00000000;  wr_data_rom[16470]='h00000000;
    rd_cycle[16471] = 1'b0;  wr_cycle[16471] = 1'b0;  addr_rom[16471]='h00000000;  wr_data_rom[16471]='h00000000;
    rd_cycle[16472] = 1'b0;  wr_cycle[16472] = 1'b0;  addr_rom[16472]='h00000000;  wr_data_rom[16472]='h00000000;
    rd_cycle[16473] = 1'b0;  wr_cycle[16473] = 1'b0;  addr_rom[16473]='h00000000;  wr_data_rom[16473]='h00000000;
    rd_cycle[16474] = 1'b0;  wr_cycle[16474] = 1'b0;  addr_rom[16474]='h00000000;  wr_data_rom[16474]='h00000000;
    rd_cycle[16475] = 1'b0;  wr_cycle[16475] = 1'b0;  addr_rom[16475]='h00000000;  wr_data_rom[16475]='h00000000;
    rd_cycle[16476] = 1'b0;  wr_cycle[16476] = 1'b0;  addr_rom[16476]='h00000000;  wr_data_rom[16476]='h00000000;
    rd_cycle[16477] = 1'b0;  wr_cycle[16477] = 1'b0;  addr_rom[16477]='h00000000;  wr_data_rom[16477]='h00000000;
    rd_cycle[16478] = 1'b0;  wr_cycle[16478] = 1'b0;  addr_rom[16478]='h00000000;  wr_data_rom[16478]='h00000000;
    rd_cycle[16479] = 1'b0;  wr_cycle[16479] = 1'b0;  addr_rom[16479]='h00000000;  wr_data_rom[16479]='h00000000;
    rd_cycle[16480] = 1'b0;  wr_cycle[16480] = 1'b0;  addr_rom[16480]='h00000000;  wr_data_rom[16480]='h00000000;
    rd_cycle[16481] = 1'b0;  wr_cycle[16481] = 1'b0;  addr_rom[16481]='h00000000;  wr_data_rom[16481]='h00000000;
    rd_cycle[16482] = 1'b0;  wr_cycle[16482] = 1'b0;  addr_rom[16482]='h00000000;  wr_data_rom[16482]='h00000000;
    rd_cycle[16483] = 1'b0;  wr_cycle[16483] = 1'b0;  addr_rom[16483]='h00000000;  wr_data_rom[16483]='h00000000;
    rd_cycle[16484] = 1'b0;  wr_cycle[16484] = 1'b0;  addr_rom[16484]='h00000000;  wr_data_rom[16484]='h00000000;
    rd_cycle[16485] = 1'b0;  wr_cycle[16485] = 1'b0;  addr_rom[16485]='h00000000;  wr_data_rom[16485]='h00000000;
    rd_cycle[16486] = 1'b0;  wr_cycle[16486] = 1'b0;  addr_rom[16486]='h00000000;  wr_data_rom[16486]='h00000000;
    rd_cycle[16487] = 1'b0;  wr_cycle[16487] = 1'b0;  addr_rom[16487]='h00000000;  wr_data_rom[16487]='h00000000;
    rd_cycle[16488] = 1'b0;  wr_cycle[16488] = 1'b0;  addr_rom[16488]='h00000000;  wr_data_rom[16488]='h00000000;
    rd_cycle[16489] = 1'b0;  wr_cycle[16489] = 1'b0;  addr_rom[16489]='h00000000;  wr_data_rom[16489]='h00000000;
    rd_cycle[16490] = 1'b0;  wr_cycle[16490] = 1'b0;  addr_rom[16490]='h00000000;  wr_data_rom[16490]='h00000000;
    rd_cycle[16491] = 1'b0;  wr_cycle[16491] = 1'b0;  addr_rom[16491]='h00000000;  wr_data_rom[16491]='h00000000;
    rd_cycle[16492] = 1'b0;  wr_cycle[16492] = 1'b0;  addr_rom[16492]='h00000000;  wr_data_rom[16492]='h00000000;
    rd_cycle[16493] = 1'b0;  wr_cycle[16493] = 1'b0;  addr_rom[16493]='h00000000;  wr_data_rom[16493]='h00000000;
    rd_cycle[16494] = 1'b0;  wr_cycle[16494] = 1'b0;  addr_rom[16494]='h00000000;  wr_data_rom[16494]='h00000000;
    rd_cycle[16495] = 1'b0;  wr_cycle[16495] = 1'b0;  addr_rom[16495]='h00000000;  wr_data_rom[16495]='h00000000;
    rd_cycle[16496] = 1'b0;  wr_cycle[16496] = 1'b0;  addr_rom[16496]='h00000000;  wr_data_rom[16496]='h00000000;
    rd_cycle[16497] = 1'b0;  wr_cycle[16497] = 1'b0;  addr_rom[16497]='h00000000;  wr_data_rom[16497]='h00000000;
    rd_cycle[16498] = 1'b0;  wr_cycle[16498] = 1'b0;  addr_rom[16498]='h00000000;  wr_data_rom[16498]='h00000000;
    rd_cycle[16499] = 1'b0;  wr_cycle[16499] = 1'b0;  addr_rom[16499]='h00000000;  wr_data_rom[16499]='h00000000;
    rd_cycle[16500] = 1'b0;  wr_cycle[16500] = 1'b0;  addr_rom[16500]='h00000000;  wr_data_rom[16500]='h00000000;
    rd_cycle[16501] = 1'b0;  wr_cycle[16501] = 1'b0;  addr_rom[16501]='h00000000;  wr_data_rom[16501]='h00000000;
    rd_cycle[16502] = 1'b0;  wr_cycle[16502] = 1'b0;  addr_rom[16502]='h00000000;  wr_data_rom[16502]='h00000000;
    rd_cycle[16503] = 1'b0;  wr_cycle[16503] = 1'b0;  addr_rom[16503]='h00000000;  wr_data_rom[16503]='h00000000;
    rd_cycle[16504] = 1'b0;  wr_cycle[16504] = 1'b0;  addr_rom[16504]='h00000000;  wr_data_rom[16504]='h00000000;
    rd_cycle[16505] = 1'b0;  wr_cycle[16505] = 1'b0;  addr_rom[16505]='h00000000;  wr_data_rom[16505]='h00000000;
    rd_cycle[16506] = 1'b0;  wr_cycle[16506] = 1'b0;  addr_rom[16506]='h00000000;  wr_data_rom[16506]='h00000000;
    rd_cycle[16507] = 1'b0;  wr_cycle[16507] = 1'b0;  addr_rom[16507]='h00000000;  wr_data_rom[16507]='h00000000;
    rd_cycle[16508] = 1'b0;  wr_cycle[16508] = 1'b0;  addr_rom[16508]='h00000000;  wr_data_rom[16508]='h00000000;
    rd_cycle[16509] = 1'b0;  wr_cycle[16509] = 1'b0;  addr_rom[16509]='h00000000;  wr_data_rom[16509]='h00000000;
    rd_cycle[16510] = 1'b0;  wr_cycle[16510] = 1'b0;  addr_rom[16510]='h00000000;  wr_data_rom[16510]='h00000000;
    rd_cycle[16511] = 1'b0;  wr_cycle[16511] = 1'b0;  addr_rom[16511]='h00000000;  wr_data_rom[16511]='h00000000;
    rd_cycle[16512] = 1'b0;  wr_cycle[16512] = 1'b0;  addr_rom[16512]='h00000000;  wr_data_rom[16512]='h00000000;
    rd_cycle[16513] = 1'b0;  wr_cycle[16513] = 1'b0;  addr_rom[16513]='h00000000;  wr_data_rom[16513]='h00000000;
    rd_cycle[16514] = 1'b0;  wr_cycle[16514] = 1'b0;  addr_rom[16514]='h00000000;  wr_data_rom[16514]='h00000000;
    rd_cycle[16515] = 1'b0;  wr_cycle[16515] = 1'b0;  addr_rom[16515]='h00000000;  wr_data_rom[16515]='h00000000;
    rd_cycle[16516] = 1'b0;  wr_cycle[16516] = 1'b0;  addr_rom[16516]='h00000000;  wr_data_rom[16516]='h00000000;
    rd_cycle[16517] = 1'b0;  wr_cycle[16517] = 1'b0;  addr_rom[16517]='h00000000;  wr_data_rom[16517]='h00000000;
    rd_cycle[16518] = 1'b0;  wr_cycle[16518] = 1'b0;  addr_rom[16518]='h00000000;  wr_data_rom[16518]='h00000000;
    rd_cycle[16519] = 1'b0;  wr_cycle[16519] = 1'b0;  addr_rom[16519]='h00000000;  wr_data_rom[16519]='h00000000;
    rd_cycle[16520] = 1'b0;  wr_cycle[16520] = 1'b0;  addr_rom[16520]='h00000000;  wr_data_rom[16520]='h00000000;
    rd_cycle[16521] = 1'b0;  wr_cycle[16521] = 1'b0;  addr_rom[16521]='h00000000;  wr_data_rom[16521]='h00000000;
    rd_cycle[16522] = 1'b0;  wr_cycle[16522] = 1'b0;  addr_rom[16522]='h00000000;  wr_data_rom[16522]='h00000000;
    rd_cycle[16523] = 1'b0;  wr_cycle[16523] = 1'b0;  addr_rom[16523]='h00000000;  wr_data_rom[16523]='h00000000;
    rd_cycle[16524] = 1'b0;  wr_cycle[16524] = 1'b0;  addr_rom[16524]='h00000000;  wr_data_rom[16524]='h00000000;
    rd_cycle[16525] = 1'b0;  wr_cycle[16525] = 1'b0;  addr_rom[16525]='h00000000;  wr_data_rom[16525]='h00000000;
    rd_cycle[16526] = 1'b0;  wr_cycle[16526] = 1'b0;  addr_rom[16526]='h00000000;  wr_data_rom[16526]='h00000000;
    rd_cycle[16527] = 1'b0;  wr_cycle[16527] = 1'b0;  addr_rom[16527]='h00000000;  wr_data_rom[16527]='h00000000;
    rd_cycle[16528] = 1'b0;  wr_cycle[16528] = 1'b0;  addr_rom[16528]='h00000000;  wr_data_rom[16528]='h00000000;
    rd_cycle[16529] = 1'b0;  wr_cycle[16529] = 1'b0;  addr_rom[16529]='h00000000;  wr_data_rom[16529]='h00000000;
    rd_cycle[16530] = 1'b0;  wr_cycle[16530] = 1'b0;  addr_rom[16530]='h00000000;  wr_data_rom[16530]='h00000000;
    rd_cycle[16531] = 1'b0;  wr_cycle[16531] = 1'b0;  addr_rom[16531]='h00000000;  wr_data_rom[16531]='h00000000;
    rd_cycle[16532] = 1'b0;  wr_cycle[16532] = 1'b0;  addr_rom[16532]='h00000000;  wr_data_rom[16532]='h00000000;
    rd_cycle[16533] = 1'b0;  wr_cycle[16533] = 1'b0;  addr_rom[16533]='h00000000;  wr_data_rom[16533]='h00000000;
    rd_cycle[16534] = 1'b0;  wr_cycle[16534] = 1'b0;  addr_rom[16534]='h00000000;  wr_data_rom[16534]='h00000000;
    rd_cycle[16535] = 1'b0;  wr_cycle[16535] = 1'b0;  addr_rom[16535]='h00000000;  wr_data_rom[16535]='h00000000;
    rd_cycle[16536] = 1'b0;  wr_cycle[16536] = 1'b0;  addr_rom[16536]='h00000000;  wr_data_rom[16536]='h00000000;
    rd_cycle[16537] = 1'b0;  wr_cycle[16537] = 1'b0;  addr_rom[16537]='h00000000;  wr_data_rom[16537]='h00000000;
    rd_cycle[16538] = 1'b0;  wr_cycle[16538] = 1'b0;  addr_rom[16538]='h00000000;  wr_data_rom[16538]='h00000000;
    rd_cycle[16539] = 1'b0;  wr_cycle[16539] = 1'b0;  addr_rom[16539]='h00000000;  wr_data_rom[16539]='h00000000;
    rd_cycle[16540] = 1'b0;  wr_cycle[16540] = 1'b0;  addr_rom[16540]='h00000000;  wr_data_rom[16540]='h00000000;
    rd_cycle[16541] = 1'b0;  wr_cycle[16541] = 1'b0;  addr_rom[16541]='h00000000;  wr_data_rom[16541]='h00000000;
    rd_cycle[16542] = 1'b0;  wr_cycle[16542] = 1'b0;  addr_rom[16542]='h00000000;  wr_data_rom[16542]='h00000000;
    rd_cycle[16543] = 1'b0;  wr_cycle[16543] = 1'b0;  addr_rom[16543]='h00000000;  wr_data_rom[16543]='h00000000;
    rd_cycle[16544] = 1'b0;  wr_cycle[16544] = 1'b0;  addr_rom[16544]='h00000000;  wr_data_rom[16544]='h00000000;
    rd_cycle[16545] = 1'b0;  wr_cycle[16545] = 1'b0;  addr_rom[16545]='h00000000;  wr_data_rom[16545]='h00000000;
    rd_cycle[16546] = 1'b0;  wr_cycle[16546] = 1'b0;  addr_rom[16546]='h00000000;  wr_data_rom[16546]='h00000000;
    rd_cycle[16547] = 1'b0;  wr_cycle[16547] = 1'b0;  addr_rom[16547]='h00000000;  wr_data_rom[16547]='h00000000;
    rd_cycle[16548] = 1'b0;  wr_cycle[16548] = 1'b0;  addr_rom[16548]='h00000000;  wr_data_rom[16548]='h00000000;
    rd_cycle[16549] = 1'b0;  wr_cycle[16549] = 1'b0;  addr_rom[16549]='h00000000;  wr_data_rom[16549]='h00000000;
    rd_cycle[16550] = 1'b0;  wr_cycle[16550] = 1'b0;  addr_rom[16550]='h00000000;  wr_data_rom[16550]='h00000000;
    rd_cycle[16551] = 1'b0;  wr_cycle[16551] = 1'b0;  addr_rom[16551]='h00000000;  wr_data_rom[16551]='h00000000;
    rd_cycle[16552] = 1'b0;  wr_cycle[16552] = 1'b0;  addr_rom[16552]='h00000000;  wr_data_rom[16552]='h00000000;
    rd_cycle[16553] = 1'b0;  wr_cycle[16553] = 1'b0;  addr_rom[16553]='h00000000;  wr_data_rom[16553]='h00000000;
    rd_cycle[16554] = 1'b0;  wr_cycle[16554] = 1'b0;  addr_rom[16554]='h00000000;  wr_data_rom[16554]='h00000000;
    rd_cycle[16555] = 1'b0;  wr_cycle[16555] = 1'b0;  addr_rom[16555]='h00000000;  wr_data_rom[16555]='h00000000;
    rd_cycle[16556] = 1'b0;  wr_cycle[16556] = 1'b0;  addr_rom[16556]='h00000000;  wr_data_rom[16556]='h00000000;
    rd_cycle[16557] = 1'b0;  wr_cycle[16557] = 1'b0;  addr_rom[16557]='h00000000;  wr_data_rom[16557]='h00000000;
    rd_cycle[16558] = 1'b0;  wr_cycle[16558] = 1'b0;  addr_rom[16558]='h00000000;  wr_data_rom[16558]='h00000000;
    rd_cycle[16559] = 1'b0;  wr_cycle[16559] = 1'b0;  addr_rom[16559]='h00000000;  wr_data_rom[16559]='h00000000;
    rd_cycle[16560] = 1'b0;  wr_cycle[16560] = 1'b0;  addr_rom[16560]='h00000000;  wr_data_rom[16560]='h00000000;
    rd_cycle[16561] = 1'b0;  wr_cycle[16561] = 1'b0;  addr_rom[16561]='h00000000;  wr_data_rom[16561]='h00000000;
    rd_cycle[16562] = 1'b0;  wr_cycle[16562] = 1'b0;  addr_rom[16562]='h00000000;  wr_data_rom[16562]='h00000000;
    rd_cycle[16563] = 1'b0;  wr_cycle[16563] = 1'b0;  addr_rom[16563]='h00000000;  wr_data_rom[16563]='h00000000;
    rd_cycle[16564] = 1'b0;  wr_cycle[16564] = 1'b0;  addr_rom[16564]='h00000000;  wr_data_rom[16564]='h00000000;
    rd_cycle[16565] = 1'b0;  wr_cycle[16565] = 1'b0;  addr_rom[16565]='h00000000;  wr_data_rom[16565]='h00000000;
    rd_cycle[16566] = 1'b0;  wr_cycle[16566] = 1'b0;  addr_rom[16566]='h00000000;  wr_data_rom[16566]='h00000000;
    rd_cycle[16567] = 1'b0;  wr_cycle[16567] = 1'b0;  addr_rom[16567]='h00000000;  wr_data_rom[16567]='h00000000;
    rd_cycle[16568] = 1'b0;  wr_cycle[16568] = 1'b0;  addr_rom[16568]='h00000000;  wr_data_rom[16568]='h00000000;
    rd_cycle[16569] = 1'b0;  wr_cycle[16569] = 1'b0;  addr_rom[16569]='h00000000;  wr_data_rom[16569]='h00000000;
    rd_cycle[16570] = 1'b0;  wr_cycle[16570] = 1'b0;  addr_rom[16570]='h00000000;  wr_data_rom[16570]='h00000000;
    rd_cycle[16571] = 1'b0;  wr_cycle[16571] = 1'b0;  addr_rom[16571]='h00000000;  wr_data_rom[16571]='h00000000;
    rd_cycle[16572] = 1'b0;  wr_cycle[16572] = 1'b0;  addr_rom[16572]='h00000000;  wr_data_rom[16572]='h00000000;
    rd_cycle[16573] = 1'b0;  wr_cycle[16573] = 1'b0;  addr_rom[16573]='h00000000;  wr_data_rom[16573]='h00000000;
    rd_cycle[16574] = 1'b0;  wr_cycle[16574] = 1'b0;  addr_rom[16574]='h00000000;  wr_data_rom[16574]='h00000000;
    rd_cycle[16575] = 1'b0;  wr_cycle[16575] = 1'b0;  addr_rom[16575]='h00000000;  wr_data_rom[16575]='h00000000;
    rd_cycle[16576] = 1'b0;  wr_cycle[16576] = 1'b0;  addr_rom[16576]='h00000000;  wr_data_rom[16576]='h00000000;
    rd_cycle[16577] = 1'b0;  wr_cycle[16577] = 1'b0;  addr_rom[16577]='h00000000;  wr_data_rom[16577]='h00000000;
    rd_cycle[16578] = 1'b0;  wr_cycle[16578] = 1'b0;  addr_rom[16578]='h00000000;  wr_data_rom[16578]='h00000000;
    rd_cycle[16579] = 1'b0;  wr_cycle[16579] = 1'b0;  addr_rom[16579]='h00000000;  wr_data_rom[16579]='h00000000;
    rd_cycle[16580] = 1'b0;  wr_cycle[16580] = 1'b0;  addr_rom[16580]='h00000000;  wr_data_rom[16580]='h00000000;
    rd_cycle[16581] = 1'b0;  wr_cycle[16581] = 1'b0;  addr_rom[16581]='h00000000;  wr_data_rom[16581]='h00000000;
    rd_cycle[16582] = 1'b0;  wr_cycle[16582] = 1'b0;  addr_rom[16582]='h00000000;  wr_data_rom[16582]='h00000000;
    rd_cycle[16583] = 1'b0;  wr_cycle[16583] = 1'b0;  addr_rom[16583]='h00000000;  wr_data_rom[16583]='h00000000;
    rd_cycle[16584] = 1'b0;  wr_cycle[16584] = 1'b0;  addr_rom[16584]='h00000000;  wr_data_rom[16584]='h00000000;
    rd_cycle[16585] = 1'b0;  wr_cycle[16585] = 1'b0;  addr_rom[16585]='h00000000;  wr_data_rom[16585]='h00000000;
    rd_cycle[16586] = 1'b0;  wr_cycle[16586] = 1'b0;  addr_rom[16586]='h00000000;  wr_data_rom[16586]='h00000000;
    rd_cycle[16587] = 1'b0;  wr_cycle[16587] = 1'b0;  addr_rom[16587]='h00000000;  wr_data_rom[16587]='h00000000;
    rd_cycle[16588] = 1'b0;  wr_cycle[16588] = 1'b0;  addr_rom[16588]='h00000000;  wr_data_rom[16588]='h00000000;
    rd_cycle[16589] = 1'b0;  wr_cycle[16589] = 1'b0;  addr_rom[16589]='h00000000;  wr_data_rom[16589]='h00000000;
    rd_cycle[16590] = 1'b0;  wr_cycle[16590] = 1'b0;  addr_rom[16590]='h00000000;  wr_data_rom[16590]='h00000000;
    rd_cycle[16591] = 1'b0;  wr_cycle[16591] = 1'b0;  addr_rom[16591]='h00000000;  wr_data_rom[16591]='h00000000;
    rd_cycle[16592] = 1'b0;  wr_cycle[16592] = 1'b0;  addr_rom[16592]='h00000000;  wr_data_rom[16592]='h00000000;
    rd_cycle[16593] = 1'b0;  wr_cycle[16593] = 1'b0;  addr_rom[16593]='h00000000;  wr_data_rom[16593]='h00000000;
    rd_cycle[16594] = 1'b0;  wr_cycle[16594] = 1'b0;  addr_rom[16594]='h00000000;  wr_data_rom[16594]='h00000000;
    rd_cycle[16595] = 1'b0;  wr_cycle[16595] = 1'b0;  addr_rom[16595]='h00000000;  wr_data_rom[16595]='h00000000;
    rd_cycle[16596] = 1'b0;  wr_cycle[16596] = 1'b0;  addr_rom[16596]='h00000000;  wr_data_rom[16596]='h00000000;
    rd_cycle[16597] = 1'b0;  wr_cycle[16597] = 1'b0;  addr_rom[16597]='h00000000;  wr_data_rom[16597]='h00000000;
    rd_cycle[16598] = 1'b0;  wr_cycle[16598] = 1'b0;  addr_rom[16598]='h00000000;  wr_data_rom[16598]='h00000000;
    rd_cycle[16599] = 1'b0;  wr_cycle[16599] = 1'b0;  addr_rom[16599]='h00000000;  wr_data_rom[16599]='h00000000;
    rd_cycle[16600] = 1'b0;  wr_cycle[16600] = 1'b0;  addr_rom[16600]='h00000000;  wr_data_rom[16600]='h00000000;
    rd_cycle[16601] = 1'b0;  wr_cycle[16601] = 1'b0;  addr_rom[16601]='h00000000;  wr_data_rom[16601]='h00000000;
    rd_cycle[16602] = 1'b0;  wr_cycle[16602] = 1'b0;  addr_rom[16602]='h00000000;  wr_data_rom[16602]='h00000000;
    rd_cycle[16603] = 1'b0;  wr_cycle[16603] = 1'b0;  addr_rom[16603]='h00000000;  wr_data_rom[16603]='h00000000;
    rd_cycle[16604] = 1'b0;  wr_cycle[16604] = 1'b0;  addr_rom[16604]='h00000000;  wr_data_rom[16604]='h00000000;
    rd_cycle[16605] = 1'b0;  wr_cycle[16605] = 1'b0;  addr_rom[16605]='h00000000;  wr_data_rom[16605]='h00000000;
    rd_cycle[16606] = 1'b0;  wr_cycle[16606] = 1'b0;  addr_rom[16606]='h00000000;  wr_data_rom[16606]='h00000000;
    rd_cycle[16607] = 1'b0;  wr_cycle[16607] = 1'b0;  addr_rom[16607]='h00000000;  wr_data_rom[16607]='h00000000;
    rd_cycle[16608] = 1'b0;  wr_cycle[16608] = 1'b0;  addr_rom[16608]='h00000000;  wr_data_rom[16608]='h00000000;
    rd_cycle[16609] = 1'b0;  wr_cycle[16609] = 1'b0;  addr_rom[16609]='h00000000;  wr_data_rom[16609]='h00000000;
    rd_cycle[16610] = 1'b0;  wr_cycle[16610] = 1'b0;  addr_rom[16610]='h00000000;  wr_data_rom[16610]='h00000000;
    rd_cycle[16611] = 1'b0;  wr_cycle[16611] = 1'b0;  addr_rom[16611]='h00000000;  wr_data_rom[16611]='h00000000;
    rd_cycle[16612] = 1'b0;  wr_cycle[16612] = 1'b0;  addr_rom[16612]='h00000000;  wr_data_rom[16612]='h00000000;
    rd_cycle[16613] = 1'b0;  wr_cycle[16613] = 1'b0;  addr_rom[16613]='h00000000;  wr_data_rom[16613]='h00000000;
    rd_cycle[16614] = 1'b0;  wr_cycle[16614] = 1'b0;  addr_rom[16614]='h00000000;  wr_data_rom[16614]='h00000000;
    rd_cycle[16615] = 1'b0;  wr_cycle[16615] = 1'b0;  addr_rom[16615]='h00000000;  wr_data_rom[16615]='h00000000;
    rd_cycle[16616] = 1'b0;  wr_cycle[16616] = 1'b0;  addr_rom[16616]='h00000000;  wr_data_rom[16616]='h00000000;
    rd_cycle[16617] = 1'b0;  wr_cycle[16617] = 1'b0;  addr_rom[16617]='h00000000;  wr_data_rom[16617]='h00000000;
    rd_cycle[16618] = 1'b0;  wr_cycle[16618] = 1'b0;  addr_rom[16618]='h00000000;  wr_data_rom[16618]='h00000000;
    rd_cycle[16619] = 1'b0;  wr_cycle[16619] = 1'b0;  addr_rom[16619]='h00000000;  wr_data_rom[16619]='h00000000;
    rd_cycle[16620] = 1'b0;  wr_cycle[16620] = 1'b0;  addr_rom[16620]='h00000000;  wr_data_rom[16620]='h00000000;
    rd_cycle[16621] = 1'b0;  wr_cycle[16621] = 1'b0;  addr_rom[16621]='h00000000;  wr_data_rom[16621]='h00000000;
    rd_cycle[16622] = 1'b0;  wr_cycle[16622] = 1'b0;  addr_rom[16622]='h00000000;  wr_data_rom[16622]='h00000000;
    rd_cycle[16623] = 1'b0;  wr_cycle[16623] = 1'b0;  addr_rom[16623]='h00000000;  wr_data_rom[16623]='h00000000;
    rd_cycle[16624] = 1'b0;  wr_cycle[16624] = 1'b0;  addr_rom[16624]='h00000000;  wr_data_rom[16624]='h00000000;
    rd_cycle[16625] = 1'b0;  wr_cycle[16625] = 1'b0;  addr_rom[16625]='h00000000;  wr_data_rom[16625]='h00000000;
    rd_cycle[16626] = 1'b0;  wr_cycle[16626] = 1'b0;  addr_rom[16626]='h00000000;  wr_data_rom[16626]='h00000000;
    rd_cycle[16627] = 1'b0;  wr_cycle[16627] = 1'b0;  addr_rom[16627]='h00000000;  wr_data_rom[16627]='h00000000;
    rd_cycle[16628] = 1'b0;  wr_cycle[16628] = 1'b0;  addr_rom[16628]='h00000000;  wr_data_rom[16628]='h00000000;
    rd_cycle[16629] = 1'b0;  wr_cycle[16629] = 1'b0;  addr_rom[16629]='h00000000;  wr_data_rom[16629]='h00000000;
    rd_cycle[16630] = 1'b0;  wr_cycle[16630] = 1'b0;  addr_rom[16630]='h00000000;  wr_data_rom[16630]='h00000000;
    rd_cycle[16631] = 1'b0;  wr_cycle[16631] = 1'b0;  addr_rom[16631]='h00000000;  wr_data_rom[16631]='h00000000;
    rd_cycle[16632] = 1'b0;  wr_cycle[16632] = 1'b0;  addr_rom[16632]='h00000000;  wr_data_rom[16632]='h00000000;
    rd_cycle[16633] = 1'b0;  wr_cycle[16633] = 1'b0;  addr_rom[16633]='h00000000;  wr_data_rom[16633]='h00000000;
    rd_cycle[16634] = 1'b0;  wr_cycle[16634] = 1'b0;  addr_rom[16634]='h00000000;  wr_data_rom[16634]='h00000000;
    rd_cycle[16635] = 1'b0;  wr_cycle[16635] = 1'b0;  addr_rom[16635]='h00000000;  wr_data_rom[16635]='h00000000;
    rd_cycle[16636] = 1'b0;  wr_cycle[16636] = 1'b0;  addr_rom[16636]='h00000000;  wr_data_rom[16636]='h00000000;
    rd_cycle[16637] = 1'b0;  wr_cycle[16637] = 1'b0;  addr_rom[16637]='h00000000;  wr_data_rom[16637]='h00000000;
    rd_cycle[16638] = 1'b0;  wr_cycle[16638] = 1'b0;  addr_rom[16638]='h00000000;  wr_data_rom[16638]='h00000000;
    rd_cycle[16639] = 1'b0;  wr_cycle[16639] = 1'b0;  addr_rom[16639]='h00000000;  wr_data_rom[16639]='h00000000;
    rd_cycle[16640] = 1'b0;  wr_cycle[16640] = 1'b0;  addr_rom[16640]='h00000000;  wr_data_rom[16640]='h00000000;
    rd_cycle[16641] = 1'b0;  wr_cycle[16641] = 1'b0;  addr_rom[16641]='h00000000;  wr_data_rom[16641]='h00000000;
    rd_cycle[16642] = 1'b0;  wr_cycle[16642] = 1'b0;  addr_rom[16642]='h00000000;  wr_data_rom[16642]='h00000000;
    rd_cycle[16643] = 1'b0;  wr_cycle[16643] = 1'b0;  addr_rom[16643]='h00000000;  wr_data_rom[16643]='h00000000;
    rd_cycle[16644] = 1'b0;  wr_cycle[16644] = 1'b0;  addr_rom[16644]='h00000000;  wr_data_rom[16644]='h00000000;
    rd_cycle[16645] = 1'b0;  wr_cycle[16645] = 1'b0;  addr_rom[16645]='h00000000;  wr_data_rom[16645]='h00000000;
    rd_cycle[16646] = 1'b0;  wr_cycle[16646] = 1'b0;  addr_rom[16646]='h00000000;  wr_data_rom[16646]='h00000000;
    rd_cycle[16647] = 1'b0;  wr_cycle[16647] = 1'b0;  addr_rom[16647]='h00000000;  wr_data_rom[16647]='h00000000;
    rd_cycle[16648] = 1'b0;  wr_cycle[16648] = 1'b0;  addr_rom[16648]='h00000000;  wr_data_rom[16648]='h00000000;
    rd_cycle[16649] = 1'b0;  wr_cycle[16649] = 1'b0;  addr_rom[16649]='h00000000;  wr_data_rom[16649]='h00000000;
    rd_cycle[16650] = 1'b0;  wr_cycle[16650] = 1'b0;  addr_rom[16650]='h00000000;  wr_data_rom[16650]='h00000000;
    rd_cycle[16651] = 1'b0;  wr_cycle[16651] = 1'b0;  addr_rom[16651]='h00000000;  wr_data_rom[16651]='h00000000;
    rd_cycle[16652] = 1'b0;  wr_cycle[16652] = 1'b0;  addr_rom[16652]='h00000000;  wr_data_rom[16652]='h00000000;
    rd_cycle[16653] = 1'b0;  wr_cycle[16653] = 1'b0;  addr_rom[16653]='h00000000;  wr_data_rom[16653]='h00000000;
    rd_cycle[16654] = 1'b0;  wr_cycle[16654] = 1'b0;  addr_rom[16654]='h00000000;  wr_data_rom[16654]='h00000000;
    rd_cycle[16655] = 1'b0;  wr_cycle[16655] = 1'b0;  addr_rom[16655]='h00000000;  wr_data_rom[16655]='h00000000;
    rd_cycle[16656] = 1'b0;  wr_cycle[16656] = 1'b0;  addr_rom[16656]='h00000000;  wr_data_rom[16656]='h00000000;
    rd_cycle[16657] = 1'b0;  wr_cycle[16657] = 1'b0;  addr_rom[16657]='h00000000;  wr_data_rom[16657]='h00000000;
    rd_cycle[16658] = 1'b0;  wr_cycle[16658] = 1'b0;  addr_rom[16658]='h00000000;  wr_data_rom[16658]='h00000000;
    rd_cycle[16659] = 1'b0;  wr_cycle[16659] = 1'b0;  addr_rom[16659]='h00000000;  wr_data_rom[16659]='h00000000;
    rd_cycle[16660] = 1'b0;  wr_cycle[16660] = 1'b0;  addr_rom[16660]='h00000000;  wr_data_rom[16660]='h00000000;
    rd_cycle[16661] = 1'b0;  wr_cycle[16661] = 1'b0;  addr_rom[16661]='h00000000;  wr_data_rom[16661]='h00000000;
    rd_cycle[16662] = 1'b0;  wr_cycle[16662] = 1'b0;  addr_rom[16662]='h00000000;  wr_data_rom[16662]='h00000000;
    rd_cycle[16663] = 1'b0;  wr_cycle[16663] = 1'b0;  addr_rom[16663]='h00000000;  wr_data_rom[16663]='h00000000;
    rd_cycle[16664] = 1'b0;  wr_cycle[16664] = 1'b0;  addr_rom[16664]='h00000000;  wr_data_rom[16664]='h00000000;
    rd_cycle[16665] = 1'b0;  wr_cycle[16665] = 1'b0;  addr_rom[16665]='h00000000;  wr_data_rom[16665]='h00000000;
    rd_cycle[16666] = 1'b0;  wr_cycle[16666] = 1'b0;  addr_rom[16666]='h00000000;  wr_data_rom[16666]='h00000000;
    rd_cycle[16667] = 1'b0;  wr_cycle[16667] = 1'b0;  addr_rom[16667]='h00000000;  wr_data_rom[16667]='h00000000;
    rd_cycle[16668] = 1'b0;  wr_cycle[16668] = 1'b0;  addr_rom[16668]='h00000000;  wr_data_rom[16668]='h00000000;
    rd_cycle[16669] = 1'b0;  wr_cycle[16669] = 1'b0;  addr_rom[16669]='h00000000;  wr_data_rom[16669]='h00000000;
    rd_cycle[16670] = 1'b0;  wr_cycle[16670] = 1'b0;  addr_rom[16670]='h00000000;  wr_data_rom[16670]='h00000000;
    rd_cycle[16671] = 1'b0;  wr_cycle[16671] = 1'b0;  addr_rom[16671]='h00000000;  wr_data_rom[16671]='h00000000;
    rd_cycle[16672] = 1'b0;  wr_cycle[16672] = 1'b0;  addr_rom[16672]='h00000000;  wr_data_rom[16672]='h00000000;
    rd_cycle[16673] = 1'b0;  wr_cycle[16673] = 1'b0;  addr_rom[16673]='h00000000;  wr_data_rom[16673]='h00000000;
    rd_cycle[16674] = 1'b0;  wr_cycle[16674] = 1'b0;  addr_rom[16674]='h00000000;  wr_data_rom[16674]='h00000000;
    rd_cycle[16675] = 1'b0;  wr_cycle[16675] = 1'b0;  addr_rom[16675]='h00000000;  wr_data_rom[16675]='h00000000;
    rd_cycle[16676] = 1'b0;  wr_cycle[16676] = 1'b0;  addr_rom[16676]='h00000000;  wr_data_rom[16676]='h00000000;
    rd_cycle[16677] = 1'b0;  wr_cycle[16677] = 1'b0;  addr_rom[16677]='h00000000;  wr_data_rom[16677]='h00000000;
    rd_cycle[16678] = 1'b0;  wr_cycle[16678] = 1'b0;  addr_rom[16678]='h00000000;  wr_data_rom[16678]='h00000000;
    rd_cycle[16679] = 1'b0;  wr_cycle[16679] = 1'b0;  addr_rom[16679]='h00000000;  wr_data_rom[16679]='h00000000;
    rd_cycle[16680] = 1'b0;  wr_cycle[16680] = 1'b0;  addr_rom[16680]='h00000000;  wr_data_rom[16680]='h00000000;
    rd_cycle[16681] = 1'b0;  wr_cycle[16681] = 1'b0;  addr_rom[16681]='h00000000;  wr_data_rom[16681]='h00000000;
    rd_cycle[16682] = 1'b0;  wr_cycle[16682] = 1'b0;  addr_rom[16682]='h00000000;  wr_data_rom[16682]='h00000000;
    rd_cycle[16683] = 1'b0;  wr_cycle[16683] = 1'b0;  addr_rom[16683]='h00000000;  wr_data_rom[16683]='h00000000;
    rd_cycle[16684] = 1'b0;  wr_cycle[16684] = 1'b0;  addr_rom[16684]='h00000000;  wr_data_rom[16684]='h00000000;
    rd_cycle[16685] = 1'b0;  wr_cycle[16685] = 1'b0;  addr_rom[16685]='h00000000;  wr_data_rom[16685]='h00000000;
    rd_cycle[16686] = 1'b0;  wr_cycle[16686] = 1'b0;  addr_rom[16686]='h00000000;  wr_data_rom[16686]='h00000000;
    rd_cycle[16687] = 1'b0;  wr_cycle[16687] = 1'b0;  addr_rom[16687]='h00000000;  wr_data_rom[16687]='h00000000;
    rd_cycle[16688] = 1'b0;  wr_cycle[16688] = 1'b0;  addr_rom[16688]='h00000000;  wr_data_rom[16688]='h00000000;
    rd_cycle[16689] = 1'b0;  wr_cycle[16689] = 1'b0;  addr_rom[16689]='h00000000;  wr_data_rom[16689]='h00000000;
    rd_cycle[16690] = 1'b0;  wr_cycle[16690] = 1'b0;  addr_rom[16690]='h00000000;  wr_data_rom[16690]='h00000000;
    rd_cycle[16691] = 1'b0;  wr_cycle[16691] = 1'b0;  addr_rom[16691]='h00000000;  wr_data_rom[16691]='h00000000;
    rd_cycle[16692] = 1'b0;  wr_cycle[16692] = 1'b0;  addr_rom[16692]='h00000000;  wr_data_rom[16692]='h00000000;
    rd_cycle[16693] = 1'b0;  wr_cycle[16693] = 1'b0;  addr_rom[16693]='h00000000;  wr_data_rom[16693]='h00000000;
    rd_cycle[16694] = 1'b0;  wr_cycle[16694] = 1'b0;  addr_rom[16694]='h00000000;  wr_data_rom[16694]='h00000000;
    rd_cycle[16695] = 1'b0;  wr_cycle[16695] = 1'b0;  addr_rom[16695]='h00000000;  wr_data_rom[16695]='h00000000;
    rd_cycle[16696] = 1'b0;  wr_cycle[16696] = 1'b0;  addr_rom[16696]='h00000000;  wr_data_rom[16696]='h00000000;
    rd_cycle[16697] = 1'b0;  wr_cycle[16697] = 1'b0;  addr_rom[16697]='h00000000;  wr_data_rom[16697]='h00000000;
    rd_cycle[16698] = 1'b0;  wr_cycle[16698] = 1'b0;  addr_rom[16698]='h00000000;  wr_data_rom[16698]='h00000000;
    rd_cycle[16699] = 1'b0;  wr_cycle[16699] = 1'b0;  addr_rom[16699]='h00000000;  wr_data_rom[16699]='h00000000;
    rd_cycle[16700] = 1'b0;  wr_cycle[16700] = 1'b0;  addr_rom[16700]='h00000000;  wr_data_rom[16700]='h00000000;
    rd_cycle[16701] = 1'b0;  wr_cycle[16701] = 1'b0;  addr_rom[16701]='h00000000;  wr_data_rom[16701]='h00000000;
    rd_cycle[16702] = 1'b0;  wr_cycle[16702] = 1'b0;  addr_rom[16702]='h00000000;  wr_data_rom[16702]='h00000000;
    rd_cycle[16703] = 1'b0;  wr_cycle[16703] = 1'b0;  addr_rom[16703]='h00000000;  wr_data_rom[16703]='h00000000;
    rd_cycle[16704] = 1'b0;  wr_cycle[16704] = 1'b0;  addr_rom[16704]='h00000000;  wr_data_rom[16704]='h00000000;
    rd_cycle[16705] = 1'b0;  wr_cycle[16705] = 1'b0;  addr_rom[16705]='h00000000;  wr_data_rom[16705]='h00000000;
    rd_cycle[16706] = 1'b0;  wr_cycle[16706] = 1'b0;  addr_rom[16706]='h00000000;  wr_data_rom[16706]='h00000000;
    rd_cycle[16707] = 1'b0;  wr_cycle[16707] = 1'b0;  addr_rom[16707]='h00000000;  wr_data_rom[16707]='h00000000;
    rd_cycle[16708] = 1'b0;  wr_cycle[16708] = 1'b0;  addr_rom[16708]='h00000000;  wr_data_rom[16708]='h00000000;
    rd_cycle[16709] = 1'b0;  wr_cycle[16709] = 1'b0;  addr_rom[16709]='h00000000;  wr_data_rom[16709]='h00000000;
    rd_cycle[16710] = 1'b0;  wr_cycle[16710] = 1'b0;  addr_rom[16710]='h00000000;  wr_data_rom[16710]='h00000000;
    rd_cycle[16711] = 1'b0;  wr_cycle[16711] = 1'b0;  addr_rom[16711]='h00000000;  wr_data_rom[16711]='h00000000;
    rd_cycle[16712] = 1'b0;  wr_cycle[16712] = 1'b0;  addr_rom[16712]='h00000000;  wr_data_rom[16712]='h00000000;
    rd_cycle[16713] = 1'b0;  wr_cycle[16713] = 1'b0;  addr_rom[16713]='h00000000;  wr_data_rom[16713]='h00000000;
    rd_cycle[16714] = 1'b0;  wr_cycle[16714] = 1'b0;  addr_rom[16714]='h00000000;  wr_data_rom[16714]='h00000000;
    rd_cycle[16715] = 1'b0;  wr_cycle[16715] = 1'b0;  addr_rom[16715]='h00000000;  wr_data_rom[16715]='h00000000;
    rd_cycle[16716] = 1'b0;  wr_cycle[16716] = 1'b0;  addr_rom[16716]='h00000000;  wr_data_rom[16716]='h00000000;
    rd_cycle[16717] = 1'b0;  wr_cycle[16717] = 1'b0;  addr_rom[16717]='h00000000;  wr_data_rom[16717]='h00000000;
    rd_cycle[16718] = 1'b0;  wr_cycle[16718] = 1'b0;  addr_rom[16718]='h00000000;  wr_data_rom[16718]='h00000000;
    rd_cycle[16719] = 1'b0;  wr_cycle[16719] = 1'b0;  addr_rom[16719]='h00000000;  wr_data_rom[16719]='h00000000;
    rd_cycle[16720] = 1'b0;  wr_cycle[16720] = 1'b0;  addr_rom[16720]='h00000000;  wr_data_rom[16720]='h00000000;
    rd_cycle[16721] = 1'b0;  wr_cycle[16721] = 1'b0;  addr_rom[16721]='h00000000;  wr_data_rom[16721]='h00000000;
    rd_cycle[16722] = 1'b0;  wr_cycle[16722] = 1'b0;  addr_rom[16722]='h00000000;  wr_data_rom[16722]='h00000000;
    rd_cycle[16723] = 1'b0;  wr_cycle[16723] = 1'b0;  addr_rom[16723]='h00000000;  wr_data_rom[16723]='h00000000;
    rd_cycle[16724] = 1'b0;  wr_cycle[16724] = 1'b0;  addr_rom[16724]='h00000000;  wr_data_rom[16724]='h00000000;
    rd_cycle[16725] = 1'b0;  wr_cycle[16725] = 1'b0;  addr_rom[16725]='h00000000;  wr_data_rom[16725]='h00000000;
    rd_cycle[16726] = 1'b0;  wr_cycle[16726] = 1'b0;  addr_rom[16726]='h00000000;  wr_data_rom[16726]='h00000000;
    rd_cycle[16727] = 1'b0;  wr_cycle[16727] = 1'b0;  addr_rom[16727]='h00000000;  wr_data_rom[16727]='h00000000;
    rd_cycle[16728] = 1'b0;  wr_cycle[16728] = 1'b0;  addr_rom[16728]='h00000000;  wr_data_rom[16728]='h00000000;
    rd_cycle[16729] = 1'b0;  wr_cycle[16729] = 1'b0;  addr_rom[16729]='h00000000;  wr_data_rom[16729]='h00000000;
    rd_cycle[16730] = 1'b0;  wr_cycle[16730] = 1'b0;  addr_rom[16730]='h00000000;  wr_data_rom[16730]='h00000000;
    rd_cycle[16731] = 1'b0;  wr_cycle[16731] = 1'b0;  addr_rom[16731]='h00000000;  wr_data_rom[16731]='h00000000;
    rd_cycle[16732] = 1'b0;  wr_cycle[16732] = 1'b0;  addr_rom[16732]='h00000000;  wr_data_rom[16732]='h00000000;
    rd_cycle[16733] = 1'b0;  wr_cycle[16733] = 1'b0;  addr_rom[16733]='h00000000;  wr_data_rom[16733]='h00000000;
    rd_cycle[16734] = 1'b0;  wr_cycle[16734] = 1'b0;  addr_rom[16734]='h00000000;  wr_data_rom[16734]='h00000000;
    rd_cycle[16735] = 1'b0;  wr_cycle[16735] = 1'b0;  addr_rom[16735]='h00000000;  wr_data_rom[16735]='h00000000;
    rd_cycle[16736] = 1'b0;  wr_cycle[16736] = 1'b0;  addr_rom[16736]='h00000000;  wr_data_rom[16736]='h00000000;
    rd_cycle[16737] = 1'b0;  wr_cycle[16737] = 1'b0;  addr_rom[16737]='h00000000;  wr_data_rom[16737]='h00000000;
    rd_cycle[16738] = 1'b0;  wr_cycle[16738] = 1'b0;  addr_rom[16738]='h00000000;  wr_data_rom[16738]='h00000000;
    rd_cycle[16739] = 1'b0;  wr_cycle[16739] = 1'b0;  addr_rom[16739]='h00000000;  wr_data_rom[16739]='h00000000;
    rd_cycle[16740] = 1'b0;  wr_cycle[16740] = 1'b0;  addr_rom[16740]='h00000000;  wr_data_rom[16740]='h00000000;
    rd_cycle[16741] = 1'b0;  wr_cycle[16741] = 1'b0;  addr_rom[16741]='h00000000;  wr_data_rom[16741]='h00000000;
    rd_cycle[16742] = 1'b0;  wr_cycle[16742] = 1'b0;  addr_rom[16742]='h00000000;  wr_data_rom[16742]='h00000000;
    rd_cycle[16743] = 1'b0;  wr_cycle[16743] = 1'b0;  addr_rom[16743]='h00000000;  wr_data_rom[16743]='h00000000;
    rd_cycle[16744] = 1'b0;  wr_cycle[16744] = 1'b0;  addr_rom[16744]='h00000000;  wr_data_rom[16744]='h00000000;
    rd_cycle[16745] = 1'b0;  wr_cycle[16745] = 1'b0;  addr_rom[16745]='h00000000;  wr_data_rom[16745]='h00000000;
    rd_cycle[16746] = 1'b0;  wr_cycle[16746] = 1'b0;  addr_rom[16746]='h00000000;  wr_data_rom[16746]='h00000000;
    rd_cycle[16747] = 1'b0;  wr_cycle[16747] = 1'b0;  addr_rom[16747]='h00000000;  wr_data_rom[16747]='h00000000;
    rd_cycle[16748] = 1'b0;  wr_cycle[16748] = 1'b0;  addr_rom[16748]='h00000000;  wr_data_rom[16748]='h00000000;
    rd_cycle[16749] = 1'b0;  wr_cycle[16749] = 1'b0;  addr_rom[16749]='h00000000;  wr_data_rom[16749]='h00000000;
    rd_cycle[16750] = 1'b0;  wr_cycle[16750] = 1'b0;  addr_rom[16750]='h00000000;  wr_data_rom[16750]='h00000000;
    rd_cycle[16751] = 1'b0;  wr_cycle[16751] = 1'b0;  addr_rom[16751]='h00000000;  wr_data_rom[16751]='h00000000;
    rd_cycle[16752] = 1'b0;  wr_cycle[16752] = 1'b0;  addr_rom[16752]='h00000000;  wr_data_rom[16752]='h00000000;
    rd_cycle[16753] = 1'b0;  wr_cycle[16753] = 1'b0;  addr_rom[16753]='h00000000;  wr_data_rom[16753]='h00000000;
    rd_cycle[16754] = 1'b0;  wr_cycle[16754] = 1'b0;  addr_rom[16754]='h00000000;  wr_data_rom[16754]='h00000000;
    rd_cycle[16755] = 1'b0;  wr_cycle[16755] = 1'b0;  addr_rom[16755]='h00000000;  wr_data_rom[16755]='h00000000;
    rd_cycle[16756] = 1'b0;  wr_cycle[16756] = 1'b0;  addr_rom[16756]='h00000000;  wr_data_rom[16756]='h00000000;
    rd_cycle[16757] = 1'b0;  wr_cycle[16757] = 1'b0;  addr_rom[16757]='h00000000;  wr_data_rom[16757]='h00000000;
    rd_cycle[16758] = 1'b0;  wr_cycle[16758] = 1'b0;  addr_rom[16758]='h00000000;  wr_data_rom[16758]='h00000000;
    rd_cycle[16759] = 1'b0;  wr_cycle[16759] = 1'b0;  addr_rom[16759]='h00000000;  wr_data_rom[16759]='h00000000;
    rd_cycle[16760] = 1'b0;  wr_cycle[16760] = 1'b0;  addr_rom[16760]='h00000000;  wr_data_rom[16760]='h00000000;
    rd_cycle[16761] = 1'b0;  wr_cycle[16761] = 1'b0;  addr_rom[16761]='h00000000;  wr_data_rom[16761]='h00000000;
    rd_cycle[16762] = 1'b0;  wr_cycle[16762] = 1'b0;  addr_rom[16762]='h00000000;  wr_data_rom[16762]='h00000000;
    rd_cycle[16763] = 1'b0;  wr_cycle[16763] = 1'b0;  addr_rom[16763]='h00000000;  wr_data_rom[16763]='h00000000;
    rd_cycle[16764] = 1'b0;  wr_cycle[16764] = 1'b0;  addr_rom[16764]='h00000000;  wr_data_rom[16764]='h00000000;
    rd_cycle[16765] = 1'b0;  wr_cycle[16765] = 1'b0;  addr_rom[16765]='h00000000;  wr_data_rom[16765]='h00000000;
    rd_cycle[16766] = 1'b0;  wr_cycle[16766] = 1'b0;  addr_rom[16766]='h00000000;  wr_data_rom[16766]='h00000000;
    rd_cycle[16767] = 1'b0;  wr_cycle[16767] = 1'b0;  addr_rom[16767]='h00000000;  wr_data_rom[16767]='h00000000;
    rd_cycle[16768] = 1'b0;  wr_cycle[16768] = 1'b0;  addr_rom[16768]='h00000000;  wr_data_rom[16768]='h00000000;
    rd_cycle[16769] = 1'b0;  wr_cycle[16769] = 1'b0;  addr_rom[16769]='h00000000;  wr_data_rom[16769]='h00000000;
    rd_cycle[16770] = 1'b0;  wr_cycle[16770] = 1'b0;  addr_rom[16770]='h00000000;  wr_data_rom[16770]='h00000000;
    rd_cycle[16771] = 1'b0;  wr_cycle[16771] = 1'b0;  addr_rom[16771]='h00000000;  wr_data_rom[16771]='h00000000;
    rd_cycle[16772] = 1'b0;  wr_cycle[16772] = 1'b0;  addr_rom[16772]='h00000000;  wr_data_rom[16772]='h00000000;
    rd_cycle[16773] = 1'b0;  wr_cycle[16773] = 1'b0;  addr_rom[16773]='h00000000;  wr_data_rom[16773]='h00000000;
    rd_cycle[16774] = 1'b0;  wr_cycle[16774] = 1'b0;  addr_rom[16774]='h00000000;  wr_data_rom[16774]='h00000000;
    rd_cycle[16775] = 1'b0;  wr_cycle[16775] = 1'b0;  addr_rom[16775]='h00000000;  wr_data_rom[16775]='h00000000;
    rd_cycle[16776] = 1'b0;  wr_cycle[16776] = 1'b0;  addr_rom[16776]='h00000000;  wr_data_rom[16776]='h00000000;
    rd_cycle[16777] = 1'b0;  wr_cycle[16777] = 1'b0;  addr_rom[16777]='h00000000;  wr_data_rom[16777]='h00000000;
    rd_cycle[16778] = 1'b0;  wr_cycle[16778] = 1'b0;  addr_rom[16778]='h00000000;  wr_data_rom[16778]='h00000000;
    rd_cycle[16779] = 1'b0;  wr_cycle[16779] = 1'b0;  addr_rom[16779]='h00000000;  wr_data_rom[16779]='h00000000;
    rd_cycle[16780] = 1'b0;  wr_cycle[16780] = 1'b0;  addr_rom[16780]='h00000000;  wr_data_rom[16780]='h00000000;
    rd_cycle[16781] = 1'b0;  wr_cycle[16781] = 1'b0;  addr_rom[16781]='h00000000;  wr_data_rom[16781]='h00000000;
    rd_cycle[16782] = 1'b0;  wr_cycle[16782] = 1'b0;  addr_rom[16782]='h00000000;  wr_data_rom[16782]='h00000000;
    rd_cycle[16783] = 1'b0;  wr_cycle[16783] = 1'b0;  addr_rom[16783]='h00000000;  wr_data_rom[16783]='h00000000;
    rd_cycle[16784] = 1'b0;  wr_cycle[16784] = 1'b0;  addr_rom[16784]='h00000000;  wr_data_rom[16784]='h00000000;
    rd_cycle[16785] = 1'b0;  wr_cycle[16785] = 1'b0;  addr_rom[16785]='h00000000;  wr_data_rom[16785]='h00000000;
    rd_cycle[16786] = 1'b0;  wr_cycle[16786] = 1'b0;  addr_rom[16786]='h00000000;  wr_data_rom[16786]='h00000000;
    rd_cycle[16787] = 1'b0;  wr_cycle[16787] = 1'b0;  addr_rom[16787]='h00000000;  wr_data_rom[16787]='h00000000;
    rd_cycle[16788] = 1'b0;  wr_cycle[16788] = 1'b0;  addr_rom[16788]='h00000000;  wr_data_rom[16788]='h00000000;
    rd_cycle[16789] = 1'b0;  wr_cycle[16789] = 1'b0;  addr_rom[16789]='h00000000;  wr_data_rom[16789]='h00000000;
    rd_cycle[16790] = 1'b0;  wr_cycle[16790] = 1'b0;  addr_rom[16790]='h00000000;  wr_data_rom[16790]='h00000000;
    rd_cycle[16791] = 1'b0;  wr_cycle[16791] = 1'b0;  addr_rom[16791]='h00000000;  wr_data_rom[16791]='h00000000;
    rd_cycle[16792] = 1'b0;  wr_cycle[16792] = 1'b0;  addr_rom[16792]='h00000000;  wr_data_rom[16792]='h00000000;
    rd_cycle[16793] = 1'b0;  wr_cycle[16793] = 1'b0;  addr_rom[16793]='h00000000;  wr_data_rom[16793]='h00000000;
    rd_cycle[16794] = 1'b0;  wr_cycle[16794] = 1'b0;  addr_rom[16794]='h00000000;  wr_data_rom[16794]='h00000000;
    rd_cycle[16795] = 1'b0;  wr_cycle[16795] = 1'b0;  addr_rom[16795]='h00000000;  wr_data_rom[16795]='h00000000;
    rd_cycle[16796] = 1'b0;  wr_cycle[16796] = 1'b0;  addr_rom[16796]='h00000000;  wr_data_rom[16796]='h00000000;
    rd_cycle[16797] = 1'b0;  wr_cycle[16797] = 1'b0;  addr_rom[16797]='h00000000;  wr_data_rom[16797]='h00000000;
    rd_cycle[16798] = 1'b0;  wr_cycle[16798] = 1'b0;  addr_rom[16798]='h00000000;  wr_data_rom[16798]='h00000000;
    rd_cycle[16799] = 1'b0;  wr_cycle[16799] = 1'b0;  addr_rom[16799]='h00000000;  wr_data_rom[16799]='h00000000;
    rd_cycle[16800] = 1'b0;  wr_cycle[16800] = 1'b0;  addr_rom[16800]='h00000000;  wr_data_rom[16800]='h00000000;
    rd_cycle[16801] = 1'b0;  wr_cycle[16801] = 1'b0;  addr_rom[16801]='h00000000;  wr_data_rom[16801]='h00000000;
    rd_cycle[16802] = 1'b0;  wr_cycle[16802] = 1'b0;  addr_rom[16802]='h00000000;  wr_data_rom[16802]='h00000000;
    rd_cycle[16803] = 1'b0;  wr_cycle[16803] = 1'b0;  addr_rom[16803]='h00000000;  wr_data_rom[16803]='h00000000;
    rd_cycle[16804] = 1'b0;  wr_cycle[16804] = 1'b0;  addr_rom[16804]='h00000000;  wr_data_rom[16804]='h00000000;
    rd_cycle[16805] = 1'b0;  wr_cycle[16805] = 1'b0;  addr_rom[16805]='h00000000;  wr_data_rom[16805]='h00000000;
    rd_cycle[16806] = 1'b0;  wr_cycle[16806] = 1'b0;  addr_rom[16806]='h00000000;  wr_data_rom[16806]='h00000000;
    rd_cycle[16807] = 1'b0;  wr_cycle[16807] = 1'b0;  addr_rom[16807]='h00000000;  wr_data_rom[16807]='h00000000;
    rd_cycle[16808] = 1'b0;  wr_cycle[16808] = 1'b0;  addr_rom[16808]='h00000000;  wr_data_rom[16808]='h00000000;
    rd_cycle[16809] = 1'b0;  wr_cycle[16809] = 1'b0;  addr_rom[16809]='h00000000;  wr_data_rom[16809]='h00000000;
    rd_cycle[16810] = 1'b0;  wr_cycle[16810] = 1'b0;  addr_rom[16810]='h00000000;  wr_data_rom[16810]='h00000000;
    rd_cycle[16811] = 1'b0;  wr_cycle[16811] = 1'b0;  addr_rom[16811]='h00000000;  wr_data_rom[16811]='h00000000;
    rd_cycle[16812] = 1'b0;  wr_cycle[16812] = 1'b0;  addr_rom[16812]='h00000000;  wr_data_rom[16812]='h00000000;
    rd_cycle[16813] = 1'b0;  wr_cycle[16813] = 1'b0;  addr_rom[16813]='h00000000;  wr_data_rom[16813]='h00000000;
    rd_cycle[16814] = 1'b0;  wr_cycle[16814] = 1'b0;  addr_rom[16814]='h00000000;  wr_data_rom[16814]='h00000000;
    rd_cycle[16815] = 1'b0;  wr_cycle[16815] = 1'b0;  addr_rom[16815]='h00000000;  wr_data_rom[16815]='h00000000;
    rd_cycle[16816] = 1'b0;  wr_cycle[16816] = 1'b0;  addr_rom[16816]='h00000000;  wr_data_rom[16816]='h00000000;
    rd_cycle[16817] = 1'b0;  wr_cycle[16817] = 1'b0;  addr_rom[16817]='h00000000;  wr_data_rom[16817]='h00000000;
    rd_cycle[16818] = 1'b0;  wr_cycle[16818] = 1'b0;  addr_rom[16818]='h00000000;  wr_data_rom[16818]='h00000000;
    rd_cycle[16819] = 1'b0;  wr_cycle[16819] = 1'b0;  addr_rom[16819]='h00000000;  wr_data_rom[16819]='h00000000;
    rd_cycle[16820] = 1'b0;  wr_cycle[16820] = 1'b0;  addr_rom[16820]='h00000000;  wr_data_rom[16820]='h00000000;
    rd_cycle[16821] = 1'b0;  wr_cycle[16821] = 1'b0;  addr_rom[16821]='h00000000;  wr_data_rom[16821]='h00000000;
    rd_cycle[16822] = 1'b0;  wr_cycle[16822] = 1'b0;  addr_rom[16822]='h00000000;  wr_data_rom[16822]='h00000000;
    rd_cycle[16823] = 1'b0;  wr_cycle[16823] = 1'b0;  addr_rom[16823]='h00000000;  wr_data_rom[16823]='h00000000;
    rd_cycle[16824] = 1'b0;  wr_cycle[16824] = 1'b0;  addr_rom[16824]='h00000000;  wr_data_rom[16824]='h00000000;
    rd_cycle[16825] = 1'b0;  wr_cycle[16825] = 1'b0;  addr_rom[16825]='h00000000;  wr_data_rom[16825]='h00000000;
    rd_cycle[16826] = 1'b0;  wr_cycle[16826] = 1'b0;  addr_rom[16826]='h00000000;  wr_data_rom[16826]='h00000000;
    rd_cycle[16827] = 1'b0;  wr_cycle[16827] = 1'b0;  addr_rom[16827]='h00000000;  wr_data_rom[16827]='h00000000;
    rd_cycle[16828] = 1'b0;  wr_cycle[16828] = 1'b0;  addr_rom[16828]='h00000000;  wr_data_rom[16828]='h00000000;
    rd_cycle[16829] = 1'b0;  wr_cycle[16829] = 1'b0;  addr_rom[16829]='h00000000;  wr_data_rom[16829]='h00000000;
    rd_cycle[16830] = 1'b0;  wr_cycle[16830] = 1'b0;  addr_rom[16830]='h00000000;  wr_data_rom[16830]='h00000000;
    rd_cycle[16831] = 1'b0;  wr_cycle[16831] = 1'b0;  addr_rom[16831]='h00000000;  wr_data_rom[16831]='h00000000;
    rd_cycle[16832] = 1'b0;  wr_cycle[16832] = 1'b0;  addr_rom[16832]='h00000000;  wr_data_rom[16832]='h00000000;
    rd_cycle[16833] = 1'b0;  wr_cycle[16833] = 1'b0;  addr_rom[16833]='h00000000;  wr_data_rom[16833]='h00000000;
    rd_cycle[16834] = 1'b0;  wr_cycle[16834] = 1'b0;  addr_rom[16834]='h00000000;  wr_data_rom[16834]='h00000000;
    rd_cycle[16835] = 1'b0;  wr_cycle[16835] = 1'b0;  addr_rom[16835]='h00000000;  wr_data_rom[16835]='h00000000;
    rd_cycle[16836] = 1'b0;  wr_cycle[16836] = 1'b0;  addr_rom[16836]='h00000000;  wr_data_rom[16836]='h00000000;
    rd_cycle[16837] = 1'b0;  wr_cycle[16837] = 1'b0;  addr_rom[16837]='h00000000;  wr_data_rom[16837]='h00000000;
    rd_cycle[16838] = 1'b0;  wr_cycle[16838] = 1'b0;  addr_rom[16838]='h00000000;  wr_data_rom[16838]='h00000000;
    rd_cycle[16839] = 1'b0;  wr_cycle[16839] = 1'b0;  addr_rom[16839]='h00000000;  wr_data_rom[16839]='h00000000;
    rd_cycle[16840] = 1'b0;  wr_cycle[16840] = 1'b0;  addr_rom[16840]='h00000000;  wr_data_rom[16840]='h00000000;
    rd_cycle[16841] = 1'b0;  wr_cycle[16841] = 1'b0;  addr_rom[16841]='h00000000;  wr_data_rom[16841]='h00000000;
    rd_cycle[16842] = 1'b0;  wr_cycle[16842] = 1'b0;  addr_rom[16842]='h00000000;  wr_data_rom[16842]='h00000000;
    rd_cycle[16843] = 1'b0;  wr_cycle[16843] = 1'b0;  addr_rom[16843]='h00000000;  wr_data_rom[16843]='h00000000;
    rd_cycle[16844] = 1'b0;  wr_cycle[16844] = 1'b0;  addr_rom[16844]='h00000000;  wr_data_rom[16844]='h00000000;
    rd_cycle[16845] = 1'b0;  wr_cycle[16845] = 1'b0;  addr_rom[16845]='h00000000;  wr_data_rom[16845]='h00000000;
    rd_cycle[16846] = 1'b0;  wr_cycle[16846] = 1'b0;  addr_rom[16846]='h00000000;  wr_data_rom[16846]='h00000000;
    rd_cycle[16847] = 1'b0;  wr_cycle[16847] = 1'b0;  addr_rom[16847]='h00000000;  wr_data_rom[16847]='h00000000;
    rd_cycle[16848] = 1'b0;  wr_cycle[16848] = 1'b0;  addr_rom[16848]='h00000000;  wr_data_rom[16848]='h00000000;
    rd_cycle[16849] = 1'b0;  wr_cycle[16849] = 1'b0;  addr_rom[16849]='h00000000;  wr_data_rom[16849]='h00000000;
    rd_cycle[16850] = 1'b0;  wr_cycle[16850] = 1'b0;  addr_rom[16850]='h00000000;  wr_data_rom[16850]='h00000000;
    rd_cycle[16851] = 1'b0;  wr_cycle[16851] = 1'b0;  addr_rom[16851]='h00000000;  wr_data_rom[16851]='h00000000;
    rd_cycle[16852] = 1'b0;  wr_cycle[16852] = 1'b0;  addr_rom[16852]='h00000000;  wr_data_rom[16852]='h00000000;
    rd_cycle[16853] = 1'b0;  wr_cycle[16853] = 1'b0;  addr_rom[16853]='h00000000;  wr_data_rom[16853]='h00000000;
    rd_cycle[16854] = 1'b0;  wr_cycle[16854] = 1'b0;  addr_rom[16854]='h00000000;  wr_data_rom[16854]='h00000000;
    rd_cycle[16855] = 1'b0;  wr_cycle[16855] = 1'b0;  addr_rom[16855]='h00000000;  wr_data_rom[16855]='h00000000;
    rd_cycle[16856] = 1'b0;  wr_cycle[16856] = 1'b0;  addr_rom[16856]='h00000000;  wr_data_rom[16856]='h00000000;
    rd_cycle[16857] = 1'b0;  wr_cycle[16857] = 1'b0;  addr_rom[16857]='h00000000;  wr_data_rom[16857]='h00000000;
    rd_cycle[16858] = 1'b0;  wr_cycle[16858] = 1'b0;  addr_rom[16858]='h00000000;  wr_data_rom[16858]='h00000000;
    rd_cycle[16859] = 1'b0;  wr_cycle[16859] = 1'b0;  addr_rom[16859]='h00000000;  wr_data_rom[16859]='h00000000;
    rd_cycle[16860] = 1'b0;  wr_cycle[16860] = 1'b0;  addr_rom[16860]='h00000000;  wr_data_rom[16860]='h00000000;
    rd_cycle[16861] = 1'b0;  wr_cycle[16861] = 1'b0;  addr_rom[16861]='h00000000;  wr_data_rom[16861]='h00000000;
    rd_cycle[16862] = 1'b0;  wr_cycle[16862] = 1'b0;  addr_rom[16862]='h00000000;  wr_data_rom[16862]='h00000000;
    rd_cycle[16863] = 1'b0;  wr_cycle[16863] = 1'b0;  addr_rom[16863]='h00000000;  wr_data_rom[16863]='h00000000;
    rd_cycle[16864] = 1'b0;  wr_cycle[16864] = 1'b0;  addr_rom[16864]='h00000000;  wr_data_rom[16864]='h00000000;
    rd_cycle[16865] = 1'b0;  wr_cycle[16865] = 1'b0;  addr_rom[16865]='h00000000;  wr_data_rom[16865]='h00000000;
    rd_cycle[16866] = 1'b0;  wr_cycle[16866] = 1'b0;  addr_rom[16866]='h00000000;  wr_data_rom[16866]='h00000000;
    rd_cycle[16867] = 1'b0;  wr_cycle[16867] = 1'b0;  addr_rom[16867]='h00000000;  wr_data_rom[16867]='h00000000;
    rd_cycle[16868] = 1'b0;  wr_cycle[16868] = 1'b0;  addr_rom[16868]='h00000000;  wr_data_rom[16868]='h00000000;
    rd_cycle[16869] = 1'b0;  wr_cycle[16869] = 1'b0;  addr_rom[16869]='h00000000;  wr_data_rom[16869]='h00000000;
    rd_cycle[16870] = 1'b0;  wr_cycle[16870] = 1'b0;  addr_rom[16870]='h00000000;  wr_data_rom[16870]='h00000000;
    rd_cycle[16871] = 1'b0;  wr_cycle[16871] = 1'b0;  addr_rom[16871]='h00000000;  wr_data_rom[16871]='h00000000;
    rd_cycle[16872] = 1'b0;  wr_cycle[16872] = 1'b0;  addr_rom[16872]='h00000000;  wr_data_rom[16872]='h00000000;
    rd_cycle[16873] = 1'b0;  wr_cycle[16873] = 1'b0;  addr_rom[16873]='h00000000;  wr_data_rom[16873]='h00000000;
    rd_cycle[16874] = 1'b0;  wr_cycle[16874] = 1'b0;  addr_rom[16874]='h00000000;  wr_data_rom[16874]='h00000000;
    rd_cycle[16875] = 1'b0;  wr_cycle[16875] = 1'b0;  addr_rom[16875]='h00000000;  wr_data_rom[16875]='h00000000;
    rd_cycle[16876] = 1'b0;  wr_cycle[16876] = 1'b0;  addr_rom[16876]='h00000000;  wr_data_rom[16876]='h00000000;
    rd_cycle[16877] = 1'b0;  wr_cycle[16877] = 1'b0;  addr_rom[16877]='h00000000;  wr_data_rom[16877]='h00000000;
    rd_cycle[16878] = 1'b0;  wr_cycle[16878] = 1'b0;  addr_rom[16878]='h00000000;  wr_data_rom[16878]='h00000000;
    rd_cycle[16879] = 1'b0;  wr_cycle[16879] = 1'b0;  addr_rom[16879]='h00000000;  wr_data_rom[16879]='h00000000;
    rd_cycle[16880] = 1'b0;  wr_cycle[16880] = 1'b0;  addr_rom[16880]='h00000000;  wr_data_rom[16880]='h00000000;
    rd_cycle[16881] = 1'b0;  wr_cycle[16881] = 1'b0;  addr_rom[16881]='h00000000;  wr_data_rom[16881]='h00000000;
    rd_cycle[16882] = 1'b0;  wr_cycle[16882] = 1'b0;  addr_rom[16882]='h00000000;  wr_data_rom[16882]='h00000000;
    rd_cycle[16883] = 1'b0;  wr_cycle[16883] = 1'b0;  addr_rom[16883]='h00000000;  wr_data_rom[16883]='h00000000;
    rd_cycle[16884] = 1'b0;  wr_cycle[16884] = 1'b0;  addr_rom[16884]='h00000000;  wr_data_rom[16884]='h00000000;
    rd_cycle[16885] = 1'b0;  wr_cycle[16885] = 1'b0;  addr_rom[16885]='h00000000;  wr_data_rom[16885]='h00000000;
    rd_cycle[16886] = 1'b0;  wr_cycle[16886] = 1'b0;  addr_rom[16886]='h00000000;  wr_data_rom[16886]='h00000000;
    rd_cycle[16887] = 1'b0;  wr_cycle[16887] = 1'b0;  addr_rom[16887]='h00000000;  wr_data_rom[16887]='h00000000;
    rd_cycle[16888] = 1'b0;  wr_cycle[16888] = 1'b0;  addr_rom[16888]='h00000000;  wr_data_rom[16888]='h00000000;
    rd_cycle[16889] = 1'b0;  wr_cycle[16889] = 1'b0;  addr_rom[16889]='h00000000;  wr_data_rom[16889]='h00000000;
    rd_cycle[16890] = 1'b0;  wr_cycle[16890] = 1'b0;  addr_rom[16890]='h00000000;  wr_data_rom[16890]='h00000000;
    rd_cycle[16891] = 1'b0;  wr_cycle[16891] = 1'b0;  addr_rom[16891]='h00000000;  wr_data_rom[16891]='h00000000;
    rd_cycle[16892] = 1'b0;  wr_cycle[16892] = 1'b0;  addr_rom[16892]='h00000000;  wr_data_rom[16892]='h00000000;
    rd_cycle[16893] = 1'b0;  wr_cycle[16893] = 1'b0;  addr_rom[16893]='h00000000;  wr_data_rom[16893]='h00000000;
    rd_cycle[16894] = 1'b0;  wr_cycle[16894] = 1'b0;  addr_rom[16894]='h00000000;  wr_data_rom[16894]='h00000000;
    rd_cycle[16895] = 1'b0;  wr_cycle[16895] = 1'b0;  addr_rom[16895]='h00000000;  wr_data_rom[16895]='h00000000;
    rd_cycle[16896] = 1'b0;  wr_cycle[16896] = 1'b0;  addr_rom[16896]='h00000000;  wr_data_rom[16896]='h00000000;
    rd_cycle[16897] = 1'b0;  wr_cycle[16897] = 1'b0;  addr_rom[16897]='h00000000;  wr_data_rom[16897]='h00000000;
    rd_cycle[16898] = 1'b0;  wr_cycle[16898] = 1'b0;  addr_rom[16898]='h00000000;  wr_data_rom[16898]='h00000000;
    rd_cycle[16899] = 1'b0;  wr_cycle[16899] = 1'b0;  addr_rom[16899]='h00000000;  wr_data_rom[16899]='h00000000;
    rd_cycle[16900] = 1'b0;  wr_cycle[16900] = 1'b0;  addr_rom[16900]='h00000000;  wr_data_rom[16900]='h00000000;
    rd_cycle[16901] = 1'b0;  wr_cycle[16901] = 1'b0;  addr_rom[16901]='h00000000;  wr_data_rom[16901]='h00000000;
    rd_cycle[16902] = 1'b0;  wr_cycle[16902] = 1'b0;  addr_rom[16902]='h00000000;  wr_data_rom[16902]='h00000000;
    rd_cycle[16903] = 1'b0;  wr_cycle[16903] = 1'b0;  addr_rom[16903]='h00000000;  wr_data_rom[16903]='h00000000;
    rd_cycle[16904] = 1'b0;  wr_cycle[16904] = 1'b0;  addr_rom[16904]='h00000000;  wr_data_rom[16904]='h00000000;
    rd_cycle[16905] = 1'b0;  wr_cycle[16905] = 1'b0;  addr_rom[16905]='h00000000;  wr_data_rom[16905]='h00000000;
    rd_cycle[16906] = 1'b0;  wr_cycle[16906] = 1'b0;  addr_rom[16906]='h00000000;  wr_data_rom[16906]='h00000000;
    rd_cycle[16907] = 1'b0;  wr_cycle[16907] = 1'b0;  addr_rom[16907]='h00000000;  wr_data_rom[16907]='h00000000;
    rd_cycle[16908] = 1'b0;  wr_cycle[16908] = 1'b0;  addr_rom[16908]='h00000000;  wr_data_rom[16908]='h00000000;
    rd_cycle[16909] = 1'b0;  wr_cycle[16909] = 1'b0;  addr_rom[16909]='h00000000;  wr_data_rom[16909]='h00000000;
    rd_cycle[16910] = 1'b0;  wr_cycle[16910] = 1'b0;  addr_rom[16910]='h00000000;  wr_data_rom[16910]='h00000000;
    rd_cycle[16911] = 1'b0;  wr_cycle[16911] = 1'b0;  addr_rom[16911]='h00000000;  wr_data_rom[16911]='h00000000;
    rd_cycle[16912] = 1'b0;  wr_cycle[16912] = 1'b0;  addr_rom[16912]='h00000000;  wr_data_rom[16912]='h00000000;
    rd_cycle[16913] = 1'b0;  wr_cycle[16913] = 1'b0;  addr_rom[16913]='h00000000;  wr_data_rom[16913]='h00000000;
    rd_cycle[16914] = 1'b0;  wr_cycle[16914] = 1'b0;  addr_rom[16914]='h00000000;  wr_data_rom[16914]='h00000000;
    rd_cycle[16915] = 1'b0;  wr_cycle[16915] = 1'b0;  addr_rom[16915]='h00000000;  wr_data_rom[16915]='h00000000;
    rd_cycle[16916] = 1'b0;  wr_cycle[16916] = 1'b0;  addr_rom[16916]='h00000000;  wr_data_rom[16916]='h00000000;
    rd_cycle[16917] = 1'b0;  wr_cycle[16917] = 1'b0;  addr_rom[16917]='h00000000;  wr_data_rom[16917]='h00000000;
    rd_cycle[16918] = 1'b0;  wr_cycle[16918] = 1'b0;  addr_rom[16918]='h00000000;  wr_data_rom[16918]='h00000000;
    rd_cycle[16919] = 1'b0;  wr_cycle[16919] = 1'b0;  addr_rom[16919]='h00000000;  wr_data_rom[16919]='h00000000;
    rd_cycle[16920] = 1'b0;  wr_cycle[16920] = 1'b0;  addr_rom[16920]='h00000000;  wr_data_rom[16920]='h00000000;
    rd_cycle[16921] = 1'b0;  wr_cycle[16921] = 1'b0;  addr_rom[16921]='h00000000;  wr_data_rom[16921]='h00000000;
    rd_cycle[16922] = 1'b0;  wr_cycle[16922] = 1'b0;  addr_rom[16922]='h00000000;  wr_data_rom[16922]='h00000000;
    rd_cycle[16923] = 1'b0;  wr_cycle[16923] = 1'b0;  addr_rom[16923]='h00000000;  wr_data_rom[16923]='h00000000;
    rd_cycle[16924] = 1'b0;  wr_cycle[16924] = 1'b0;  addr_rom[16924]='h00000000;  wr_data_rom[16924]='h00000000;
    rd_cycle[16925] = 1'b0;  wr_cycle[16925] = 1'b0;  addr_rom[16925]='h00000000;  wr_data_rom[16925]='h00000000;
    rd_cycle[16926] = 1'b0;  wr_cycle[16926] = 1'b0;  addr_rom[16926]='h00000000;  wr_data_rom[16926]='h00000000;
    rd_cycle[16927] = 1'b0;  wr_cycle[16927] = 1'b0;  addr_rom[16927]='h00000000;  wr_data_rom[16927]='h00000000;
    rd_cycle[16928] = 1'b0;  wr_cycle[16928] = 1'b0;  addr_rom[16928]='h00000000;  wr_data_rom[16928]='h00000000;
    rd_cycle[16929] = 1'b0;  wr_cycle[16929] = 1'b0;  addr_rom[16929]='h00000000;  wr_data_rom[16929]='h00000000;
    rd_cycle[16930] = 1'b0;  wr_cycle[16930] = 1'b0;  addr_rom[16930]='h00000000;  wr_data_rom[16930]='h00000000;
    rd_cycle[16931] = 1'b0;  wr_cycle[16931] = 1'b0;  addr_rom[16931]='h00000000;  wr_data_rom[16931]='h00000000;
    rd_cycle[16932] = 1'b0;  wr_cycle[16932] = 1'b0;  addr_rom[16932]='h00000000;  wr_data_rom[16932]='h00000000;
    rd_cycle[16933] = 1'b0;  wr_cycle[16933] = 1'b0;  addr_rom[16933]='h00000000;  wr_data_rom[16933]='h00000000;
    rd_cycle[16934] = 1'b0;  wr_cycle[16934] = 1'b0;  addr_rom[16934]='h00000000;  wr_data_rom[16934]='h00000000;
    rd_cycle[16935] = 1'b0;  wr_cycle[16935] = 1'b0;  addr_rom[16935]='h00000000;  wr_data_rom[16935]='h00000000;
    rd_cycle[16936] = 1'b0;  wr_cycle[16936] = 1'b0;  addr_rom[16936]='h00000000;  wr_data_rom[16936]='h00000000;
    rd_cycle[16937] = 1'b0;  wr_cycle[16937] = 1'b0;  addr_rom[16937]='h00000000;  wr_data_rom[16937]='h00000000;
    rd_cycle[16938] = 1'b0;  wr_cycle[16938] = 1'b0;  addr_rom[16938]='h00000000;  wr_data_rom[16938]='h00000000;
    rd_cycle[16939] = 1'b0;  wr_cycle[16939] = 1'b0;  addr_rom[16939]='h00000000;  wr_data_rom[16939]='h00000000;
    rd_cycle[16940] = 1'b0;  wr_cycle[16940] = 1'b0;  addr_rom[16940]='h00000000;  wr_data_rom[16940]='h00000000;
    rd_cycle[16941] = 1'b0;  wr_cycle[16941] = 1'b0;  addr_rom[16941]='h00000000;  wr_data_rom[16941]='h00000000;
    rd_cycle[16942] = 1'b0;  wr_cycle[16942] = 1'b0;  addr_rom[16942]='h00000000;  wr_data_rom[16942]='h00000000;
    rd_cycle[16943] = 1'b0;  wr_cycle[16943] = 1'b0;  addr_rom[16943]='h00000000;  wr_data_rom[16943]='h00000000;
    rd_cycle[16944] = 1'b0;  wr_cycle[16944] = 1'b0;  addr_rom[16944]='h00000000;  wr_data_rom[16944]='h00000000;
    rd_cycle[16945] = 1'b0;  wr_cycle[16945] = 1'b0;  addr_rom[16945]='h00000000;  wr_data_rom[16945]='h00000000;
    rd_cycle[16946] = 1'b0;  wr_cycle[16946] = 1'b0;  addr_rom[16946]='h00000000;  wr_data_rom[16946]='h00000000;
    rd_cycle[16947] = 1'b0;  wr_cycle[16947] = 1'b0;  addr_rom[16947]='h00000000;  wr_data_rom[16947]='h00000000;
    rd_cycle[16948] = 1'b0;  wr_cycle[16948] = 1'b0;  addr_rom[16948]='h00000000;  wr_data_rom[16948]='h00000000;
    rd_cycle[16949] = 1'b0;  wr_cycle[16949] = 1'b0;  addr_rom[16949]='h00000000;  wr_data_rom[16949]='h00000000;
    rd_cycle[16950] = 1'b0;  wr_cycle[16950] = 1'b0;  addr_rom[16950]='h00000000;  wr_data_rom[16950]='h00000000;
    rd_cycle[16951] = 1'b0;  wr_cycle[16951] = 1'b0;  addr_rom[16951]='h00000000;  wr_data_rom[16951]='h00000000;
    rd_cycle[16952] = 1'b0;  wr_cycle[16952] = 1'b0;  addr_rom[16952]='h00000000;  wr_data_rom[16952]='h00000000;
    rd_cycle[16953] = 1'b0;  wr_cycle[16953] = 1'b0;  addr_rom[16953]='h00000000;  wr_data_rom[16953]='h00000000;
    rd_cycle[16954] = 1'b0;  wr_cycle[16954] = 1'b0;  addr_rom[16954]='h00000000;  wr_data_rom[16954]='h00000000;
    rd_cycle[16955] = 1'b0;  wr_cycle[16955] = 1'b0;  addr_rom[16955]='h00000000;  wr_data_rom[16955]='h00000000;
    rd_cycle[16956] = 1'b0;  wr_cycle[16956] = 1'b0;  addr_rom[16956]='h00000000;  wr_data_rom[16956]='h00000000;
    rd_cycle[16957] = 1'b0;  wr_cycle[16957] = 1'b0;  addr_rom[16957]='h00000000;  wr_data_rom[16957]='h00000000;
    rd_cycle[16958] = 1'b0;  wr_cycle[16958] = 1'b0;  addr_rom[16958]='h00000000;  wr_data_rom[16958]='h00000000;
    rd_cycle[16959] = 1'b0;  wr_cycle[16959] = 1'b0;  addr_rom[16959]='h00000000;  wr_data_rom[16959]='h00000000;
    rd_cycle[16960] = 1'b0;  wr_cycle[16960] = 1'b0;  addr_rom[16960]='h00000000;  wr_data_rom[16960]='h00000000;
    rd_cycle[16961] = 1'b0;  wr_cycle[16961] = 1'b0;  addr_rom[16961]='h00000000;  wr_data_rom[16961]='h00000000;
    rd_cycle[16962] = 1'b0;  wr_cycle[16962] = 1'b0;  addr_rom[16962]='h00000000;  wr_data_rom[16962]='h00000000;
    rd_cycle[16963] = 1'b0;  wr_cycle[16963] = 1'b0;  addr_rom[16963]='h00000000;  wr_data_rom[16963]='h00000000;
    rd_cycle[16964] = 1'b0;  wr_cycle[16964] = 1'b0;  addr_rom[16964]='h00000000;  wr_data_rom[16964]='h00000000;
    rd_cycle[16965] = 1'b0;  wr_cycle[16965] = 1'b0;  addr_rom[16965]='h00000000;  wr_data_rom[16965]='h00000000;
    rd_cycle[16966] = 1'b0;  wr_cycle[16966] = 1'b0;  addr_rom[16966]='h00000000;  wr_data_rom[16966]='h00000000;
    rd_cycle[16967] = 1'b0;  wr_cycle[16967] = 1'b0;  addr_rom[16967]='h00000000;  wr_data_rom[16967]='h00000000;
    rd_cycle[16968] = 1'b0;  wr_cycle[16968] = 1'b0;  addr_rom[16968]='h00000000;  wr_data_rom[16968]='h00000000;
    rd_cycle[16969] = 1'b0;  wr_cycle[16969] = 1'b0;  addr_rom[16969]='h00000000;  wr_data_rom[16969]='h00000000;
    rd_cycle[16970] = 1'b0;  wr_cycle[16970] = 1'b0;  addr_rom[16970]='h00000000;  wr_data_rom[16970]='h00000000;
    rd_cycle[16971] = 1'b0;  wr_cycle[16971] = 1'b0;  addr_rom[16971]='h00000000;  wr_data_rom[16971]='h00000000;
    rd_cycle[16972] = 1'b0;  wr_cycle[16972] = 1'b0;  addr_rom[16972]='h00000000;  wr_data_rom[16972]='h00000000;
    rd_cycle[16973] = 1'b0;  wr_cycle[16973] = 1'b0;  addr_rom[16973]='h00000000;  wr_data_rom[16973]='h00000000;
    rd_cycle[16974] = 1'b0;  wr_cycle[16974] = 1'b0;  addr_rom[16974]='h00000000;  wr_data_rom[16974]='h00000000;
    rd_cycle[16975] = 1'b0;  wr_cycle[16975] = 1'b0;  addr_rom[16975]='h00000000;  wr_data_rom[16975]='h00000000;
    rd_cycle[16976] = 1'b0;  wr_cycle[16976] = 1'b0;  addr_rom[16976]='h00000000;  wr_data_rom[16976]='h00000000;
    rd_cycle[16977] = 1'b0;  wr_cycle[16977] = 1'b0;  addr_rom[16977]='h00000000;  wr_data_rom[16977]='h00000000;
    rd_cycle[16978] = 1'b0;  wr_cycle[16978] = 1'b0;  addr_rom[16978]='h00000000;  wr_data_rom[16978]='h00000000;
    rd_cycle[16979] = 1'b0;  wr_cycle[16979] = 1'b0;  addr_rom[16979]='h00000000;  wr_data_rom[16979]='h00000000;
    rd_cycle[16980] = 1'b0;  wr_cycle[16980] = 1'b0;  addr_rom[16980]='h00000000;  wr_data_rom[16980]='h00000000;
    rd_cycle[16981] = 1'b0;  wr_cycle[16981] = 1'b0;  addr_rom[16981]='h00000000;  wr_data_rom[16981]='h00000000;
    rd_cycle[16982] = 1'b0;  wr_cycle[16982] = 1'b0;  addr_rom[16982]='h00000000;  wr_data_rom[16982]='h00000000;
    rd_cycle[16983] = 1'b0;  wr_cycle[16983] = 1'b0;  addr_rom[16983]='h00000000;  wr_data_rom[16983]='h00000000;
    rd_cycle[16984] = 1'b0;  wr_cycle[16984] = 1'b0;  addr_rom[16984]='h00000000;  wr_data_rom[16984]='h00000000;
    rd_cycle[16985] = 1'b0;  wr_cycle[16985] = 1'b0;  addr_rom[16985]='h00000000;  wr_data_rom[16985]='h00000000;
    rd_cycle[16986] = 1'b0;  wr_cycle[16986] = 1'b0;  addr_rom[16986]='h00000000;  wr_data_rom[16986]='h00000000;
    rd_cycle[16987] = 1'b0;  wr_cycle[16987] = 1'b0;  addr_rom[16987]='h00000000;  wr_data_rom[16987]='h00000000;
    rd_cycle[16988] = 1'b0;  wr_cycle[16988] = 1'b0;  addr_rom[16988]='h00000000;  wr_data_rom[16988]='h00000000;
    rd_cycle[16989] = 1'b0;  wr_cycle[16989] = 1'b0;  addr_rom[16989]='h00000000;  wr_data_rom[16989]='h00000000;
    rd_cycle[16990] = 1'b0;  wr_cycle[16990] = 1'b0;  addr_rom[16990]='h00000000;  wr_data_rom[16990]='h00000000;
    rd_cycle[16991] = 1'b0;  wr_cycle[16991] = 1'b0;  addr_rom[16991]='h00000000;  wr_data_rom[16991]='h00000000;
    rd_cycle[16992] = 1'b0;  wr_cycle[16992] = 1'b0;  addr_rom[16992]='h00000000;  wr_data_rom[16992]='h00000000;
    rd_cycle[16993] = 1'b0;  wr_cycle[16993] = 1'b0;  addr_rom[16993]='h00000000;  wr_data_rom[16993]='h00000000;
    rd_cycle[16994] = 1'b0;  wr_cycle[16994] = 1'b0;  addr_rom[16994]='h00000000;  wr_data_rom[16994]='h00000000;
    rd_cycle[16995] = 1'b0;  wr_cycle[16995] = 1'b0;  addr_rom[16995]='h00000000;  wr_data_rom[16995]='h00000000;
    rd_cycle[16996] = 1'b0;  wr_cycle[16996] = 1'b0;  addr_rom[16996]='h00000000;  wr_data_rom[16996]='h00000000;
    rd_cycle[16997] = 1'b0;  wr_cycle[16997] = 1'b0;  addr_rom[16997]='h00000000;  wr_data_rom[16997]='h00000000;
    rd_cycle[16998] = 1'b0;  wr_cycle[16998] = 1'b0;  addr_rom[16998]='h00000000;  wr_data_rom[16998]='h00000000;
    rd_cycle[16999] = 1'b0;  wr_cycle[16999] = 1'b0;  addr_rom[16999]='h00000000;  wr_data_rom[16999]='h00000000;
    rd_cycle[17000] = 1'b0;  wr_cycle[17000] = 1'b0;  addr_rom[17000]='h00000000;  wr_data_rom[17000]='h00000000;
    rd_cycle[17001] = 1'b0;  wr_cycle[17001] = 1'b0;  addr_rom[17001]='h00000000;  wr_data_rom[17001]='h00000000;
    rd_cycle[17002] = 1'b0;  wr_cycle[17002] = 1'b0;  addr_rom[17002]='h00000000;  wr_data_rom[17002]='h00000000;
    rd_cycle[17003] = 1'b0;  wr_cycle[17003] = 1'b0;  addr_rom[17003]='h00000000;  wr_data_rom[17003]='h00000000;
    rd_cycle[17004] = 1'b0;  wr_cycle[17004] = 1'b0;  addr_rom[17004]='h00000000;  wr_data_rom[17004]='h00000000;
    rd_cycle[17005] = 1'b0;  wr_cycle[17005] = 1'b0;  addr_rom[17005]='h00000000;  wr_data_rom[17005]='h00000000;
    rd_cycle[17006] = 1'b0;  wr_cycle[17006] = 1'b0;  addr_rom[17006]='h00000000;  wr_data_rom[17006]='h00000000;
    rd_cycle[17007] = 1'b0;  wr_cycle[17007] = 1'b0;  addr_rom[17007]='h00000000;  wr_data_rom[17007]='h00000000;
    rd_cycle[17008] = 1'b0;  wr_cycle[17008] = 1'b0;  addr_rom[17008]='h00000000;  wr_data_rom[17008]='h00000000;
    rd_cycle[17009] = 1'b0;  wr_cycle[17009] = 1'b0;  addr_rom[17009]='h00000000;  wr_data_rom[17009]='h00000000;
    rd_cycle[17010] = 1'b0;  wr_cycle[17010] = 1'b0;  addr_rom[17010]='h00000000;  wr_data_rom[17010]='h00000000;
    rd_cycle[17011] = 1'b0;  wr_cycle[17011] = 1'b0;  addr_rom[17011]='h00000000;  wr_data_rom[17011]='h00000000;
    rd_cycle[17012] = 1'b0;  wr_cycle[17012] = 1'b0;  addr_rom[17012]='h00000000;  wr_data_rom[17012]='h00000000;
    rd_cycle[17013] = 1'b0;  wr_cycle[17013] = 1'b0;  addr_rom[17013]='h00000000;  wr_data_rom[17013]='h00000000;
    rd_cycle[17014] = 1'b0;  wr_cycle[17014] = 1'b0;  addr_rom[17014]='h00000000;  wr_data_rom[17014]='h00000000;
    rd_cycle[17015] = 1'b0;  wr_cycle[17015] = 1'b0;  addr_rom[17015]='h00000000;  wr_data_rom[17015]='h00000000;
    rd_cycle[17016] = 1'b0;  wr_cycle[17016] = 1'b0;  addr_rom[17016]='h00000000;  wr_data_rom[17016]='h00000000;
    rd_cycle[17017] = 1'b0;  wr_cycle[17017] = 1'b0;  addr_rom[17017]='h00000000;  wr_data_rom[17017]='h00000000;
    rd_cycle[17018] = 1'b0;  wr_cycle[17018] = 1'b0;  addr_rom[17018]='h00000000;  wr_data_rom[17018]='h00000000;
    rd_cycle[17019] = 1'b0;  wr_cycle[17019] = 1'b0;  addr_rom[17019]='h00000000;  wr_data_rom[17019]='h00000000;
    rd_cycle[17020] = 1'b0;  wr_cycle[17020] = 1'b0;  addr_rom[17020]='h00000000;  wr_data_rom[17020]='h00000000;
    rd_cycle[17021] = 1'b0;  wr_cycle[17021] = 1'b0;  addr_rom[17021]='h00000000;  wr_data_rom[17021]='h00000000;
    rd_cycle[17022] = 1'b0;  wr_cycle[17022] = 1'b0;  addr_rom[17022]='h00000000;  wr_data_rom[17022]='h00000000;
    rd_cycle[17023] = 1'b0;  wr_cycle[17023] = 1'b0;  addr_rom[17023]='h00000000;  wr_data_rom[17023]='h00000000;
    rd_cycle[17024] = 1'b0;  wr_cycle[17024] = 1'b0;  addr_rom[17024]='h00000000;  wr_data_rom[17024]='h00000000;
    rd_cycle[17025] = 1'b0;  wr_cycle[17025] = 1'b0;  addr_rom[17025]='h00000000;  wr_data_rom[17025]='h00000000;
    rd_cycle[17026] = 1'b0;  wr_cycle[17026] = 1'b0;  addr_rom[17026]='h00000000;  wr_data_rom[17026]='h00000000;
    rd_cycle[17027] = 1'b0;  wr_cycle[17027] = 1'b0;  addr_rom[17027]='h00000000;  wr_data_rom[17027]='h00000000;
    rd_cycle[17028] = 1'b0;  wr_cycle[17028] = 1'b0;  addr_rom[17028]='h00000000;  wr_data_rom[17028]='h00000000;
    rd_cycle[17029] = 1'b0;  wr_cycle[17029] = 1'b0;  addr_rom[17029]='h00000000;  wr_data_rom[17029]='h00000000;
    rd_cycle[17030] = 1'b0;  wr_cycle[17030] = 1'b0;  addr_rom[17030]='h00000000;  wr_data_rom[17030]='h00000000;
    rd_cycle[17031] = 1'b0;  wr_cycle[17031] = 1'b0;  addr_rom[17031]='h00000000;  wr_data_rom[17031]='h00000000;
    rd_cycle[17032] = 1'b0;  wr_cycle[17032] = 1'b0;  addr_rom[17032]='h00000000;  wr_data_rom[17032]='h00000000;
    rd_cycle[17033] = 1'b0;  wr_cycle[17033] = 1'b0;  addr_rom[17033]='h00000000;  wr_data_rom[17033]='h00000000;
    rd_cycle[17034] = 1'b0;  wr_cycle[17034] = 1'b0;  addr_rom[17034]='h00000000;  wr_data_rom[17034]='h00000000;
    rd_cycle[17035] = 1'b0;  wr_cycle[17035] = 1'b0;  addr_rom[17035]='h00000000;  wr_data_rom[17035]='h00000000;
    rd_cycle[17036] = 1'b0;  wr_cycle[17036] = 1'b0;  addr_rom[17036]='h00000000;  wr_data_rom[17036]='h00000000;
    rd_cycle[17037] = 1'b0;  wr_cycle[17037] = 1'b0;  addr_rom[17037]='h00000000;  wr_data_rom[17037]='h00000000;
    rd_cycle[17038] = 1'b0;  wr_cycle[17038] = 1'b0;  addr_rom[17038]='h00000000;  wr_data_rom[17038]='h00000000;
    rd_cycle[17039] = 1'b0;  wr_cycle[17039] = 1'b0;  addr_rom[17039]='h00000000;  wr_data_rom[17039]='h00000000;
    rd_cycle[17040] = 1'b0;  wr_cycle[17040] = 1'b0;  addr_rom[17040]='h00000000;  wr_data_rom[17040]='h00000000;
    rd_cycle[17041] = 1'b0;  wr_cycle[17041] = 1'b0;  addr_rom[17041]='h00000000;  wr_data_rom[17041]='h00000000;
    rd_cycle[17042] = 1'b0;  wr_cycle[17042] = 1'b0;  addr_rom[17042]='h00000000;  wr_data_rom[17042]='h00000000;
    rd_cycle[17043] = 1'b0;  wr_cycle[17043] = 1'b0;  addr_rom[17043]='h00000000;  wr_data_rom[17043]='h00000000;
    rd_cycle[17044] = 1'b0;  wr_cycle[17044] = 1'b0;  addr_rom[17044]='h00000000;  wr_data_rom[17044]='h00000000;
    rd_cycle[17045] = 1'b0;  wr_cycle[17045] = 1'b0;  addr_rom[17045]='h00000000;  wr_data_rom[17045]='h00000000;
    rd_cycle[17046] = 1'b0;  wr_cycle[17046] = 1'b0;  addr_rom[17046]='h00000000;  wr_data_rom[17046]='h00000000;
    rd_cycle[17047] = 1'b0;  wr_cycle[17047] = 1'b0;  addr_rom[17047]='h00000000;  wr_data_rom[17047]='h00000000;
    rd_cycle[17048] = 1'b0;  wr_cycle[17048] = 1'b0;  addr_rom[17048]='h00000000;  wr_data_rom[17048]='h00000000;
    rd_cycle[17049] = 1'b0;  wr_cycle[17049] = 1'b0;  addr_rom[17049]='h00000000;  wr_data_rom[17049]='h00000000;
    rd_cycle[17050] = 1'b0;  wr_cycle[17050] = 1'b0;  addr_rom[17050]='h00000000;  wr_data_rom[17050]='h00000000;
    rd_cycle[17051] = 1'b0;  wr_cycle[17051] = 1'b0;  addr_rom[17051]='h00000000;  wr_data_rom[17051]='h00000000;
    rd_cycle[17052] = 1'b0;  wr_cycle[17052] = 1'b0;  addr_rom[17052]='h00000000;  wr_data_rom[17052]='h00000000;
    rd_cycle[17053] = 1'b0;  wr_cycle[17053] = 1'b0;  addr_rom[17053]='h00000000;  wr_data_rom[17053]='h00000000;
    rd_cycle[17054] = 1'b0;  wr_cycle[17054] = 1'b0;  addr_rom[17054]='h00000000;  wr_data_rom[17054]='h00000000;
    rd_cycle[17055] = 1'b0;  wr_cycle[17055] = 1'b0;  addr_rom[17055]='h00000000;  wr_data_rom[17055]='h00000000;
    rd_cycle[17056] = 1'b0;  wr_cycle[17056] = 1'b0;  addr_rom[17056]='h00000000;  wr_data_rom[17056]='h00000000;
    rd_cycle[17057] = 1'b0;  wr_cycle[17057] = 1'b0;  addr_rom[17057]='h00000000;  wr_data_rom[17057]='h00000000;
    rd_cycle[17058] = 1'b0;  wr_cycle[17058] = 1'b0;  addr_rom[17058]='h00000000;  wr_data_rom[17058]='h00000000;
    rd_cycle[17059] = 1'b0;  wr_cycle[17059] = 1'b0;  addr_rom[17059]='h00000000;  wr_data_rom[17059]='h00000000;
    rd_cycle[17060] = 1'b0;  wr_cycle[17060] = 1'b0;  addr_rom[17060]='h00000000;  wr_data_rom[17060]='h00000000;
    rd_cycle[17061] = 1'b0;  wr_cycle[17061] = 1'b0;  addr_rom[17061]='h00000000;  wr_data_rom[17061]='h00000000;
    rd_cycle[17062] = 1'b0;  wr_cycle[17062] = 1'b0;  addr_rom[17062]='h00000000;  wr_data_rom[17062]='h00000000;
    rd_cycle[17063] = 1'b0;  wr_cycle[17063] = 1'b0;  addr_rom[17063]='h00000000;  wr_data_rom[17063]='h00000000;
    rd_cycle[17064] = 1'b0;  wr_cycle[17064] = 1'b0;  addr_rom[17064]='h00000000;  wr_data_rom[17064]='h00000000;
    rd_cycle[17065] = 1'b0;  wr_cycle[17065] = 1'b0;  addr_rom[17065]='h00000000;  wr_data_rom[17065]='h00000000;
    rd_cycle[17066] = 1'b0;  wr_cycle[17066] = 1'b0;  addr_rom[17066]='h00000000;  wr_data_rom[17066]='h00000000;
    rd_cycle[17067] = 1'b0;  wr_cycle[17067] = 1'b0;  addr_rom[17067]='h00000000;  wr_data_rom[17067]='h00000000;
    rd_cycle[17068] = 1'b0;  wr_cycle[17068] = 1'b0;  addr_rom[17068]='h00000000;  wr_data_rom[17068]='h00000000;
    rd_cycle[17069] = 1'b0;  wr_cycle[17069] = 1'b0;  addr_rom[17069]='h00000000;  wr_data_rom[17069]='h00000000;
    rd_cycle[17070] = 1'b0;  wr_cycle[17070] = 1'b0;  addr_rom[17070]='h00000000;  wr_data_rom[17070]='h00000000;
    rd_cycle[17071] = 1'b0;  wr_cycle[17071] = 1'b0;  addr_rom[17071]='h00000000;  wr_data_rom[17071]='h00000000;
    rd_cycle[17072] = 1'b0;  wr_cycle[17072] = 1'b0;  addr_rom[17072]='h00000000;  wr_data_rom[17072]='h00000000;
    rd_cycle[17073] = 1'b0;  wr_cycle[17073] = 1'b0;  addr_rom[17073]='h00000000;  wr_data_rom[17073]='h00000000;
    rd_cycle[17074] = 1'b0;  wr_cycle[17074] = 1'b0;  addr_rom[17074]='h00000000;  wr_data_rom[17074]='h00000000;
    rd_cycle[17075] = 1'b0;  wr_cycle[17075] = 1'b0;  addr_rom[17075]='h00000000;  wr_data_rom[17075]='h00000000;
    rd_cycle[17076] = 1'b0;  wr_cycle[17076] = 1'b0;  addr_rom[17076]='h00000000;  wr_data_rom[17076]='h00000000;
    rd_cycle[17077] = 1'b0;  wr_cycle[17077] = 1'b0;  addr_rom[17077]='h00000000;  wr_data_rom[17077]='h00000000;
    rd_cycle[17078] = 1'b0;  wr_cycle[17078] = 1'b0;  addr_rom[17078]='h00000000;  wr_data_rom[17078]='h00000000;
    rd_cycle[17079] = 1'b0;  wr_cycle[17079] = 1'b0;  addr_rom[17079]='h00000000;  wr_data_rom[17079]='h00000000;
    rd_cycle[17080] = 1'b0;  wr_cycle[17080] = 1'b0;  addr_rom[17080]='h00000000;  wr_data_rom[17080]='h00000000;
    rd_cycle[17081] = 1'b0;  wr_cycle[17081] = 1'b0;  addr_rom[17081]='h00000000;  wr_data_rom[17081]='h00000000;
    rd_cycle[17082] = 1'b0;  wr_cycle[17082] = 1'b0;  addr_rom[17082]='h00000000;  wr_data_rom[17082]='h00000000;
    rd_cycle[17083] = 1'b0;  wr_cycle[17083] = 1'b0;  addr_rom[17083]='h00000000;  wr_data_rom[17083]='h00000000;
    rd_cycle[17084] = 1'b0;  wr_cycle[17084] = 1'b0;  addr_rom[17084]='h00000000;  wr_data_rom[17084]='h00000000;
    rd_cycle[17085] = 1'b0;  wr_cycle[17085] = 1'b0;  addr_rom[17085]='h00000000;  wr_data_rom[17085]='h00000000;
    rd_cycle[17086] = 1'b0;  wr_cycle[17086] = 1'b0;  addr_rom[17086]='h00000000;  wr_data_rom[17086]='h00000000;
    rd_cycle[17087] = 1'b0;  wr_cycle[17087] = 1'b0;  addr_rom[17087]='h00000000;  wr_data_rom[17087]='h00000000;
    rd_cycle[17088] = 1'b0;  wr_cycle[17088] = 1'b0;  addr_rom[17088]='h00000000;  wr_data_rom[17088]='h00000000;
    rd_cycle[17089] = 1'b0;  wr_cycle[17089] = 1'b0;  addr_rom[17089]='h00000000;  wr_data_rom[17089]='h00000000;
    rd_cycle[17090] = 1'b0;  wr_cycle[17090] = 1'b0;  addr_rom[17090]='h00000000;  wr_data_rom[17090]='h00000000;
    rd_cycle[17091] = 1'b0;  wr_cycle[17091] = 1'b0;  addr_rom[17091]='h00000000;  wr_data_rom[17091]='h00000000;
    rd_cycle[17092] = 1'b0;  wr_cycle[17092] = 1'b0;  addr_rom[17092]='h00000000;  wr_data_rom[17092]='h00000000;
    rd_cycle[17093] = 1'b0;  wr_cycle[17093] = 1'b0;  addr_rom[17093]='h00000000;  wr_data_rom[17093]='h00000000;
    rd_cycle[17094] = 1'b0;  wr_cycle[17094] = 1'b0;  addr_rom[17094]='h00000000;  wr_data_rom[17094]='h00000000;
    rd_cycle[17095] = 1'b0;  wr_cycle[17095] = 1'b0;  addr_rom[17095]='h00000000;  wr_data_rom[17095]='h00000000;
    rd_cycle[17096] = 1'b0;  wr_cycle[17096] = 1'b0;  addr_rom[17096]='h00000000;  wr_data_rom[17096]='h00000000;
    rd_cycle[17097] = 1'b0;  wr_cycle[17097] = 1'b0;  addr_rom[17097]='h00000000;  wr_data_rom[17097]='h00000000;
    rd_cycle[17098] = 1'b0;  wr_cycle[17098] = 1'b0;  addr_rom[17098]='h00000000;  wr_data_rom[17098]='h00000000;
    rd_cycle[17099] = 1'b0;  wr_cycle[17099] = 1'b0;  addr_rom[17099]='h00000000;  wr_data_rom[17099]='h00000000;
    rd_cycle[17100] = 1'b0;  wr_cycle[17100] = 1'b0;  addr_rom[17100]='h00000000;  wr_data_rom[17100]='h00000000;
    rd_cycle[17101] = 1'b0;  wr_cycle[17101] = 1'b0;  addr_rom[17101]='h00000000;  wr_data_rom[17101]='h00000000;
    rd_cycle[17102] = 1'b0;  wr_cycle[17102] = 1'b0;  addr_rom[17102]='h00000000;  wr_data_rom[17102]='h00000000;
    rd_cycle[17103] = 1'b0;  wr_cycle[17103] = 1'b0;  addr_rom[17103]='h00000000;  wr_data_rom[17103]='h00000000;
    rd_cycle[17104] = 1'b0;  wr_cycle[17104] = 1'b0;  addr_rom[17104]='h00000000;  wr_data_rom[17104]='h00000000;
    rd_cycle[17105] = 1'b0;  wr_cycle[17105] = 1'b0;  addr_rom[17105]='h00000000;  wr_data_rom[17105]='h00000000;
    rd_cycle[17106] = 1'b0;  wr_cycle[17106] = 1'b0;  addr_rom[17106]='h00000000;  wr_data_rom[17106]='h00000000;
    rd_cycle[17107] = 1'b0;  wr_cycle[17107] = 1'b0;  addr_rom[17107]='h00000000;  wr_data_rom[17107]='h00000000;
    rd_cycle[17108] = 1'b0;  wr_cycle[17108] = 1'b0;  addr_rom[17108]='h00000000;  wr_data_rom[17108]='h00000000;
    rd_cycle[17109] = 1'b0;  wr_cycle[17109] = 1'b0;  addr_rom[17109]='h00000000;  wr_data_rom[17109]='h00000000;
    rd_cycle[17110] = 1'b0;  wr_cycle[17110] = 1'b0;  addr_rom[17110]='h00000000;  wr_data_rom[17110]='h00000000;
    rd_cycle[17111] = 1'b0;  wr_cycle[17111] = 1'b0;  addr_rom[17111]='h00000000;  wr_data_rom[17111]='h00000000;
    rd_cycle[17112] = 1'b0;  wr_cycle[17112] = 1'b0;  addr_rom[17112]='h00000000;  wr_data_rom[17112]='h00000000;
    rd_cycle[17113] = 1'b0;  wr_cycle[17113] = 1'b0;  addr_rom[17113]='h00000000;  wr_data_rom[17113]='h00000000;
    rd_cycle[17114] = 1'b0;  wr_cycle[17114] = 1'b0;  addr_rom[17114]='h00000000;  wr_data_rom[17114]='h00000000;
    rd_cycle[17115] = 1'b0;  wr_cycle[17115] = 1'b0;  addr_rom[17115]='h00000000;  wr_data_rom[17115]='h00000000;
    rd_cycle[17116] = 1'b0;  wr_cycle[17116] = 1'b0;  addr_rom[17116]='h00000000;  wr_data_rom[17116]='h00000000;
    rd_cycle[17117] = 1'b0;  wr_cycle[17117] = 1'b0;  addr_rom[17117]='h00000000;  wr_data_rom[17117]='h00000000;
    rd_cycle[17118] = 1'b0;  wr_cycle[17118] = 1'b0;  addr_rom[17118]='h00000000;  wr_data_rom[17118]='h00000000;
    rd_cycle[17119] = 1'b0;  wr_cycle[17119] = 1'b0;  addr_rom[17119]='h00000000;  wr_data_rom[17119]='h00000000;
    rd_cycle[17120] = 1'b0;  wr_cycle[17120] = 1'b0;  addr_rom[17120]='h00000000;  wr_data_rom[17120]='h00000000;
    rd_cycle[17121] = 1'b0;  wr_cycle[17121] = 1'b0;  addr_rom[17121]='h00000000;  wr_data_rom[17121]='h00000000;
    rd_cycle[17122] = 1'b0;  wr_cycle[17122] = 1'b0;  addr_rom[17122]='h00000000;  wr_data_rom[17122]='h00000000;
    rd_cycle[17123] = 1'b0;  wr_cycle[17123] = 1'b0;  addr_rom[17123]='h00000000;  wr_data_rom[17123]='h00000000;
    rd_cycle[17124] = 1'b0;  wr_cycle[17124] = 1'b0;  addr_rom[17124]='h00000000;  wr_data_rom[17124]='h00000000;
    rd_cycle[17125] = 1'b0;  wr_cycle[17125] = 1'b0;  addr_rom[17125]='h00000000;  wr_data_rom[17125]='h00000000;
    rd_cycle[17126] = 1'b0;  wr_cycle[17126] = 1'b0;  addr_rom[17126]='h00000000;  wr_data_rom[17126]='h00000000;
    rd_cycle[17127] = 1'b0;  wr_cycle[17127] = 1'b0;  addr_rom[17127]='h00000000;  wr_data_rom[17127]='h00000000;
    rd_cycle[17128] = 1'b0;  wr_cycle[17128] = 1'b0;  addr_rom[17128]='h00000000;  wr_data_rom[17128]='h00000000;
    rd_cycle[17129] = 1'b0;  wr_cycle[17129] = 1'b0;  addr_rom[17129]='h00000000;  wr_data_rom[17129]='h00000000;
    rd_cycle[17130] = 1'b0;  wr_cycle[17130] = 1'b0;  addr_rom[17130]='h00000000;  wr_data_rom[17130]='h00000000;
    rd_cycle[17131] = 1'b0;  wr_cycle[17131] = 1'b0;  addr_rom[17131]='h00000000;  wr_data_rom[17131]='h00000000;
    rd_cycle[17132] = 1'b0;  wr_cycle[17132] = 1'b0;  addr_rom[17132]='h00000000;  wr_data_rom[17132]='h00000000;
    rd_cycle[17133] = 1'b0;  wr_cycle[17133] = 1'b0;  addr_rom[17133]='h00000000;  wr_data_rom[17133]='h00000000;
    rd_cycle[17134] = 1'b0;  wr_cycle[17134] = 1'b0;  addr_rom[17134]='h00000000;  wr_data_rom[17134]='h00000000;
    rd_cycle[17135] = 1'b0;  wr_cycle[17135] = 1'b0;  addr_rom[17135]='h00000000;  wr_data_rom[17135]='h00000000;
    rd_cycle[17136] = 1'b0;  wr_cycle[17136] = 1'b0;  addr_rom[17136]='h00000000;  wr_data_rom[17136]='h00000000;
    rd_cycle[17137] = 1'b0;  wr_cycle[17137] = 1'b0;  addr_rom[17137]='h00000000;  wr_data_rom[17137]='h00000000;
    rd_cycle[17138] = 1'b0;  wr_cycle[17138] = 1'b0;  addr_rom[17138]='h00000000;  wr_data_rom[17138]='h00000000;
    rd_cycle[17139] = 1'b0;  wr_cycle[17139] = 1'b0;  addr_rom[17139]='h00000000;  wr_data_rom[17139]='h00000000;
    rd_cycle[17140] = 1'b0;  wr_cycle[17140] = 1'b0;  addr_rom[17140]='h00000000;  wr_data_rom[17140]='h00000000;
    rd_cycle[17141] = 1'b0;  wr_cycle[17141] = 1'b0;  addr_rom[17141]='h00000000;  wr_data_rom[17141]='h00000000;
    rd_cycle[17142] = 1'b0;  wr_cycle[17142] = 1'b0;  addr_rom[17142]='h00000000;  wr_data_rom[17142]='h00000000;
    rd_cycle[17143] = 1'b0;  wr_cycle[17143] = 1'b0;  addr_rom[17143]='h00000000;  wr_data_rom[17143]='h00000000;
    rd_cycle[17144] = 1'b0;  wr_cycle[17144] = 1'b0;  addr_rom[17144]='h00000000;  wr_data_rom[17144]='h00000000;
    rd_cycle[17145] = 1'b0;  wr_cycle[17145] = 1'b0;  addr_rom[17145]='h00000000;  wr_data_rom[17145]='h00000000;
    rd_cycle[17146] = 1'b0;  wr_cycle[17146] = 1'b0;  addr_rom[17146]='h00000000;  wr_data_rom[17146]='h00000000;
    rd_cycle[17147] = 1'b0;  wr_cycle[17147] = 1'b0;  addr_rom[17147]='h00000000;  wr_data_rom[17147]='h00000000;
    rd_cycle[17148] = 1'b0;  wr_cycle[17148] = 1'b0;  addr_rom[17148]='h00000000;  wr_data_rom[17148]='h00000000;
    rd_cycle[17149] = 1'b0;  wr_cycle[17149] = 1'b0;  addr_rom[17149]='h00000000;  wr_data_rom[17149]='h00000000;
    rd_cycle[17150] = 1'b0;  wr_cycle[17150] = 1'b0;  addr_rom[17150]='h00000000;  wr_data_rom[17150]='h00000000;
    rd_cycle[17151] = 1'b0;  wr_cycle[17151] = 1'b0;  addr_rom[17151]='h00000000;  wr_data_rom[17151]='h00000000;
    rd_cycle[17152] = 1'b0;  wr_cycle[17152] = 1'b0;  addr_rom[17152]='h00000000;  wr_data_rom[17152]='h00000000;
    rd_cycle[17153] = 1'b0;  wr_cycle[17153] = 1'b0;  addr_rom[17153]='h00000000;  wr_data_rom[17153]='h00000000;
    rd_cycle[17154] = 1'b0;  wr_cycle[17154] = 1'b0;  addr_rom[17154]='h00000000;  wr_data_rom[17154]='h00000000;
    rd_cycle[17155] = 1'b0;  wr_cycle[17155] = 1'b0;  addr_rom[17155]='h00000000;  wr_data_rom[17155]='h00000000;
    rd_cycle[17156] = 1'b0;  wr_cycle[17156] = 1'b0;  addr_rom[17156]='h00000000;  wr_data_rom[17156]='h00000000;
    rd_cycle[17157] = 1'b0;  wr_cycle[17157] = 1'b0;  addr_rom[17157]='h00000000;  wr_data_rom[17157]='h00000000;
    rd_cycle[17158] = 1'b0;  wr_cycle[17158] = 1'b0;  addr_rom[17158]='h00000000;  wr_data_rom[17158]='h00000000;
    rd_cycle[17159] = 1'b0;  wr_cycle[17159] = 1'b0;  addr_rom[17159]='h00000000;  wr_data_rom[17159]='h00000000;
    rd_cycle[17160] = 1'b0;  wr_cycle[17160] = 1'b0;  addr_rom[17160]='h00000000;  wr_data_rom[17160]='h00000000;
    rd_cycle[17161] = 1'b0;  wr_cycle[17161] = 1'b0;  addr_rom[17161]='h00000000;  wr_data_rom[17161]='h00000000;
    rd_cycle[17162] = 1'b0;  wr_cycle[17162] = 1'b0;  addr_rom[17162]='h00000000;  wr_data_rom[17162]='h00000000;
    rd_cycle[17163] = 1'b0;  wr_cycle[17163] = 1'b0;  addr_rom[17163]='h00000000;  wr_data_rom[17163]='h00000000;
    rd_cycle[17164] = 1'b0;  wr_cycle[17164] = 1'b0;  addr_rom[17164]='h00000000;  wr_data_rom[17164]='h00000000;
    rd_cycle[17165] = 1'b0;  wr_cycle[17165] = 1'b0;  addr_rom[17165]='h00000000;  wr_data_rom[17165]='h00000000;
    rd_cycle[17166] = 1'b0;  wr_cycle[17166] = 1'b0;  addr_rom[17166]='h00000000;  wr_data_rom[17166]='h00000000;
    rd_cycle[17167] = 1'b0;  wr_cycle[17167] = 1'b0;  addr_rom[17167]='h00000000;  wr_data_rom[17167]='h00000000;
    rd_cycle[17168] = 1'b0;  wr_cycle[17168] = 1'b0;  addr_rom[17168]='h00000000;  wr_data_rom[17168]='h00000000;
    rd_cycle[17169] = 1'b0;  wr_cycle[17169] = 1'b0;  addr_rom[17169]='h00000000;  wr_data_rom[17169]='h00000000;
    rd_cycle[17170] = 1'b0;  wr_cycle[17170] = 1'b0;  addr_rom[17170]='h00000000;  wr_data_rom[17170]='h00000000;
    rd_cycle[17171] = 1'b0;  wr_cycle[17171] = 1'b0;  addr_rom[17171]='h00000000;  wr_data_rom[17171]='h00000000;
    rd_cycle[17172] = 1'b0;  wr_cycle[17172] = 1'b0;  addr_rom[17172]='h00000000;  wr_data_rom[17172]='h00000000;
    rd_cycle[17173] = 1'b0;  wr_cycle[17173] = 1'b0;  addr_rom[17173]='h00000000;  wr_data_rom[17173]='h00000000;
    rd_cycle[17174] = 1'b0;  wr_cycle[17174] = 1'b0;  addr_rom[17174]='h00000000;  wr_data_rom[17174]='h00000000;
    rd_cycle[17175] = 1'b0;  wr_cycle[17175] = 1'b0;  addr_rom[17175]='h00000000;  wr_data_rom[17175]='h00000000;
    rd_cycle[17176] = 1'b0;  wr_cycle[17176] = 1'b0;  addr_rom[17176]='h00000000;  wr_data_rom[17176]='h00000000;
    rd_cycle[17177] = 1'b0;  wr_cycle[17177] = 1'b0;  addr_rom[17177]='h00000000;  wr_data_rom[17177]='h00000000;
    rd_cycle[17178] = 1'b0;  wr_cycle[17178] = 1'b0;  addr_rom[17178]='h00000000;  wr_data_rom[17178]='h00000000;
    rd_cycle[17179] = 1'b0;  wr_cycle[17179] = 1'b0;  addr_rom[17179]='h00000000;  wr_data_rom[17179]='h00000000;
    rd_cycle[17180] = 1'b0;  wr_cycle[17180] = 1'b0;  addr_rom[17180]='h00000000;  wr_data_rom[17180]='h00000000;
    rd_cycle[17181] = 1'b0;  wr_cycle[17181] = 1'b0;  addr_rom[17181]='h00000000;  wr_data_rom[17181]='h00000000;
    rd_cycle[17182] = 1'b0;  wr_cycle[17182] = 1'b0;  addr_rom[17182]='h00000000;  wr_data_rom[17182]='h00000000;
    rd_cycle[17183] = 1'b0;  wr_cycle[17183] = 1'b0;  addr_rom[17183]='h00000000;  wr_data_rom[17183]='h00000000;
    rd_cycle[17184] = 1'b0;  wr_cycle[17184] = 1'b0;  addr_rom[17184]='h00000000;  wr_data_rom[17184]='h00000000;
    rd_cycle[17185] = 1'b0;  wr_cycle[17185] = 1'b0;  addr_rom[17185]='h00000000;  wr_data_rom[17185]='h00000000;
    rd_cycle[17186] = 1'b0;  wr_cycle[17186] = 1'b0;  addr_rom[17186]='h00000000;  wr_data_rom[17186]='h00000000;
    rd_cycle[17187] = 1'b0;  wr_cycle[17187] = 1'b0;  addr_rom[17187]='h00000000;  wr_data_rom[17187]='h00000000;
    rd_cycle[17188] = 1'b0;  wr_cycle[17188] = 1'b0;  addr_rom[17188]='h00000000;  wr_data_rom[17188]='h00000000;
    rd_cycle[17189] = 1'b0;  wr_cycle[17189] = 1'b0;  addr_rom[17189]='h00000000;  wr_data_rom[17189]='h00000000;
    rd_cycle[17190] = 1'b0;  wr_cycle[17190] = 1'b0;  addr_rom[17190]='h00000000;  wr_data_rom[17190]='h00000000;
    rd_cycle[17191] = 1'b0;  wr_cycle[17191] = 1'b0;  addr_rom[17191]='h00000000;  wr_data_rom[17191]='h00000000;
    rd_cycle[17192] = 1'b0;  wr_cycle[17192] = 1'b0;  addr_rom[17192]='h00000000;  wr_data_rom[17192]='h00000000;
    rd_cycle[17193] = 1'b0;  wr_cycle[17193] = 1'b0;  addr_rom[17193]='h00000000;  wr_data_rom[17193]='h00000000;
    rd_cycle[17194] = 1'b0;  wr_cycle[17194] = 1'b0;  addr_rom[17194]='h00000000;  wr_data_rom[17194]='h00000000;
    rd_cycle[17195] = 1'b0;  wr_cycle[17195] = 1'b0;  addr_rom[17195]='h00000000;  wr_data_rom[17195]='h00000000;
    rd_cycle[17196] = 1'b0;  wr_cycle[17196] = 1'b0;  addr_rom[17196]='h00000000;  wr_data_rom[17196]='h00000000;
    rd_cycle[17197] = 1'b0;  wr_cycle[17197] = 1'b0;  addr_rom[17197]='h00000000;  wr_data_rom[17197]='h00000000;
    rd_cycle[17198] = 1'b0;  wr_cycle[17198] = 1'b0;  addr_rom[17198]='h00000000;  wr_data_rom[17198]='h00000000;
    rd_cycle[17199] = 1'b0;  wr_cycle[17199] = 1'b0;  addr_rom[17199]='h00000000;  wr_data_rom[17199]='h00000000;
    rd_cycle[17200] = 1'b0;  wr_cycle[17200] = 1'b0;  addr_rom[17200]='h00000000;  wr_data_rom[17200]='h00000000;
    rd_cycle[17201] = 1'b0;  wr_cycle[17201] = 1'b0;  addr_rom[17201]='h00000000;  wr_data_rom[17201]='h00000000;
    rd_cycle[17202] = 1'b0;  wr_cycle[17202] = 1'b0;  addr_rom[17202]='h00000000;  wr_data_rom[17202]='h00000000;
    rd_cycle[17203] = 1'b0;  wr_cycle[17203] = 1'b0;  addr_rom[17203]='h00000000;  wr_data_rom[17203]='h00000000;
    rd_cycle[17204] = 1'b0;  wr_cycle[17204] = 1'b0;  addr_rom[17204]='h00000000;  wr_data_rom[17204]='h00000000;
    rd_cycle[17205] = 1'b0;  wr_cycle[17205] = 1'b0;  addr_rom[17205]='h00000000;  wr_data_rom[17205]='h00000000;
    rd_cycle[17206] = 1'b0;  wr_cycle[17206] = 1'b0;  addr_rom[17206]='h00000000;  wr_data_rom[17206]='h00000000;
    rd_cycle[17207] = 1'b0;  wr_cycle[17207] = 1'b0;  addr_rom[17207]='h00000000;  wr_data_rom[17207]='h00000000;
    rd_cycle[17208] = 1'b0;  wr_cycle[17208] = 1'b0;  addr_rom[17208]='h00000000;  wr_data_rom[17208]='h00000000;
    rd_cycle[17209] = 1'b0;  wr_cycle[17209] = 1'b0;  addr_rom[17209]='h00000000;  wr_data_rom[17209]='h00000000;
    rd_cycle[17210] = 1'b0;  wr_cycle[17210] = 1'b0;  addr_rom[17210]='h00000000;  wr_data_rom[17210]='h00000000;
    rd_cycle[17211] = 1'b0;  wr_cycle[17211] = 1'b0;  addr_rom[17211]='h00000000;  wr_data_rom[17211]='h00000000;
    rd_cycle[17212] = 1'b0;  wr_cycle[17212] = 1'b0;  addr_rom[17212]='h00000000;  wr_data_rom[17212]='h00000000;
    rd_cycle[17213] = 1'b0;  wr_cycle[17213] = 1'b0;  addr_rom[17213]='h00000000;  wr_data_rom[17213]='h00000000;
    rd_cycle[17214] = 1'b0;  wr_cycle[17214] = 1'b0;  addr_rom[17214]='h00000000;  wr_data_rom[17214]='h00000000;
    rd_cycle[17215] = 1'b0;  wr_cycle[17215] = 1'b0;  addr_rom[17215]='h00000000;  wr_data_rom[17215]='h00000000;
    rd_cycle[17216] = 1'b0;  wr_cycle[17216] = 1'b0;  addr_rom[17216]='h00000000;  wr_data_rom[17216]='h00000000;
    rd_cycle[17217] = 1'b0;  wr_cycle[17217] = 1'b0;  addr_rom[17217]='h00000000;  wr_data_rom[17217]='h00000000;
    rd_cycle[17218] = 1'b0;  wr_cycle[17218] = 1'b0;  addr_rom[17218]='h00000000;  wr_data_rom[17218]='h00000000;
    rd_cycle[17219] = 1'b0;  wr_cycle[17219] = 1'b0;  addr_rom[17219]='h00000000;  wr_data_rom[17219]='h00000000;
    rd_cycle[17220] = 1'b0;  wr_cycle[17220] = 1'b0;  addr_rom[17220]='h00000000;  wr_data_rom[17220]='h00000000;
    rd_cycle[17221] = 1'b0;  wr_cycle[17221] = 1'b0;  addr_rom[17221]='h00000000;  wr_data_rom[17221]='h00000000;
    rd_cycle[17222] = 1'b0;  wr_cycle[17222] = 1'b0;  addr_rom[17222]='h00000000;  wr_data_rom[17222]='h00000000;
    rd_cycle[17223] = 1'b0;  wr_cycle[17223] = 1'b0;  addr_rom[17223]='h00000000;  wr_data_rom[17223]='h00000000;
    rd_cycle[17224] = 1'b0;  wr_cycle[17224] = 1'b0;  addr_rom[17224]='h00000000;  wr_data_rom[17224]='h00000000;
    rd_cycle[17225] = 1'b0;  wr_cycle[17225] = 1'b0;  addr_rom[17225]='h00000000;  wr_data_rom[17225]='h00000000;
    rd_cycle[17226] = 1'b0;  wr_cycle[17226] = 1'b0;  addr_rom[17226]='h00000000;  wr_data_rom[17226]='h00000000;
    rd_cycle[17227] = 1'b0;  wr_cycle[17227] = 1'b0;  addr_rom[17227]='h00000000;  wr_data_rom[17227]='h00000000;
    rd_cycle[17228] = 1'b0;  wr_cycle[17228] = 1'b0;  addr_rom[17228]='h00000000;  wr_data_rom[17228]='h00000000;
    rd_cycle[17229] = 1'b0;  wr_cycle[17229] = 1'b0;  addr_rom[17229]='h00000000;  wr_data_rom[17229]='h00000000;
    rd_cycle[17230] = 1'b0;  wr_cycle[17230] = 1'b0;  addr_rom[17230]='h00000000;  wr_data_rom[17230]='h00000000;
    rd_cycle[17231] = 1'b0;  wr_cycle[17231] = 1'b0;  addr_rom[17231]='h00000000;  wr_data_rom[17231]='h00000000;
    rd_cycle[17232] = 1'b0;  wr_cycle[17232] = 1'b0;  addr_rom[17232]='h00000000;  wr_data_rom[17232]='h00000000;
    rd_cycle[17233] = 1'b0;  wr_cycle[17233] = 1'b0;  addr_rom[17233]='h00000000;  wr_data_rom[17233]='h00000000;
    rd_cycle[17234] = 1'b0;  wr_cycle[17234] = 1'b0;  addr_rom[17234]='h00000000;  wr_data_rom[17234]='h00000000;
    rd_cycle[17235] = 1'b0;  wr_cycle[17235] = 1'b0;  addr_rom[17235]='h00000000;  wr_data_rom[17235]='h00000000;
    rd_cycle[17236] = 1'b0;  wr_cycle[17236] = 1'b0;  addr_rom[17236]='h00000000;  wr_data_rom[17236]='h00000000;
    rd_cycle[17237] = 1'b0;  wr_cycle[17237] = 1'b0;  addr_rom[17237]='h00000000;  wr_data_rom[17237]='h00000000;
    rd_cycle[17238] = 1'b0;  wr_cycle[17238] = 1'b0;  addr_rom[17238]='h00000000;  wr_data_rom[17238]='h00000000;
    rd_cycle[17239] = 1'b0;  wr_cycle[17239] = 1'b0;  addr_rom[17239]='h00000000;  wr_data_rom[17239]='h00000000;
    rd_cycle[17240] = 1'b0;  wr_cycle[17240] = 1'b0;  addr_rom[17240]='h00000000;  wr_data_rom[17240]='h00000000;
    rd_cycle[17241] = 1'b0;  wr_cycle[17241] = 1'b0;  addr_rom[17241]='h00000000;  wr_data_rom[17241]='h00000000;
    rd_cycle[17242] = 1'b0;  wr_cycle[17242] = 1'b0;  addr_rom[17242]='h00000000;  wr_data_rom[17242]='h00000000;
    rd_cycle[17243] = 1'b0;  wr_cycle[17243] = 1'b0;  addr_rom[17243]='h00000000;  wr_data_rom[17243]='h00000000;
    rd_cycle[17244] = 1'b0;  wr_cycle[17244] = 1'b0;  addr_rom[17244]='h00000000;  wr_data_rom[17244]='h00000000;
    rd_cycle[17245] = 1'b0;  wr_cycle[17245] = 1'b0;  addr_rom[17245]='h00000000;  wr_data_rom[17245]='h00000000;
    rd_cycle[17246] = 1'b0;  wr_cycle[17246] = 1'b0;  addr_rom[17246]='h00000000;  wr_data_rom[17246]='h00000000;
    rd_cycle[17247] = 1'b0;  wr_cycle[17247] = 1'b0;  addr_rom[17247]='h00000000;  wr_data_rom[17247]='h00000000;
    rd_cycle[17248] = 1'b0;  wr_cycle[17248] = 1'b0;  addr_rom[17248]='h00000000;  wr_data_rom[17248]='h00000000;
    rd_cycle[17249] = 1'b0;  wr_cycle[17249] = 1'b0;  addr_rom[17249]='h00000000;  wr_data_rom[17249]='h00000000;
    rd_cycle[17250] = 1'b0;  wr_cycle[17250] = 1'b0;  addr_rom[17250]='h00000000;  wr_data_rom[17250]='h00000000;
    rd_cycle[17251] = 1'b0;  wr_cycle[17251] = 1'b0;  addr_rom[17251]='h00000000;  wr_data_rom[17251]='h00000000;
    rd_cycle[17252] = 1'b0;  wr_cycle[17252] = 1'b0;  addr_rom[17252]='h00000000;  wr_data_rom[17252]='h00000000;
    rd_cycle[17253] = 1'b0;  wr_cycle[17253] = 1'b0;  addr_rom[17253]='h00000000;  wr_data_rom[17253]='h00000000;
    rd_cycle[17254] = 1'b0;  wr_cycle[17254] = 1'b0;  addr_rom[17254]='h00000000;  wr_data_rom[17254]='h00000000;
    rd_cycle[17255] = 1'b0;  wr_cycle[17255] = 1'b0;  addr_rom[17255]='h00000000;  wr_data_rom[17255]='h00000000;
    rd_cycle[17256] = 1'b0;  wr_cycle[17256] = 1'b0;  addr_rom[17256]='h00000000;  wr_data_rom[17256]='h00000000;
    rd_cycle[17257] = 1'b0;  wr_cycle[17257] = 1'b0;  addr_rom[17257]='h00000000;  wr_data_rom[17257]='h00000000;
    rd_cycle[17258] = 1'b0;  wr_cycle[17258] = 1'b0;  addr_rom[17258]='h00000000;  wr_data_rom[17258]='h00000000;
    rd_cycle[17259] = 1'b0;  wr_cycle[17259] = 1'b0;  addr_rom[17259]='h00000000;  wr_data_rom[17259]='h00000000;
    rd_cycle[17260] = 1'b0;  wr_cycle[17260] = 1'b0;  addr_rom[17260]='h00000000;  wr_data_rom[17260]='h00000000;
    rd_cycle[17261] = 1'b0;  wr_cycle[17261] = 1'b0;  addr_rom[17261]='h00000000;  wr_data_rom[17261]='h00000000;
    rd_cycle[17262] = 1'b0;  wr_cycle[17262] = 1'b0;  addr_rom[17262]='h00000000;  wr_data_rom[17262]='h00000000;
    rd_cycle[17263] = 1'b0;  wr_cycle[17263] = 1'b0;  addr_rom[17263]='h00000000;  wr_data_rom[17263]='h00000000;
    rd_cycle[17264] = 1'b0;  wr_cycle[17264] = 1'b0;  addr_rom[17264]='h00000000;  wr_data_rom[17264]='h00000000;
    rd_cycle[17265] = 1'b0;  wr_cycle[17265] = 1'b0;  addr_rom[17265]='h00000000;  wr_data_rom[17265]='h00000000;
    rd_cycle[17266] = 1'b0;  wr_cycle[17266] = 1'b0;  addr_rom[17266]='h00000000;  wr_data_rom[17266]='h00000000;
    rd_cycle[17267] = 1'b0;  wr_cycle[17267] = 1'b0;  addr_rom[17267]='h00000000;  wr_data_rom[17267]='h00000000;
    rd_cycle[17268] = 1'b0;  wr_cycle[17268] = 1'b0;  addr_rom[17268]='h00000000;  wr_data_rom[17268]='h00000000;
    rd_cycle[17269] = 1'b0;  wr_cycle[17269] = 1'b0;  addr_rom[17269]='h00000000;  wr_data_rom[17269]='h00000000;
    rd_cycle[17270] = 1'b0;  wr_cycle[17270] = 1'b0;  addr_rom[17270]='h00000000;  wr_data_rom[17270]='h00000000;
    rd_cycle[17271] = 1'b0;  wr_cycle[17271] = 1'b0;  addr_rom[17271]='h00000000;  wr_data_rom[17271]='h00000000;
    rd_cycle[17272] = 1'b0;  wr_cycle[17272] = 1'b0;  addr_rom[17272]='h00000000;  wr_data_rom[17272]='h00000000;
    rd_cycle[17273] = 1'b0;  wr_cycle[17273] = 1'b0;  addr_rom[17273]='h00000000;  wr_data_rom[17273]='h00000000;
    rd_cycle[17274] = 1'b0;  wr_cycle[17274] = 1'b0;  addr_rom[17274]='h00000000;  wr_data_rom[17274]='h00000000;
    rd_cycle[17275] = 1'b0;  wr_cycle[17275] = 1'b0;  addr_rom[17275]='h00000000;  wr_data_rom[17275]='h00000000;
    rd_cycle[17276] = 1'b0;  wr_cycle[17276] = 1'b0;  addr_rom[17276]='h00000000;  wr_data_rom[17276]='h00000000;
    rd_cycle[17277] = 1'b0;  wr_cycle[17277] = 1'b0;  addr_rom[17277]='h00000000;  wr_data_rom[17277]='h00000000;
    rd_cycle[17278] = 1'b0;  wr_cycle[17278] = 1'b0;  addr_rom[17278]='h00000000;  wr_data_rom[17278]='h00000000;
    rd_cycle[17279] = 1'b0;  wr_cycle[17279] = 1'b0;  addr_rom[17279]='h00000000;  wr_data_rom[17279]='h00000000;
    rd_cycle[17280] = 1'b0;  wr_cycle[17280] = 1'b0;  addr_rom[17280]='h00000000;  wr_data_rom[17280]='h00000000;
    rd_cycle[17281] = 1'b0;  wr_cycle[17281] = 1'b0;  addr_rom[17281]='h00000000;  wr_data_rom[17281]='h00000000;
    rd_cycle[17282] = 1'b0;  wr_cycle[17282] = 1'b0;  addr_rom[17282]='h00000000;  wr_data_rom[17282]='h00000000;
    rd_cycle[17283] = 1'b0;  wr_cycle[17283] = 1'b0;  addr_rom[17283]='h00000000;  wr_data_rom[17283]='h00000000;
    rd_cycle[17284] = 1'b0;  wr_cycle[17284] = 1'b0;  addr_rom[17284]='h00000000;  wr_data_rom[17284]='h00000000;
    rd_cycle[17285] = 1'b0;  wr_cycle[17285] = 1'b0;  addr_rom[17285]='h00000000;  wr_data_rom[17285]='h00000000;
    rd_cycle[17286] = 1'b0;  wr_cycle[17286] = 1'b0;  addr_rom[17286]='h00000000;  wr_data_rom[17286]='h00000000;
    rd_cycle[17287] = 1'b0;  wr_cycle[17287] = 1'b0;  addr_rom[17287]='h00000000;  wr_data_rom[17287]='h00000000;
    rd_cycle[17288] = 1'b0;  wr_cycle[17288] = 1'b0;  addr_rom[17288]='h00000000;  wr_data_rom[17288]='h00000000;
    rd_cycle[17289] = 1'b0;  wr_cycle[17289] = 1'b0;  addr_rom[17289]='h00000000;  wr_data_rom[17289]='h00000000;
    rd_cycle[17290] = 1'b0;  wr_cycle[17290] = 1'b0;  addr_rom[17290]='h00000000;  wr_data_rom[17290]='h00000000;
    rd_cycle[17291] = 1'b0;  wr_cycle[17291] = 1'b0;  addr_rom[17291]='h00000000;  wr_data_rom[17291]='h00000000;
    rd_cycle[17292] = 1'b0;  wr_cycle[17292] = 1'b0;  addr_rom[17292]='h00000000;  wr_data_rom[17292]='h00000000;
    rd_cycle[17293] = 1'b0;  wr_cycle[17293] = 1'b0;  addr_rom[17293]='h00000000;  wr_data_rom[17293]='h00000000;
    rd_cycle[17294] = 1'b0;  wr_cycle[17294] = 1'b0;  addr_rom[17294]='h00000000;  wr_data_rom[17294]='h00000000;
    rd_cycle[17295] = 1'b0;  wr_cycle[17295] = 1'b0;  addr_rom[17295]='h00000000;  wr_data_rom[17295]='h00000000;
    rd_cycle[17296] = 1'b0;  wr_cycle[17296] = 1'b0;  addr_rom[17296]='h00000000;  wr_data_rom[17296]='h00000000;
    rd_cycle[17297] = 1'b0;  wr_cycle[17297] = 1'b0;  addr_rom[17297]='h00000000;  wr_data_rom[17297]='h00000000;
    rd_cycle[17298] = 1'b0;  wr_cycle[17298] = 1'b0;  addr_rom[17298]='h00000000;  wr_data_rom[17298]='h00000000;
    rd_cycle[17299] = 1'b0;  wr_cycle[17299] = 1'b0;  addr_rom[17299]='h00000000;  wr_data_rom[17299]='h00000000;
    rd_cycle[17300] = 1'b0;  wr_cycle[17300] = 1'b0;  addr_rom[17300]='h00000000;  wr_data_rom[17300]='h00000000;
    rd_cycle[17301] = 1'b0;  wr_cycle[17301] = 1'b0;  addr_rom[17301]='h00000000;  wr_data_rom[17301]='h00000000;
    rd_cycle[17302] = 1'b0;  wr_cycle[17302] = 1'b0;  addr_rom[17302]='h00000000;  wr_data_rom[17302]='h00000000;
    rd_cycle[17303] = 1'b0;  wr_cycle[17303] = 1'b0;  addr_rom[17303]='h00000000;  wr_data_rom[17303]='h00000000;
    rd_cycle[17304] = 1'b0;  wr_cycle[17304] = 1'b0;  addr_rom[17304]='h00000000;  wr_data_rom[17304]='h00000000;
    rd_cycle[17305] = 1'b0;  wr_cycle[17305] = 1'b0;  addr_rom[17305]='h00000000;  wr_data_rom[17305]='h00000000;
    rd_cycle[17306] = 1'b0;  wr_cycle[17306] = 1'b0;  addr_rom[17306]='h00000000;  wr_data_rom[17306]='h00000000;
    rd_cycle[17307] = 1'b0;  wr_cycle[17307] = 1'b0;  addr_rom[17307]='h00000000;  wr_data_rom[17307]='h00000000;
    rd_cycle[17308] = 1'b0;  wr_cycle[17308] = 1'b0;  addr_rom[17308]='h00000000;  wr_data_rom[17308]='h00000000;
    rd_cycle[17309] = 1'b0;  wr_cycle[17309] = 1'b0;  addr_rom[17309]='h00000000;  wr_data_rom[17309]='h00000000;
    rd_cycle[17310] = 1'b0;  wr_cycle[17310] = 1'b0;  addr_rom[17310]='h00000000;  wr_data_rom[17310]='h00000000;
    rd_cycle[17311] = 1'b0;  wr_cycle[17311] = 1'b0;  addr_rom[17311]='h00000000;  wr_data_rom[17311]='h00000000;
    rd_cycle[17312] = 1'b0;  wr_cycle[17312] = 1'b0;  addr_rom[17312]='h00000000;  wr_data_rom[17312]='h00000000;
    rd_cycle[17313] = 1'b0;  wr_cycle[17313] = 1'b0;  addr_rom[17313]='h00000000;  wr_data_rom[17313]='h00000000;
    rd_cycle[17314] = 1'b0;  wr_cycle[17314] = 1'b0;  addr_rom[17314]='h00000000;  wr_data_rom[17314]='h00000000;
    rd_cycle[17315] = 1'b0;  wr_cycle[17315] = 1'b0;  addr_rom[17315]='h00000000;  wr_data_rom[17315]='h00000000;
    rd_cycle[17316] = 1'b0;  wr_cycle[17316] = 1'b0;  addr_rom[17316]='h00000000;  wr_data_rom[17316]='h00000000;
    rd_cycle[17317] = 1'b0;  wr_cycle[17317] = 1'b0;  addr_rom[17317]='h00000000;  wr_data_rom[17317]='h00000000;
    rd_cycle[17318] = 1'b0;  wr_cycle[17318] = 1'b0;  addr_rom[17318]='h00000000;  wr_data_rom[17318]='h00000000;
    rd_cycle[17319] = 1'b0;  wr_cycle[17319] = 1'b0;  addr_rom[17319]='h00000000;  wr_data_rom[17319]='h00000000;
    rd_cycle[17320] = 1'b0;  wr_cycle[17320] = 1'b0;  addr_rom[17320]='h00000000;  wr_data_rom[17320]='h00000000;
    rd_cycle[17321] = 1'b0;  wr_cycle[17321] = 1'b0;  addr_rom[17321]='h00000000;  wr_data_rom[17321]='h00000000;
    rd_cycle[17322] = 1'b0;  wr_cycle[17322] = 1'b0;  addr_rom[17322]='h00000000;  wr_data_rom[17322]='h00000000;
    rd_cycle[17323] = 1'b0;  wr_cycle[17323] = 1'b0;  addr_rom[17323]='h00000000;  wr_data_rom[17323]='h00000000;
    rd_cycle[17324] = 1'b0;  wr_cycle[17324] = 1'b0;  addr_rom[17324]='h00000000;  wr_data_rom[17324]='h00000000;
    rd_cycle[17325] = 1'b0;  wr_cycle[17325] = 1'b0;  addr_rom[17325]='h00000000;  wr_data_rom[17325]='h00000000;
    rd_cycle[17326] = 1'b0;  wr_cycle[17326] = 1'b0;  addr_rom[17326]='h00000000;  wr_data_rom[17326]='h00000000;
    rd_cycle[17327] = 1'b0;  wr_cycle[17327] = 1'b0;  addr_rom[17327]='h00000000;  wr_data_rom[17327]='h00000000;
    rd_cycle[17328] = 1'b0;  wr_cycle[17328] = 1'b0;  addr_rom[17328]='h00000000;  wr_data_rom[17328]='h00000000;
    rd_cycle[17329] = 1'b0;  wr_cycle[17329] = 1'b0;  addr_rom[17329]='h00000000;  wr_data_rom[17329]='h00000000;
    rd_cycle[17330] = 1'b0;  wr_cycle[17330] = 1'b0;  addr_rom[17330]='h00000000;  wr_data_rom[17330]='h00000000;
    rd_cycle[17331] = 1'b0;  wr_cycle[17331] = 1'b0;  addr_rom[17331]='h00000000;  wr_data_rom[17331]='h00000000;
    rd_cycle[17332] = 1'b0;  wr_cycle[17332] = 1'b0;  addr_rom[17332]='h00000000;  wr_data_rom[17332]='h00000000;
    rd_cycle[17333] = 1'b0;  wr_cycle[17333] = 1'b0;  addr_rom[17333]='h00000000;  wr_data_rom[17333]='h00000000;
    rd_cycle[17334] = 1'b0;  wr_cycle[17334] = 1'b0;  addr_rom[17334]='h00000000;  wr_data_rom[17334]='h00000000;
    rd_cycle[17335] = 1'b0;  wr_cycle[17335] = 1'b0;  addr_rom[17335]='h00000000;  wr_data_rom[17335]='h00000000;
    rd_cycle[17336] = 1'b0;  wr_cycle[17336] = 1'b0;  addr_rom[17336]='h00000000;  wr_data_rom[17336]='h00000000;
    rd_cycle[17337] = 1'b0;  wr_cycle[17337] = 1'b0;  addr_rom[17337]='h00000000;  wr_data_rom[17337]='h00000000;
    rd_cycle[17338] = 1'b0;  wr_cycle[17338] = 1'b0;  addr_rom[17338]='h00000000;  wr_data_rom[17338]='h00000000;
    rd_cycle[17339] = 1'b0;  wr_cycle[17339] = 1'b0;  addr_rom[17339]='h00000000;  wr_data_rom[17339]='h00000000;
    rd_cycle[17340] = 1'b0;  wr_cycle[17340] = 1'b0;  addr_rom[17340]='h00000000;  wr_data_rom[17340]='h00000000;
    rd_cycle[17341] = 1'b0;  wr_cycle[17341] = 1'b0;  addr_rom[17341]='h00000000;  wr_data_rom[17341]='h00000000;
    rd_cycle[17342] = 1'b0;  wr_cycle[17342] = 1'b0;  addr_rom[17342]='h00000000;  wr_data_rom[17342]='h00000000;
    rd_cycle[17343] = 1'b0;  wr_cycle[17343] = 1'b0;  addr_rom[17343]='h00000000;  wr_data_rom[17343]='h00000000;
    rd_cycle[17344] = 1'b0;  wr_cycle[17344] = 1'b0;  addr_rom[17344]='h00000000;  wr_data_rom[17344]='h00000000;
    rd_cycle[17345] = 1'b0;  wr_cycle[17345] = 1'b0;  addr_rom[17345]='h00000000;  wr_data_rom[17345]='h00000000;
    rd_cycle[17346] = 1'b0;  wr_cycle[17346] = 1'b0;  addr_rom[17346]='h00000000;  wr_data_rom[17346]='h00000000;
    rd_cycle[17347] = 1'b0;  wr_cycle[17347] = 1'b0;  addr_rom[17347]='h00000000;  wr_data_rom[17347]='h00000000;
    rd_cycle[17348] = 1'b0;  wr_cycle[17348] = 1'b0;  addr_rom[17348]='h00000000;  wr_data_rom[17348]='h00000000;
    rd_cycle[17349] = 1'b0;  wr_cycle[17349] = 1'b0;  addr_rom[17349]='h00000000;  wr_data_rom[17349]='h00000000;
    rd_cycle[17350] = 1'b0;  wr_cycle[17350] = 1'b0;  addr_rom[17350]='h00000000;  wr_data_rom[17350]='h00000000;
    rd_cycle[17351] = 1'b0;  wr_cycle[17351] = 1'b0;  addr_rom[17351]='h00000000;  wr_data_rom[17351]='h00000000;
    rd_cycle[17352] = 1'b0;  wr_cycle[17352] = 1'b0;  addr_rom[17352]='h00000000;  wr_data_rom[17352]='h00000000;
    rd_cycle[17353] = 1'b0;  wr_cycle[17353] = 1'b0;  addr_rom[17353]='h00000000;  wr_data_rom[17353]='h00000000;
    rd_cycle[17354] = 1'b0;  wr_cycle[17354] = 1'b0;  addr_rom[17354]='h00000000;  wr_data_rom[17354]='h00000000;
    rd_cycle[17355] = 1'b0;  wr_cycle[17355] = 1'b0;  addr_rom[17355]='h00000000;  wr_data_rom[17355]='h00000000;
    rd_cycle[17356] = 1'b0;  wr_cycle[17356] = 1'b0;  addr_rom[17356]='h00000000;  wr_data_rom[17356]='h00000000;
    rd_cycle[17357] = 1'b0;  wr_cycle[17357] = 1'b0;  addr_rom[17357]='h00000000;  wr_data_rom[17357]='h00000000;
    rd_cycle[17358] = 1'b0;  wr_cycle[17358] = 1'b0;  addr_rom[17358]='h00000000;  wr_data_rom[17358]='h00000000;
    rd_cycle[17359] = 1'b0;  wr_cycle[17359] = 1'b0;  addr_rom[17359]='h00000000;  wr_data_rom[17359]='h00000000;
    rd_cycle[17360] = 1'b0;  wr_cycle[17360] = 1'b0;  addr_rom[17360]='h00000000;  wr_data_rom[17360]='h00000000;
    rd_cycle[17361] = 1'b0;  wr_cycle[17361] = 1'b0;  addr_rom[17361]='h00000000;  wr_data_rom[17361]='h00000000;
    rd_cycle[17362] = 1'b0;  wr_cycle[17362] = 1'b0;  addr_rom[17362]='h00000000;  wr_data_rom[17362]='h00000000;
    rd_cycle[17363] = 1'b0;  wr_cycle[17363] = 1'b0;  addr_rom[17363]='h00000000;  wr_data_rom[17363]='h00000000;
    rd_cycle[17364] = 1'b0;  wr_cycle[17364] = 1'b0;  addr_rom[17364]='h00000000;  wr_data_rom[17364]='h00000000;
    rd_cycle[17365] = 1'b0;  wr_cycle[17365] = 1'b0;  addr_rom[17365]='h00000000;  wr_data_rom[17365]='h00000000;
    rd_cycle[17366] = 1'b0;  wr_cycle[17366] = 1'b0;  addr_rom[17366]='h00000000;  wr_data_rom[17366]='h00000000;
    rd_cycle[17367] = 1'b0;  wr_cycle[17367] = 1'b0;  addr_rom[17367]='h00000000;  wr_data_rom[17367]='h00000000;
    rd_cycle[17368] = 1'b0;  wr_cycle[17368] = 1'b0;  addr_rom[17368]='h00000000;  wr_data_rom[17368]='h00000000;
    rd_cycle[17369] = 1'b0;  wr_cycle[17369] = 1'b0;  addr_rom[17369]='h00000000;  wr_data_rom[17369]='h00000000;
    rd_cycle[17370] = 1'b0;  wr_cycle[17370] = 1'b0;  addr_rom[17370]='h00000000;  wr_data_rom[17370]='h00000000;
    rd_cycle[17371] = 1'b0;  wr_cycle[17371] = 1'b0;  addr_rom[17371]='h00000000;  wr_data_rom[17371]='h00000000;
    rd_cycle[17372] = 1'b0;  wr_cycle[17372] = 1'b0;  addr_rom[17372]='h00000000;  wr_data_rom[17372]='h00000000;
    rd_cycle[17373] = 1'b0;  wr_cycle[17373] = 1'b0;  addr_rom[17373]='h00000000;  wr_data_rom[17373]='h00000000;
    rd_cycle[17374] = 1'b0;  wr_cycle[17374] = 1'b0;  addr_rom[17374]='h00000000;  wr_data_rom[17374]='h00000000;
    rd_cycle[17375] = 1'b0;  wr_cycle[17375] = 1'b0;  addr_rom[17375]='h00000000;  wr_data_rom[17375]='h00000000;
    rd_cycle[17376] = 1'b0;  wr_cycle[17376] = 1'b0;  addr_rom[17376]='h00000000;  wr_data_rom[17376]='h00000000;
    rd_cycle[17377] = 1'b0;  wr_cycle[17377] = 1'b0;  addr_rom[17377]='h00000000;  wr_data_rom[17377]='h00000000;
    rd_cycle[17378] = 1'b0;  wr_cycle[17378] = 1'b0;  addr_rom[17378]='h00000000;  wr_data_rom[17378]='h00000000;
    rd_cycle[17379] = 1'b0;  wr_cycle[17379] = 1'b0;  addr_rom[17379]='h00000000;  wr_data_rom[17379]='h00000000;
    rd_cycle[17380] = 1'b0;  wr_cycle[17380] = 1'b0;  addr_rom[17380]='h00000000;  wr_data_rom[17380]='h00000000;
    rd_cycle[17381] = 1'b0;  wr_cycle[17381] = 1'b0;  addr_rom[17381]='h00000000;  wr_data_rom[17381]='h00000000;
    rd_cycle[17382] = 1'b0;  wr_cycle[17382] = 1'b0;  addr_rom[17382]='h00000000;  wr_data_rom[17382]='h00000000;
    rd_cycle[17383] = 1'b0;  wr_cycle[17383] = 1'b0;  addr_rom[17383]='h00000000;  wr_data_rom[17383]='h00000000;
    rd_cycle[17384] = 1'b0;  wr_cycle[17384] = 1'b0;  addr_rom[17384]='h00000000;  wr_data_rom[17384]='h00000000;
    rd_cycle[17385] = 1'b0;  wr_cycle[17385] = 1'b0;  addr_rom[17385]='h00000000;  wr_data_rom[17385]='h00000000;
    rd_cycle[17386] = 1'b0;  wr_cycle[17386] = 1'b0;  addr_rom[17386]='h00000000;  wr_data_rom[17386]='h00000000;
    rd_cycle[17387] = 1'b0;  wr_cycle[17387] = 1'b0;  addr_rom[17387]='h00000000;  wr_data_rom[17387]='h00000000;
    rd_cycle[17388] = 1'b0;  wr_cycle[17388] = 1'b0;  addr_rom[17388]='h00000000;  wr_data_rom[17388]='h00000000;
    rd_cycle[17389] = 1'b0;  wr_cycle[17389] = 1'b0;  addr_rom[17389]='h00000000;  wr_data_rom[17389]='h00000000;
    rd_cycle[17390] = 1'b0;  wr_cycle[17390] = 1'b0;  addr_rom[17390]='h00000000;  wr_data_rom[17390]='h00000000;
    rd_cycle[17391] = 1'b0;  wr_cycle[17391] = 1'b0;  addr_rom[17391]='h00000000;  wr_data_rom[17391]='h00000000;
    rd_cycle[17392] = 1'b0;  wr_cycle[17392] = 1'b0;  addr_rom[17392]='h00000000;  wr_data_rom[17392]='h00000000;
    rd_cycle[17393] = 1'b0;  wr_cycle[17393] = 1'b0;  addr_rom[17393]='h00000000;  wr_data_rom[17393]='h00000000;
    rd_cycle[17394] = 1'b0;  wr_cycle[17394] = 1'b0;  addr_rom[17394]='h00000000;  wr_data_rom[17394]='h00000000;
    rd_cycle[17395] = 1'b0;  wr_cycle[17395] = 1'b0;  addr_rom[17395]='h00000000;  wr_data_rom[17395]='h00000000;
    rd_cycle[17396] = 1'b0;  wr_cycle[17396] = 1'b0;  addr_rom[17396]='h00000000;  wr_data_rom[17396]='h00000000;
    rd_cycle[17397] = 1'b0;  wr_cycle[17397] = 1'b0;  addr_rom[17397]='h00000000;  wr_data_rom[17397]='h00000000;
    rd_cycle[17398] = 1'b0;  wr_cycle[17398] = 1'b0;  addr_rom[17398]='h00000000;  wr_data_rom[17398]='h00000000;
    rd_cycle[17399] = 1'b0;  wr_cycle[17399] = 1'b0;  addr_rom[17399]='h00000000;  wr_data_rom[17399]='h00000000;
    rd_cycle[17400] = 1'b0;  wr_cycle[17400] = 1'b0;  addr_rom[17400]='h00000000;  wr_data_rom[17400]='h00000000;
    rd_cycle[17401] = 1'b0;  wr_cycle[17401] = 1'b0;  addr_rom[17401]='h00000000;  wr_data_rom[17401]='h00000000;
    rd_cycle[17402] = 1'b0;  wr_cycle[17402] = 1'b0;  addr_rom[17402]='h00000000;  wr_data_rom[17402]='h00000000;
    rd_cycle[17403] = 1'b0;  wr_cycle[17403] = 1'b0;  addr_rom[17403]='h00000000;  wr_data_rom[17403]='h00000000;
    rd_cycle[17404] = 1'b0;  wr_cycle[17404] = 1'b0;  addr_rom[17404]='h00000000;  wr_data_rom[17404]='h00000000;
    rd_cycle[17405] = 1'b0;  wr_cycle[17405] = 1'b0;  addr_rom[17405]='h00000000;  wr_data_rom[17405]='h00000000;
    rd_cycle[17406] = 1'b0;  wr_cycle[17406] = 1'b0;  addr_rom[17406]='h00000000;  wr_data_rom[17406]='h00000000;
    rd_cycle[17407] = 1'b0;  wr_cycle[17407] = 1'b0;  addr_rom[17407]='h00000000;  wr_data_rom[17407]='h00000000;
    rd_cycle[17408] = 1'b0;  wr_cycle[17408] = 1'b0;  addr_rom[17408]='h00000000;  wr_data_rom[17408]='h00000000;
    rd_cycle[17409] = 1'b0;  wr_cycle[17409] = 1'b0;  addr_rom[17409]='h00000000;  wr_data_rom[17409]='h00000000;
    rd_cycle[17410] = 1'b0;  wr_cycle[17410] = 1'b0;  addr_rom[17410]='h00000000;  wr_data_rom[17410]='h00000000;
    rd_cycle[17411] = 1'b0;  wr_cycle[17411] = 1'b0;  addr_rom[17411]='h00000000;  wr_data_rom[17411]='h00000000;
    rd_cycle[17412] = 1'b0;  wr_cycle[17412] = 1'b0;  addr_rom[17412]='h00000000;  wr_data_rom[17412]='h00000000;
    rd_cycle[17413] = 1'b0;  wr_cycle[17413] = 1'b0;  addr_rom[17413]='h00000000;  wr_data_rom[17413]='h00000000;
    rd_cycle[17414] = 1'b0;  wr_cycle[17414] = 1'b0;  addr_rom[17414]='h00000000;  wr_data_rom[17414]='h00000000;
    rd_cycle[17415] = 1'b0;  wr_cycle[17415] = 1'b0;  addr_rom[17415]='h00000000;  wr_data_rom[17415]='h00000000;
    rd_cycle[17416] = 1'b0;  wr_cycle[17416] = 1'b0;  addr_rom[17416]='h00000000;  wr_data_rom[17416]='h00000000;
    rd_cycle[17417] = 1'b0;  wr_cycle[17417] = 1'b0;  addr_rom[17417]='h00000000;  wr_data_rom[17417]='h00000000;
    rd_cycle[17418] = 1'b0;  wr_cycle[17418] = 1'b0;  addr_rom[17418]='h00000000;  wr_data_rom[17418]='h00000000;
    rd_cycle[17419] = 1'b0;  wr_cycle[17419] = 1'b0;  addr_rom[17419]='h00000000;  wr_data_rom[17419]='h00000000;
    rd_cycle[17420] = 1'b0;  wr_cycle[17420] = 1'b0;  addr_rom[17420]='h00000000;  wr_data_rom[17420]='h00000000;
    rd_cycle[17421] = 1'b0;  wr_cycle[17421] = 1'b0;  addr_rom[17421]='h00000000;  wr_data_rom[17421]='h00000000;
    rd_cycle[17422] = 1'b0;  wr_cycle[17422] = 1'b0;  addr_rom[17422]='h00000000;  wr_data_rom[17422]='h00000000;
    rd_cycle[17423] = 1'b0;  wr_cycle[17423] = 1'b0;  addr_rom[17423]='h00000000;  wr_data_rom[17423]='h00000000;
    rd_cycle[17424] = 1'b0;  wr_cycle[17424] = 1'b0;  addr_rom[17424]='h00000000;  wr_data_rom[17424]='h00000000;
    rd_cycle[17425] = 1'b0;  wr_cycle[17425] = 1'b0;  addr_rom[17425]='h00000000;  wr_data_rom[17425]='h00000000;
    rd_cycle[17426] = 1'b0;  wr_cycle[17426] = 1'b0;  addr_rom[17426]='h00000000;  wr_data_rom[17426]='h00000000;
    rd_cycle[17427] = 1'b0;  wr_cycle[17427] = 1'b0;  addr_rom[17427]='h00000000;  wr_data_rom[17427]='h00000000;
    rd_cycle[17428] = 1'b0;  wr_cycle[17428] = 1'b0;  addr_rom[17428]='h00000000;  wr_data_rom[17428]='h00000000;
    rd_cycle[17429] = 1'b0;  wr_cycle[17429] = 1'b0;  addr_rom[17429]='h00000000;  wr_data_rom[17429]='h00000000;
    rd_cycle[17430] = 1'b0;  wr_cycle[17430] = 1'b0;  addr_rom[17430]='h00000000;  wr_data_rom[17430]='h00000000;
    rd_cycle[17431] = 1'b0;  wr_cycle[17431] = 1'b0;  addr_rom[17431]='h00000000;  wr_data_rom[17431]='h00000000;
    rd_cycle[17432] = 1'b0;  wr_cycle[17432] = 1'b0;  addr_rom[17432]='h00000000;  wr_data_rom[17432]='h00000000;
    rd_cycle[17433] = 1'b0;  wr_cycle[17433] = 1'b0;  addr_rom[17433]='h00000000;  wr_data_rom[17433]='h00000000;
    rd_cycle[17434] = 1'b0;  wr_cycle[17434] = 1'b0;  addr_rom[17434]='h00000000;  wr_data_rom[17434]='h00000000;
    rd_cycle[17435] = 1'b0;  wr_cycle[17435] = 1'b0;  addr_rom[17435]='h00000000;  wr_data_rom[17435]='h00000000;
    rd_cycle[17436] = 1'b0;  wr_cycle[17436] = 1'b0;  addr_rom[17436]='h00000000;  wr_data_rom[17436]='h00000000;
    rd_cycle[17437] = 1'b0;  wr_cycle[17437] = 1'b0;  addr_rom[17437]='h00000000;  wr_data_rom[17437]='h00000000;
    rd_cycle[17438] = 1'b0;  wr_cycle[17438] = 1'b0;  addr_rom[17438]='h00000000;  wr_data_rom[17438]='h00000000;
    rd_cycle[17439] = 1'b0;  wr_cycle[17439] = 1'b0;  addr_rom[17439]='h00000000;  wr_data_rom[17439]='h00000000;
    rd_cycle[17440] = 1'b0;  wr_cycle[17440] = 1'b0;  addr_rom[17440]='h00000000;  wr_data_rom[17440]='h00000000;
    rd_cycle[17441] = 1'b0;  wr_cycle[17441] = 1'b0;  addr_rom[17441]='h00000000;  wr_data_rom[17441]='h00000000;
    rd_cycle[17442] = 1'b0;  wr_cycle[17442] = 1'b0;  addr_rom[17442]='h00000000;  wr_data_rom[17442]='h00000000;
    rd_cycle[17443] = 1'b0;  wr_cycle[17443] = 1'b0;  addr_rom[17443]='h00000000;  wr_data_rom[17443]='h00000000;
    rd_cycle[17444] = 1'b0;  wr_cycle[17444] = 1'b0;  addr_rom[17444]='h00000000;  wr_data_rom[17444]='h00000000;
    rd_cycle[17445] = 1'b0;  wr_cycle[17445] = 1'b0;  addr_rom[17445]='h00000000;  wr_data_rom[17445]='h00000000;
    rd_cycle[17446] = 1'b0;  wr_cycle[17446] = 1'b0;  addr_rom[17446]='h00000000;  wr_data_rom[17446]='h00000000;
    rd_cycle[17447] = 1'b0;  wr_cycle[17447] = 1'b0;  addr_rom[17447]='h00000000;  wr_data_rom[17447]='h00000000;
    rd_cycle[17448] = 1'b0;  wr_cycle[17448] = 1'b0;  addr_rom[17448]='h00000000;  wr_data_rom[17448]='h00000000;
    rd_cycle[17449] = 1'b0;  wr_cycle[17449] = 1'b0;  addr_rom[17449]='h00000000;  wr_data_rom[17449]='h00000000;
    rd_cycle[17450] = 1'b0;  wr_cycle[17450] = 1'b0;  addr_rom[17450]='h00000000;  wr_data_rom[17450]='h00000000;
    rd_cycle[17451] = 1'b0;  wr_cycle[17451] = 1'b0;  addr_rom[17451]='h00000000;  wr_data_rom[17451]='h00000000;
    rd_cycle[17452] = 1'b0;  wr_cycle[17452] = 1'b0;  addr_rom[17452]='h00000000;  wr_data_rom[17452]='h00000000;
    rd_cycle[17453] = 1'b0;  wr_cycle[17453] = 1'b0;  addr_rom[17453]='h00000000;  wr_data_rom[17453]='h00000000;
    rd_cycle[17454] = 1'b0;  wr_cycle[17454] = 1'b0;  addr_rom[17454]='h00000000;  wr_data_rom[17454]='h00000000;
    rd_cycle[17455] = 1'b0;  wr_cycle[17455] = 1'b0;  addr_rom[17455]='h00000000;  wr_data_rom[17455]='h00000000;
    rd_cycle[17456] = 1'b0;  wr_cycle[17456] = 1'b0;  addr_rom[17456]='h00000000;  wr_data_rom[17456]='h00000000;
    rd_cycle[17457] = 1'b0;  wr_cycle[17457] = 1'b0;  addr_rom[17457]='h00000000;  wr_data_rom[17457]='h00000000;
    rd_cycle[17458] = 1'b0;  wr_cycle[17458] = 1'b0;  addr_rom[17458]='h00000000;  wr_data_rom[17458]='h00000000;
    rd_cycle[17459] = 1'b0;  wr_cycle[17459] = 1'b0;  addr_rom[17459]='h00000000;  wr_data_rom[17459]='h00000000;
    rd_cycle[17460] = 1'b0;  wr_cycle[17460] = 1'b0;  addr_rom[17460]='h00000000;  wr_data_rom[17460]='h00000000;
    rd_cycle[17461] = 1'b0;  wr_cycle[17461] = 1'b0;  addr_rom[17461]='h00000000;  wr_data_rom[17461]='h00000000;
    rd_cycle[17462] = 1'b0;  wr_cycle[17462] = 1'b0;  addr_rom[17462]='h00000000;  wr_data_rom[17462]='h00000000;
    rd_cycle[17463] = 1'b0;  wr_cycle[17463] = 1'b0;  addr_rom[17463]='h00000000;  wr_data_rom[17463]='h00000000;
    rd_cycle[17464] = 1'b0;  wr_cycle[17464] = 1'b0;  addr_rom[17464]='h00000000;  wr_data_rom[17464]='h00000000;
    rd_cycle[17465] = 1'b0;  wr_cycle[17465] = 1'b0;  addr_rom[17465]='h00000000;  wr_data_rom[17465]='h00000000;
    rd_cycle[17466] = 1'b0;  wr_cycle[17466] = 1'b0;  addr_rom[17466]='h00000000;  wr_data_rom[17466]='h00000000;
    rd_cycle[17467] = 1'b0;  wr_cycle[17467] = 1'b0;  addr_rom[17467]='h00000000;  wr_data_rom[17467]='h00000000;
    rd_cycle[17468] = 1'b0;  wr_cycle[17468] = 1'b0;  addr_rom[17468]='h00000000;  wr_data_rom[17468]='h00000000;
    rd_cycle[17469] = 1'b0;  wr_cycle[17469] = 1'b0;  addr_rom[17469]='h00000000;  wr_data_rom[17469]='h00000000;
    rd_cycle[17470] = 1'b0;  wr_cycle[17470] = 1'b0;  addr_rom[17470]='h00000000;  wr_data_rom[17470]='h00000000;
    rd_cycle[17471] = 1'b0;  wr_cycle[17471] = 1'b0;  addr_rom[17471]='h00000000;  wr_data_rom[17471]='h00000000;
    rd_cycle[17472] = 1'b0;  wr_cycle[17472] = 1'b0;  addr_rom[17472]='h00000000;  wr_data_rom[17472]='h00000000;
    rd_cycle[17473] = 1'b0;  wr_cycle[17473] = 1'b0;  addr_rom[17473]='h00000000;  wr_data_rom[17473]='h00000000;
    rd_cycle[17474] = 1'b0;  wr_cycle[17474] = 1'b0;  addr_rom[17474]='h00000000;  wr_data_rom[17474]='h00000000;
    rd_cycle[17475] = 1'b0;  wr_cycle[17475] = 1'b0;  addr_rom[17475]='h00000000;  wr_data_rom[17475]='h00000000;
    rd_cycle[17476] = 1'b0;  wr_cycle[17476] = 1'b0;  addr_rom[17476]='h00000000;  wr_data_rom[17476]='h00000000;
    rd_cycle[17477] = 1'b0;  wr_cycle[17477] = 1'b0;  addr_rom[17477]='h00000000;  wr_data_rom[17477]='h00000000;
    rd_cycle[17478] = 1'b0;  wr_cycle[17478] = 1'b0;  addr_rom[17478]='h00000000;  wr_data_rom[17478]='h00000000;
    rd_cycle[17479] = 1'b0;  wr_cycle[17479] = 1'b0;  addr_rom[17479]='h00000000;  wr_data_rom[17479]='h00000000;
    rd_cycle[17480] = 1'b0;  wr_cycle[17480] = 1'b0;  addr_rom[17480]='h00000000;  wr_data_rom[17480]='h00000000;
    rd_cycle[17481] = 1'b0;  wr_cycle[17481] = 1'b0;  addr_rom[17481]='h00000000;  wr_data_rom[17481]='h00000000;
    rd_cycle[17482] = 1'b0;  wr_cycle[17482] = 1'b0;  addr_rom[17482]='h00000000;  wr_data_rom[17482]='h00000000;
    rd_cycle[17483] = 1'b0;  wr_cycle[17483] = 1'b0;  addr_rom[17483]='h00000000;  wr_data_rom[17483]='h00000000;
    rd_cycle[17484] = 1'b0;  wr_cycle[17484] = 1'b0;  addr_rom[17484]='h00000000;  wr_data_rom[17484]='h00000000;
    rd_cycle[17485] = 1'b0;  wr_cycle[17485] = 1'b0;  addr_rom[17485]='h00000000;  wr_data_rom[17485]='h00000000;
    rd_cycle[17486] = 1'b0;  wr_cycle[17486] = 1'b0;  addr_rom[17486]='h00000000;  wr_data_rom[17486]='h00000000;
    rd_cycle[17487] = 1'b0;  wr_cycle[17487] = 1'b0;  addr_rom[17487]='h00000000;  wr_data_rom[17487]='h00000000;
    rd_cycle[17488] = 1'b0;  wr_cycle[17488] = 1'b0;  addr_rom[17488]='h00000000;  wr_data_rom[17488]='h00000000;
    rd_cycle[17489] = 1'b0;  wr_cycle[17489] = 1'b0;  addr_rom[17489]='h00000000;  wr_data_rom[17489]='h00000000;
    rd_cycle[17490] = 1'b0;  wr_cycle[17490] = 1'b0;  addr_rom[17490]='h00000000;  wr_data_rom[17490]='h00000000;
    rd_cycle[17491] = 1'b0;  wr_cycle[17491] = 1'b0;  addr_rom[17491]='h00000000;  wr_data_rom[17491]='h00000000;
    rd_cycle[17492] = 1'b0;  wr_cycle[17492] = 1'b0;  addr_rom[17492]='h00000000;  wr_data_rom[17492]='h00000000;
    rd_cycle[17493] = 1'b0;  wr_cycle[17493] = 1'b0;  addr_rom[17493]='h00000000;  wr_data_rom[17493]='h00000000;
    rd_cycle[17494] = 1'b0;  wr_cycle[17494] = 1'b0;  addr_rom[17494]='h00000000;  wr_data_rom[17494]='h00000000;
    rd_cycle[17495] = 1'b0;  wr_cycle[17495] = 1'b0;  addr_rom[17495]='h00000000;  wr_data_rom[17495]='h00000000;
    rd_cycle[17496] = 1'b0;  wr_cycle[17496] = 1'b0;  addr_rom[17496]='h00000000;  wr_data_rom[17496]='h00000000;
    rd_cycle[17497] = 1'b0;  wr_cycle[17497] = 1'b0;  addr_rom[17497]='h00000000;  wr_data_rom[17497]='h00000000;
    rd_cycle[17498] = 1'b0;  wr_cycle[17498] = 1'b0;  addr_rom[17498]='h00000000;  wr_data_rom[17498]='h00000000;
    rd_cycle[17499] = 1'b0;  wr_cycle[17499] = 1'b0;  addr_rom[17499]='h00000000;  wr_data_rom[17499]='h00000000;
    rd_cycle[17500] = 1'b0;  wr_cycle[17500] = 1'b0;  addr_rom[17500]='h00000000;  wr_data_rom[17500]='h00000000;
    rd_cycle[17501] = 1'b0;  wr_cycle[17501] = 1'b0;  addr_rom[17501]='h00000000;  wr_data_rom[17501]='h00000000;
    rd_cycle[17502] = 1'b0;  wr_cycle[17502] = 1'b0;  addr_rom[17502]='h00000000;  wr_data_rom[17502]='h00000000;
    rd_cycle[17503] = 1'b0;  wr_cycle[17503] = 1'b0;  addr_rom[17503]='h00000000;  wr_data_rom[17503]='h00000000;
    rd_cycle[17504] = 1'b0;  wr_cycle[17504] = 1'b0;  addr_rom[17504]='h00000000;  wr_data_rom[17504]='h00000000;
    rd_cycle[17505] = 1'b0;  wr_cycle[17505] = 1'b0;  addr_rom[17505]='h00000000;  wr_data_rom[17505]='h00000000;
    rd_cycle[17506] = 1'b0;  wr_cycle[17506] = 1'b0;  addr_rom[17506]='h00000000;  wr_data_rom[17506]='h00000000;
    rd_cycle[17507] = 1'b0;  wr_cycle[17507] = 1'b0;  addr_rom[17507]='h00000000;  wr_data_rom[17507]='h00000000;
    rd_cycle[17508] = 1'b0;  wr_cycle[17508] = 1'b0;  addr_rom[17508]='h00000000;  wr_data_rom[17508]='h00000000;
    rd_cycle[17509] = 1'b0;  wr_cycle[17509] = 1'b0;  addr_rom[17509]='h00000000;  wr_data_rom[17509]='h00000000;
    rd_cycle[17510] = 1'b0;  wr_cycle[17510] = 1'b0;  addr_rom[17510]='h00000000;  wr_data_rom[17510]='h00000000;
    rd_cycle[17511] = 1'b0;  wr_cycle[17511] = 1'b0;  addr_rom[17511]='h00000000;  wr_data_rom[17511]='h00000000;
    rd_cycle[17512] = 1'b0;  wr_cycle[17512] = 1'b0;  addr_rom[17512]='h00000000;  wr_data_rom[17512]='h00000000;
    rd_cycle[17513] = 1'b0;  wr_cycle[17513] = 1'b0;  addr_rom[17513]='h00000000;  wr_data_rom[17513]='h00000000;
    rd_cycle[17514] = 1'b0;  wr_cycle[17514] = 1'b0;  addr_rom[17514]='h00000000;  wr_data_rom[17514]='h00000000;
    rd_cycle[17515] = 1'b0;  wr_cycle[17515] = 1'b0;  addr_rom[17515]='h00000000;  wr_data_rom[17515]='h00000000;
    rd_cycle[17516] = 1'b0;  wr_cycle[17516] = 1'b0;  addr_rom[17516]='h00000000;  wr_data_rom[17516]='h00000000;
    rd_cycle[17517] = 1'b0;  wr_cycle[17517] = 1'b0;  addr_rom[17517]='h00000000;  wr_data_rom[17517]='h00000000;
    rd_cycle[17518] = 1'b0;  wr_cycle[17518] = 1'b0;  addr_rom[17518]='h00000000;  wr_data_rom[17518]='h00000000;
    rd_cycle[17519] = 1'b0;  wr_cycle[17519] = 1'b0;  addr_rom[17519]='h00000000;  wr_data_rom[17519]='h00000000;
    rd_cycle[17520] = 1'b0;  wr_cycle[17520] = 1'b0;  addr_rom[17520]='h00000000;  wr_data_rom[17520]='h00000000;
    rd_cycle[17521] = 1'b0;  wr_cycle[17521] = 1'b0;  addr_rom[17521]='h00000000;  wr_data_rom[17521]='h00000000;
    rd_cycle[17522] = 1'b0;  wr_cycle[17522] = 1'b0;  addr_rom[17522]='h00000000;  wr_data_rom[17522]='h00000000;
    rd_cycle[17523] = 1'b0;  wr_cycle[17523] = 1'b0;  addr_rom[17523]='h00000000;  wr_data_rom[17523]='h00000000;
    rd_cycle[17524] = 1'b0;  wr_cycle[17524] = 1'b0;  addr_rom[17524]='h00000000;  wr_data_rom[17524]='h00000000;
    rd_cycle[17525] = 1'b0;  wr_cycle[17525] = 1'b0;  addr_rom[17525]='h00000000;  wr_data_rom[17525]='h00000000;
    rd_cycle[17526] = 1'b0;  wr_cycle[17526] = 1'b0;  addr_rom[17526]='h00000000;  wr_data_rom[17526]='h00000000;
    rd_cycle[17527] = 1'b0;  wr_cycle[17527] = 1'b0;  addr_rom[17527]='h00000000;  wr_data_rom[17527]='h00000000;
    rd_cycle[17528] = 1'b0;  wr_cycle[17528] = 1'b0;  addr_rom[17528]='h00000000;  wr_data_rom[17528]='h00000000;
    rd_cycle[17529] = 1'b0;  wr_cycle[17529] = 1'b0;  addr_rom[17529]='h00000000;  wr_data_rom[17529]='h00000000;
    rd_cycle[17530] = 1'b0;  wr_cycle[17530] = 1'b0;  addr_rom[17530]='h00000000;  wr_data_rom[17530]='h00000000;
    rd_cycle[17531] = 1'b0;  wr_cycle[17531] = 1'b0;  addr_rom[17531]='h00000000;  wr_data_rom[17531]='h00000000;
    rd_cycle[17532] = 1'b0;  wr_cycle[17532] = 1'b0;  addr_rom[17532]='h00000000;  wr_data_rom[17532]='h00000000;
    rd_cycle[17533] = 1'b0;  wr_cycle[17533] = 1'b0;  addr_rom[17533]='h00000000;  wr_data_rom[17533]='h00000000;
    rd_cycle[17534] = 1'b0;  wr_cycle[17534] = 1'b0;  addr_rom[17534]='h00000000;  wr_data_rom[17534]='h00000000;
    rd_cycle[17535] = 1'b0;  wr_cycle[17535] = 1'b0;  addr_rom[17535]='h00000000;  wr_data_rom[17535]='h00000000;
    rd_cycle[17536] = 1'b0;  wr_cycle[17536] = 1'b0;  addr_rom[17536]='h00000000;  wr_data_rom[17536]='h00000000;
    rd_cycle[17537] = 1'b0;  wr_cycle[17537] = 1'b0;  addr_rom[17537]='h00000000;  wr_data_rom[17537]='h00000000;
    rd_cycle[17538] = 1'b0;  wr_cycle[17538] = 1'b0;  addr_rom[17538]='h00000000;  wr_data_rom[17538]='h00000000;
    rd_cycle[17539] = 1'b0;  wr_cycle[17539] = 1'b0;  addr_rom[17539]='h00000000;  wr_data_rom[17539]='h00000000;
    rd_cycle[17540] = 1'b0;  wr_cycle[17540] = 1'b0;  addr_rom[17540]='h00000000;  wr_data_rom[17540]='h00000000;
    rd_cycle[17541] = 1'b0;  wr_cycle[17541] = 1'b0;  addr_rom[17541]='h00000000;  wr_data_rom[17541]='h00000000;
    rd_cycle[17542] = 1'b0;  wr_cycle[17542] = 1'b0;  addr_rom[17542]='h00000000;  wr_data_rom[17542]='h00000000;
    rd_cycle[17543] = 1'b0;  wr_cycle[17543] = 1'b0;  addr_rom[17543]='h00000000;  wr_data_rom[17543]='h00000000;
    rd_cycle[17544] = 1'b0;  wr_cycle[17544] = 1'b0;  addr_rom[17544]='h00000000;  wr_data_rom[17544]='h00000000;
    rd_cycle[17545] = 1'b0;  wr_cycle[17545] = 1'b0;  addr_rom[17545]='h00000000;  wr_data_rom[17545]='h00000000;
    rd_cycle[17546] = 1'b0;  wr_cycle[17546] = 1'b0;  addr_rom[17546]='h00000000;  wr_data_rom[17546]='h00000000;
    rd_cycle[17547] = 1'b0;  wr_cycle[17547] = 1'b0;  addr_rom[17547]='h00000000;  wr_data_rom[17547]='h00000000;
    rd_cycle[17548] = 1'b0;  wr_cycle[17548] = 1'b0;  addr_rom[17548]='h00000000;  wr_data_rom[17548]='h00000000;
    rd_cycle[17549] = 1'b0;  wr_cycle[17549] = 1'b0;  addr_rom[17549]='h00000000;  wr_data_rom[17549]='h00000000;
    rd_cycle[17550] = 1'b0;  wr_cycle[17550] = 1'b0;  addr_rom[17550]='h00000000;  wr_data_rom[17550]='h00000000;
    rd_cycle[17551] = 1'b0;  wr_cycle[17551] = 1'b0;  addr_rom[17551]='h00000000;  wr_data_rom[17551]='h00000000;
    rd_cycle[17552] = 1'b0;  wr_cycle[17552] = 1'b0;  addr_rom[17552]='h00000000;  wr_data_rom[17552]='h00000000;
    rd_cycle[17553] = 1'b0;  wr_cycle[17553] = 1'b0;  addr_rom[17553]='h00000000;  wr_data_rom[17553]='h00000000;
    rd_cycle[17554] = 1'b0;  wr_cycle[17554] = 1'b0;  addr_rom[17554]='h00000000;  wr_data_rom[17554]='h00000000;
    rd_cycle[17555] = 1'b0;  wr_cycle[17555] = 1'b0;  addr_rom[17555]='h00000000;  wr_data_rom[17555]='h00000000;
    rd_cycle[17556] = 1'b0;  wr_cycle[17556] = 1'b0;  addr_rom[17556]='h00000000;  wr_data_rom[17556]='h00000000;
    rd_cycle[17557] = 1'b0;  wr_cycle[17557] = 1'b0;  addr_rom[17557]='h00000000;  wr_data_rom[17557]='h00000000;
    rd_cycle[17558] = 1'b0;  wr_cycle[17558] = 1'b0;  addr_rom[17558]='h00000000;  wr_data_rom[17558]='h00000000;
    rd_cycle[17559] = 1'b0;  wr_cycle[17559] = 1'b0;  addr_rom[17559]='h00000000;  wr_data_rom[17559]='h00000000;
    rd_cycle[17560] = 1'b0;  wr_cycle[17560] = 1'b0;  addr_rom[17560]='h00000000;  wr_data_rom[17560]='h00000000;
    rd_cycle[17561] = 1'b0;  wr_cycle[17561] = 1'b0;  addr_rom[17561]='h00000000;  wr_data_rom[17561]='h00000000;
    rd_cycle[17562] = 1'b0;  wr_cycle[17562] = 1'b0;  addr_rom[17562]='h00000000;  wr_data_rom[17562]='h00000000;
    rd_cycle[17563] = 1'b0;  wr_cycle[17563] = 1'b0;  addr_rom[17563]='h00000000;  wr_data_rom[17563]='h00000000;
    rd_cycle[17564] = 1'b0;  wr_cycle[17564] = 1'b0;  addr_rom[17564]='h00000000;  wr_data_rom[17564]='h00000000;
    rd_cycle[17565] = 1'b0;  wr_cycle[17565] = 1'b0;  addr_rom[17565]='h00000000;  wr_data_rom[17565]='h00000000;
    rd_cycle[17566] = 1'b0;  wr_cycle[17566] = 1'b0;  addr_rom[17566]='h00000000;  wr_data_rom[17566]='h00000000;
    rd_cycle[17567] = 1'b0;  wr_cycle[17567] = 1'b0;  addr_rom[17567]='h00000000;  wr_data_rom[17567]='h00000000;
    rd_cycle[17568] = 1'b0;  wr_cycle[17568] = 1'b0;  addr_rom[17568]='h00000000;  wr_data_rom[17568]='h00000000;
    rd_cycle[17569] = 1'b0;  wr_cycle[17569] = 1'b0;  addr_rom[17569]='h00000000;  wr_data_rom[17569]='h00000000;
    rd_cycle[17570] = 1'b0;  wr_cycle[17570] = 1'b0;  addr_rom[17570]='h00000000;  wr_data_rom[17570]='h00000000;
    rd_cycle[17571] = 1'b0;  wr_cycle[17571] = 1'b0;  addr_rom[17571]='h00000000;  wr_data_rom[17571]='h00000000;
    rd_cycle[17572] = 1'b0;  wr_cycle[17572] = 1'b0;  addr_rom[17572]='h00000000;  wr_data_rom[17572]='h00000000;
    rd_cycle[17573] = 1'b0;  wr_cycle[17573] = 1'b0;  addr_rom[17573]='h00000000;  wr_data_rom[17573]='h00000000;
    rd_cycle[17574] = 1'b0;  wr_cycle[17574] = 1'b0;  addr_rom[17574]='h00000000;  wr_data_rom[17574]='h00000000;
    rd_cycle[17575] = 1'b0;  wr_cycle[17575] = 1'b0;  addr_rom[17575]='h00000000;  wr_data_rom[17575]='h00000000;
    rd_cycle[17576] = 1'b0;  wr_cycle[17576] = 1'b0;  addr_rom[17576]='h00000000;  wr_data_rom[17576]='h00000000;
    rd_cycle[17577] = 1'b0;  wr_cycle[17577] = 1'b0;  addr_rom[17577]='h00000000;  wr_data_rom[17577]='h00000000;
    rd_cycle[17578] = 1'b0;  wr_cycle[17578] = 1'b0;  addr_rom[17578]='h00000000;  wr_data_rom[17578]='h00000000;
    rd_cycle[17579] = 1'b0;  wr_cycle[17579] = 1'b0;  addr_rom[17579]='h00000000;  wr_data_rom[17579]='h00000000;
    rd_cycle[17580] = 1'b0;  wr_cycle[17580] = 1'b0;  addr_rom[17580]='h00000000;  wr_data_rom[17580]='h00000000;
    rd_cycle[17581] = 1'b0;  wr_cycle[17581] = 1'b0;  addr_rom[17581]='h00000000;  wr_data_rom[17581]='h00000000;
    rd_cycle[17582] = 1'b0;  wr_cycle[17582] = 1'b0;  addr_rom[17582]='h00000000;  wr_data_rom[17582]='h00000000;
    rd_cycle[17583] = 1'b0;  wr_cycle[17583] = 1'b0;  addr_rom[17583]='h00000000;  wr_data_rom[17583]='h00000000;
    rd_cycle[17584] = 1'b0;  wr_cycle[17584] = 1'b0;  addr_rom[17584]='h00000000;  wr_data_rom[17584]='h00000000;
    rd_cycle[17585] = 1'b0;  wr_cycle[17585] = 1'b0;  addr_rom[17585]='h00000000;  wr_data_rom[17585]='h00000000;
    rd_cycle[17586] = 1'b0;  wr_cycle[17586] = 1'b0;  addr_rom[17586]='h00000000;  wr_data_rom[17586]='h00000000;
    rd_cycle[17587] = 1'b0;  wr_cycle[17587] = 1'b0;  addr_rom[17587]='h00000000;  wr_data_rom[17587]='h00000000;
    rd_cycle[17588] = 1'b0;  wr_cycle[17588] = 1'b0;  addr_rom[17588]='h00000000;  wr_data_rom[17588]='h00000000;
    rd_cycle[17589] = 1'b0;  wr_cycle[17589] = 1'b0;  addr_rom[17589]='h00000000;  wr_data_rom[17589]='h00000000;
    rd_cycle[17590] = 1'b0;  wr_cycle[17590] = 1'b0;  addr_rom[17590]='h00000000;  wr_data_rom[17590]='h00000000;
    rd_cycle[17591] = 1'b0;  wr_cycle[17591] = 1'b0;  addr_rom[17591]='h00000000;  wr_data_rom[17591]='h00000000;
    rd_cycle[17592] = 1'b0;  wr_cycle[17592] = 1'b0;  addr_rom[17592]='h00000000;  wr_data_rom[17592]='h00000000;
    rd_cycle[17593] = 1'b0;  wr_cycle[17593] = 1'b0;  addr_rom[17593]='h00000000;  wr_data_rom[17593]='h00000000;
    rd_cycle[17594] = 1'b0;  wr_cycle[17594] = 1'b0;  addr_rom[17594]='h00000000;  wr_data_rom[17594]='h00000000;
    rd_cycle[17595] = 1'b0;  wr_cycle[17595] = 1'b0;  addr_rom[17595]='h00000000;  wr_data_rom[17595]='h00000000;
    rd_cycle[17596] = 1'b0;  wr_cycle[17596] = 1'b0;  addr_rom[17596]='h00000000;  wr_data_rom[17596]='h00000000;
    rd_cycle[17597] = 1'b0;  wr_cycle[17597] = 1'b0;  addr_rom[17597]='h00000000;  wr_data_rom[17597]='h00000000;
    rd_cycle[17598] = 1'b0;  wr_cycle[17598] = 1'b0;  addr_rom[17598]='h00000000;  wr_data_rom[17598]='h00000000;
    rd_cycle[17599] = 1'b0;  wr_cycle[17599] = 1'b0;  addr_rom[17599]='h00000000;  wr_data_rom[17599]='h00000000;
    rd_cycle[17600] = 1'b0;  wr_cycle[17600] = 1'b0;  addr_rom[17600]='h00000000;  wr_data_rom[17600]='h00000000;
    rd_cycle[17601] = 1'b0;  wr_cycle[17601] = 1'b0;  addr_rom[17601]='h00000000;  wr_data_rom[17601]='h00000000;
    rd_cycle[17602] = 1'b0;  wr_cycle[17602] = 1'b0;  addr_rom[17602]='h00000000;  wr_data_rom[17602]='h00000000;
    rd_cycle[17603] = 1'b0;  wr_cycle[17603] = 1'b0;  addr_rom[17603]='h00000000;  wr_data_rom[17603]='h00000000;
    rd_cycle[17604] = 1'b0;  wr_cycle[17604] = 1'b0;  addr_rom[17604]='h00000000;  wr_data_rom[17604]='h00000000;
    rd_cycle[17605] = 1'b0;  wr_cycle[17605] = 1'b0;  addr_rom[17605]='h00000000;  wr_data_rom[17605]='h00000000;
    rd_cycle[17606] = 1'b0;  wr_cycle[17606] = 1'b0;  addr_rom[17606]='h00000000;  wr_data_rom[17606]='h00000000;
    rd_cycle[17607] = 1'b0;  wr_cycle[17607] = 1'b0;  addr_rom[17607]='h00000000;  wr_data_rom[17607]='h00000000;
    rd_cycle[17608] = 1'b0;  wr_cycle[17608] = 1'b0;  addr_rom[17608]='h00000000;  wr_data_rom[17608]='h00000000;
    rd_cycle[17609] = 1'b0;  wr_cycle[17609] = 1'b0;  addr_rom[17609]='h00000000;  wr_data_rom[17609]='h00000000;
    rd_cycle[17610] = 1'b0;  wr_cycle[17610] = 1'b0;  addr_rom[17610]='h00000000;  wr_data_rom[17610]='h00000000;
    rd_cycle[17611] = 1'b0;  wr_cycle[17611] = 1'b0;  addr_rom[17611]='h00000000;  wr_data_rom[17611]='h00000000;
    rd_cycle[17612] = 1'b0;  wr_cycle[17612] = 1'b0;  addr_rom[17612]='h00000000;  wr_data_rom[17612]='h00000000;
    rd_cycle[17613] = 1'b0;  wr_cycle[17613] = 1'b0;  addr_rom[17613]='h00000000;  wr_data_rom[17613]='h00000000;
    rd_cycle[17614] = 1'b0;  wr_cycle[17614] = 1'b0;  addr_rom[17614]='h00000000;  wr_data_rom[17614]='h00000000;
    rd_cycle[17615] = 1'b0;  wr_cycle[17615] = 1'b0;  addr_rom[17615]='h00000000;  wr_data_rom[17615]='h00000000;
    rd_cycle[17616] = 1'b0;  wr_cycle[17616] = 1'b0;  addr_rom[17616]='h00000000;  wr_data_rom[17616]='h00000000;
    rd_cycle[17617] = 1'b0;  wr_cycle[17617] = 1'b0;  addr_rom[17617]='h00000000;  wr_data_rom[17617]='h00000000;
    rd_cycle[17618] = 1'b0;  wr_cycle[17618] = 1'b0;  addr_rom[17618]='h00000000;  wr_data_rom[17618]='h00000000;
    rd_cycle[17619] = 1'b0;  wr_cycle[17619] = 1'b0;  addr_rom[17619]='h00000000;  wr_data_rom[17619]='h00000000;
    rd_cycle[17620] = 1'b0;  wr_cycle[17620] = 1'b0;  addr_rom[17620]='h00000000;  wr_data_rom[17620]='h00000000;
    rd_cycle[17621] = 1'b0;  wr_cycle[17621] = 1'b0;  addr_rom[17621]='h00000000;  wr_data_rom[17621]='h00000000;
    rd_cycle[17622] = 1'b0;  wr_cycle[17622] = 1'b0;  addr_rom[17622]='h00000000;  wr_data_rom[17622]='h00000000;
    rd_cycle[17623] = 1'b0;  wr_cycle[17623] = 1'b0;  addr_rom[17623]='h00000000;  wr_data_rom[17623]='h00000000;
    rd_cycle[17624] = 1'b0;  wr_cycle[17624] = 1'b0;  addr_rom[17624]='h00000000;  wr_data_rom[17624]='h00000000;
    rd_cycle[17625] = 1'b0;  wr_cycle[17625] = 1'b0;  addr_rom[17625]='h00000000;  wr_data_rom[17625]='h00000000;
    rd_cycle[17626] = 1'b0;  wr_cycle[17626] = 1'b0;  addr_rom[17626]='h00000000;  wr_data_rom[17626]='h00000000;
    rd_cycle[17627] = 1'b0;  wr_cycle[17627] = 1'b0;  addr_rom[17627]='h00000000;  wr_data_rom[17627]='h00000000;
    rd_cycle[17628] = 1'b0;  wr_cycle[17628] = 1'b0;  addr_rom[17628]='h00000000;  wr_data_rom[17628]='h00000000;
    rd_cycle[17629] = 1'b0;  wr_cycle[17629] = 1'b0;  addr_rom[17629]='h00000000;  wr_data_rom[17629]='h00000000;
    rd_cycle[17630] = 1'b0;  wr_cycle[17630] = 1'b0;  addr_rom[17630]='h00000000;  wr_data_rom[17630]='h00000000;
    rd_cycle[17631] = 1'b0;  wr_cycle[17631] = 1'b0;  addr_rom[17631]='h00000000;  wr_data_rom[17631]='h00000000;
    rd_cycle[17632] = 1'b0;  wr_cycle[17632] = 1'b0;  addr_rom[17632]='h00000000;  wr_data_rom[17632]='h00000000;
    rd_cycle[17633] = 1'b0;  wr_cycle[17633] = 1'b0;  addr_rom[17633]='h00000000;  wr_data_rom[17633]='h00000000;
    rd_cycle[17634] = 1'b0;  wr_cycle[17634] = 1'b0;  addr_rom[17634]='h00000000;  wr_data_rom[17634]='h00000000;
    rd_cycle[17635] = 1'b0;  wr_cycle[17635] = 1'b0;  addr_rom[17635]='h00000000;  wr_data_rom[17635]='h00000000;
    rd_cycle[17636] = 1'b0;  wr_cycle[17636] = 1'b0;  addr_rom[17636]='h00000000;  wr_data_rom[17636]='h00000000;
    rd_cycle[17637] = 1'b0;  wr_cycle[17637] = 1'b0;  addr_rom[17637]='h00000000;  wr_data_rom[17637]='h00000000;
    rd_cycle[17638] = 1'b0;  wr_cycle[17638] = 1'b0;  addr_rom[17638]='h00000000;  wr_data_rom[17638]='h00000000;
    rd_cycle[17639] = 1'b0;  wr_cycle[17639] = 1'b0;  addr_rom[17639]='h00000000;  wr_data_rom[17639]='h00000000;
    rd_cycle[17640] = 1'b0;  wr_cycle[17640] = 1'b0;  addr_rom[17640]='h00000000;  wr_data_rom[17640]='h00000000;
    rd_cycle[17641] = 1'b0;  wr_cycle[17641] = 1'b0;  addr_rom[17641]='h00000000;  wr_data_rom[17641]='h00000000;
    rd_cycle[17642] = 1'b0;  wr_cycle[17642] = 1'b0;  addr_rom[17642]='h00000000;  wr_data_rom[17642]='h00000000;
    rd_cycle[17643] = 1'b0;  wr_cycle[17643] = 1'b0;  addr_rom[17643]='h00000000;  wr_data_rom[17643]='h00000000;
    rd_cycle[17644] = 1'b0;  wr_cycle[17644] = 1'b0;  addr_rom[17644]='h00000000;  wr_data_rom[17644]='h00000000;
    rd_cycle[17645] = 1'b0;  wr_cycle[17645] = 1'b0;  addr_rom[17645]='h00000000;  wr_data_rom[17645]='h00000000;
    rd_cycle[17646] = 1'b0;  wr_cycle[17646] = 1'b0;  addr_rom[17646]='h00000000;  wr_data_rom[17646]='h00000000;
    rd_cycle[17647] = 1'b0;  wr_cycle[17647] = 1'b0;  addr_rom[17647]='h00000000;  wr_data_rom[17647]='h00000000;
    rd_cycle[17648] = 1'b0;  wr_cycle[17648] = 1'b0;  addr_rom[17648]='h00000000;  wr_data_rom[17648]='h00000000;
    rd_cycle[17649] = 1'b0;  wr_cycle[17649] = 1'b0;  addr_rom[17649]='h00000000;  wr_data_rom[17649]='h00000000;
    rd_cycle[17650] = 1'b0;  wr_cycle[17650] = 1'b0;  addr_rom[17650]='h00000000;  wr_data_rom[17650]='h00000000;
    rd_cycle[17651] = 1'b0;  wr_cycle[17651] = 1'b0;  addr_rom[17651]='h00000000;  wr_data_rom[17651]='h00000000;
    rd_cycle[17652] = 1'b0;  wr_cycle[17652] = 1'b0;  addr_rom[17652]='h00000000;  wr_data_rom[17652]='h00000000;
    rd_cycle[17653] = 1'b0;  wr_cycle[17653] = 1'b0;  addr_rom[17653]='h00000000;  wr_data_rom[17653]='h00000000;
    rd_cycle[17654] = 1'b0;  wr_cycle[17654] = 1'b0;  addr_rom[17654]='h00000000;  wr_data_rom[17654]='h00000000;
    rd_cycle[17655] = 1'b0;  wr_cycle[17655] = 1'b0;  addr_rom[17655]='h00000000;  wr_data_rom[17655]='h00000000;
    rd_cycle[17656] = 1'b0;  wr_cycle[17656] = 1'b0;  addr_rom[17656]='h00000000;  wr_data_rom[17656]='h00000000;
    rd_cycle[17657] = 1'b0;  wr_cycle[17657] = 1'b0;  addr_rom[17657]='h00000000;  wr_data_rom[17657]='h00000000;
    rd_cycle[17658] = 1'b0;  wr_cycle[17658] = 1'b0;  addr_rom[17658]='h00000000;  wr_data_rom[17658]='h00000000;
    rd_cycle[17659] = 1'b0;  wr_cycle[17659] = 1'b0;  addr_rom[17659]='h00000000;  wr_data_rom[17659]='h00000000;
    rd_cycle[17660] = 1'b0;  wr_cycle[17660] = 1'b0;  addr_rom[17660]='h00000000;  wr_data_rom[17660]='h00000000;
    rd_cycle[17661] = 1'b0;  wr_cycle[17661] = 1'b0;  addr_rom[17661]='h00000000;  wr_data_rom[17661]='h00000000;
    rd_cycle[17662] = 1'b0;  wr_cycle[17662] = 1'b0;  addr_rom[17662]='h00000000;  wr_data_rom[17662]='h00000000;
    rd_cycle[17663] = 1'b0;  wr_cycle[17663] = 1'b0;  addr_rom[17663]='h00000000;  wr_data_rom[17663]='h00000000;
    rd_cycle[17664] = 1'b0;  wr_cycle[17664] = 1'b0;  addr_rom[17664]='h00000000;  wr_data_rom[17664]='h00000000;
    rd_cycle[17665] = 1'b0;  wr_cycle[17665] = 1'b0;  addr_rom[17665]='h00000000;  wr_data_rom[17665]='h00000000;
    rd_cycle[17666] = 1'b0;  wr_cycle[17666] = 1'b0;  addr_rom[17666]='h00000000;  wr_data_rom[17666]='h00000000;
    rd_cycle[17667] = 1'b0;  wr_cycle[17667] = 1'b0;  addr_rom[17667]='h00000000;  wr_data_rom[17667]='h00000000;
    rd_cycle[17668] = 1'b0;  wr_cycle[17668] = 1'b0;  addr_rom[17668]='h00000000;  wr_data_rom[17668]='h00000000;
    rd_cycle[17669] = 1'b0;  wr_cycle[17669] = 1'b0;  addr_rom[17669]='h00000000;  wr_data_rom[17669]='h00000000;
    rd_cycle[17670] = 1'b0;  wr_cycle[17670] = 1'b0;  addr_rom[17670]='h00000000;  wr_data_rom[17670]='h00000000;
    rd_cycle[17671] = 1'b0;  wr_cycle[17671] = 1'b0;  addr_rom[17671]='h00000000;  wr_data_rom[17671]='h00000000;
    rd_cycle[17672] = 1'b0;  wr_cycle[17672] = 1'b0;  addr_rom[17672]='h00000000;  wr_data_rom[17672]='h00000000;
    rd_cycle[17673] = 1'b0;  wr_cycle[17673] = 1'b0;  addr_rom[17673]='h00000000;  wr_data_rom[17673]='h00000000;
    rd_cycle[17674] = 1'b0;  wr_cycle[17674] = 1'b0;  addr_rom[17674]='h00000000;  wr_data_rom[17674]='h00000000;
    rd_cycle[17675] = 1'b0;  wr_cycle[17675] = 1'b0;  addr_rom[17675]='h00000000;  wr_data_rom[17675]='h00000000;
    rd_cycle[17676] = 1'b0;  wr_cycle[17676] = 1'b0;  addr_rom[17676]='h00000000;  wr_data_rom[17676]='h00000000;
    rd_cycle[17677] = 1'b0;  wr_cycle[17677] = 1'b0;  addr_rom[17677]='h00000000;  wr_data_rom[17677]='h00000000;
    rd_cycle[17678] = 1'b0;  wr_cycle[17678] = 1'b0;  addr_rom[17678]='h00000000;  wr_data_rom[17678]='h00000000;
    rd_cycle[17679] = 1'b0;  wr_cycle[17679] = 1'b0;  addr_rom[17679]='h00000000;  wr_data_rom[17679]='h00000000;
    rd_cycle[17680] = 1'b0;  wr_cycle[17680] = 1'b0;  addr_rom[17680]='h00000000;  wr_data_rom[17680]='h00000000;
    rd_cycle[17681] = 1'b0;  wr_cycle[17681] = 1'b0;  addr_rom[17681]='h00000000;  wr_data_rom[17681]='h00000000;
    rd_cycle[17682] = 1'b0;  wr_cycle[17682] = 1'b0;  addr_rom[17682]='h00000000;  wr_data_rom[17682]='h00000000;
    rd_cycle[17683] = 1'b0;  wr_cycle[17683] = 1'b0;  addr_rom[17683]='h00000000;  wr_data_rom[17683]='h00000000;
    rd_cycle[17684] = 1'b0;  wr_cycle[17684] = 1'b0;  addr_rom[17684]='h00000000;  wr_data_rom[17684]='h00000000;
    rd_cycle[17685] = 1'b0;  wr_cycle[17685] = 1'b0;  addr_rom[17685]='h00000000;  wr_data_rom[17685]='h00000000;
    rd_cycle[17686] = 1'b0;  wr_cycle[17686] = 1'b0;  addr_rom[17686]='h00000000;  wr_data_rom[17686]='h00000000;
    rd_cycle[17687] = 1'b0;  wr_cycle[17687] = 1'b0;  addr_rom[17687]='h00000000;  wr_data_rom[17687]='h00000000;
    rd_cycle[17688] = 1'b0;  wr_cycle[17688] = 1'b0;  addr_rom[17688]='h00000000;  wr_data_rom[17688]='h00000000;
    rd_cycle[17689] = 1'b0;  wr_cycle[17689] = 1'b0;  addr_rom[17689]='h00000000;  wr_data_rom[17689]='h00000000;
    rd_cycle[17690] = 1'b0;  wr_cycle[17690] = 1'b0;  addr_rom[17690]='h00000000;  wr_data_rom[17690]='h00000000;
    rd_cycle[17691] = 1'b0;  wr_cycle[17691] = 1'b0;  addr_rom[17691]='h00000000;  wr_data_rom[17691]='h00000000;
    rd_cycle[17692] = 1'b0;  wr_cycle[17692] = 1'b0;  addr_rom[17692]='h00000000;  wr_data_rom[17692]='h00000000;
    rd_cycle[17693] = 1'b0;  wr_cycle[17693] = 1'b0;  addr_rom[17693]='h00000000;  wr_data_rom[17693]='h00000000;
    rd_cycle[17694] = 1'b0;  wr_cycle[17694] = 1'b0;  addr_rom[17694]='h00000000;  wr_data_rom[17694]='h00000000;
    rd_cycle[17695] = 1'b0;  wr_cycle[17695] = 1'b0;  addr_rom[17695]='h00000000;  wr_data_rom[17695]='h00000000;
    rd_cycle[17696] = 1'b0;  wr_cycle[17696] = 1'b0;  addr_rom[17696]='h00000000;  wr_data_rom[17696]='h00000000;
    rd_cycle[17697] = 1'b0;  wr_cycle[17697] = 1'b0;  addr_rom[17697]='h00000000;  wr_data_rom[17697]='h00000000;
    rd_cycle[17698] = 1'b0;  wr_cycle[17698] = 1'b0;  addr_rom[17698]='h00000000;  wr_data_rom[17698]='h00000000;
    rd_cycle[17699] = 1'b0;  wr_cycle[17699] = 1'b0;  addr_rom[17699]='h00000000;  wr_data_rom[17699]='h00000000;
    rd_cycle[17700] = 1'b0;  wr_cycle[17700] = 1'b0;  addr_rom[17700]='h00000000;  wr_data_rom[17700]='h00000000;
    rd_cycle[17701] = 1'b0;  wr_cycle[17701] = 1'b0;  addr_rom[17701]='h00000000;  wr_data_rom[17701]='h00000000;
    rd_cycle[17702] = 1'b0;  wr_cycle[17702] = 1'b0;  addr_rom[17702]='h00000000;  wr_data_rom[17702]='h00000000;
    rd_cycle[17703] = 1'b0;  wr_cycle[17703] = 1'b0;  addr_rom[17703]='h00000000;  wr_data_rom[17703]='h00000000;
    rd_cycle[17704] = 1'b0;  wr_cycle[17704] = 1'b0;  addr_rom[17704]='h00000000;  wr_data_rom[17704]='h00000000;
    rd_cycle[17705] = 1'b0;  wr_cycle[17705] = 1'b0;  addr_rom[17705]='h00000000;  wr_data_rom[17705]='h00000000;
    rd_cycle[17706] = 1'b0;  wr_cycle[17706] = 1'b0;  addr_rom[17706]='h00000000;  wr_data_rom[17706]='h00000000;
    rd_cycle[17707] = 1'b0;  wr_cycle[17707] = 1'b0;  addr_rom[17707]='h00000000;  wr_data_rom[17707]='h00000000;
    rd_cycle[17708] = 1'b0;  wr_cycle[17708] = 1'b0;  addr_rom[17708]='h00000000;  wr_data_rom[17708]='h00000000;
    rd_cycle[17709] = 1'b0;  wr_cycle[17709] = 1'b0;  addr_rom[17709]='h00000000;  wr_data_rom[17709]='h00000000;
    rd_cycle[17710] = 1'b0;  wr_cycle[17710] = 1'b0;  addr_rom[17710]='h00000000;  wr_data_rom[17710]='h00000000;
    rd_cycle[17711] = 1'b0;  wr_cycle[17711] = 1'b0;  addr_rom[17711]='h00000000;  wr_data_rom[17711]='h00000000;
    rd_cycle[17712] = 1'b0;  wr_cycle[17712] = 1'b0;  addr_rom[17712]='h00000000;  wr_data_rom[17712]='h00000000;
    rd_cycle[17713] = 1'b0;  wr_cycle[17713] = 1'b0;  addr_rom[17713]='h00000000;  wr_data_rom[17713]='h00000000;
    rd_cycle[17714] = 1'b0;  wr_cycle[17714] = 1'b0;  addr_rom[17714]='h00000000;  wr_data_rom[17714]='h00000000;
    rd_cycle[17715] = 1'b0;  wr_cycle[17715] = 1'b0;  addr_rom[17715]='h00000000;  wr_data_rom[17715]='h00000000;
    rd_cycle[17716] = 1'b0;  wr_cycle[17716] = 1'b0;  addr_rom[17716]='h00000000;  wr_data_rom[17716]='h00000000;
    rd_cycle[17717] = 1'b0;  wr_cycle[17717] = 1'b0;  addr_rom[17717]='h00000000;  wr_data_rom[17717]='h00000000;
    rd_cycle[17718] = 1'b0;  wr_cycle[17718] = 1'b0;  addr_rom[17718]='h00000000;  wr_data_rom[17718]='h00000000;
    rd_cycle[17719] = 1'b0;  wr_cycle[17719] = 1'b0;  addr_rom[17719]='h00000000;  wr_data_rom[17719]='h00000000;
    rd_cycle[17720] = 1'b0;  wr_cycle[17720] = 1'b0;  addr_rom[17720]='h00000000;  wr_data_rom[17720]='h00000000;
    rd_cycle[17721] = 1'b0;  wr_cycle[17721] = 1'b0;  addr_rom[17721]='h00000000;  wr_data_rom[17721]='h00000000;
    rd_cycle[17722] = 1'b0;  wr_cycle[17722] = 1'b0;  addr_rom[17722]='h00000000;  wr_data_rom[17722]='h00000000;
    rd_cycle[17723] = 1'b0;  wr_cycle[17723] = 1'b0;  addr_rom[17723]='h00000000;  wr_data_rom[17723]='h00000000;
    rd_cycle[17724] = 1'b0;  wr_cycle[17724] = 1'b0;  addr_rom[17724]='h00000000;  wr_data_rom[17724]='h00000000;
    rd_cycle[17725] = 1'b0;  wr_cycle[17725] = 1'b0;  addr_rom[17725]='h00000000;  wr_data_rom[17725]='h00000000;
    rd_cycle[17726] = 1'b0;  wr_cycle[17726] = 1'b0;  addr_rom[17726]='h00000000;  wr_data_rom[17726]='h00000000;
    rd_cycle[17727] = 1'b0;  wr_cycle[17727] = 1'b0;  addr_rom[17727]='h00000000;  wr_data_rom[17727]='h00000000;
    rd_cycle[17728] = 1'b0;  wr_cycle[17728] = 1'b0;  addr_rom[17728]='h00000000;  wr_data_rom[17728]='h00000000;
    rd_cycle[17729] = 1'b0;  wr_cycle[17729] = 1'b0;  addr_rom[17729]='h00000000;  wr_data_rom[17729]='h00000000;
    rd_cycle[17730] = 1'b0;  wr_cycle[17730] = 1'b0;  addr_rom[17730]='h00000000;  wr_data_rom[17730]='h00000000;
    rd_cycle[17731] = 1'b0;  wr_cycle[17731] = 1'b0;  addr_rom[17731]='h00000000;  wr_data_rom[17731]='h00000000;
    rd_cycle[17732] = 1'b0;  wr_cycle[17732] = 1'b0;  addr_rom[17732]='h00000000;  wr_data_rom[17732]='h00000000;
    rd_cycle[17733] = 1'b0;  wr_cycle[17733] = 1'b0;  addr_rom[17733]='h00000000;  wr_data_rom[17733]='h00000000;
    rd_cycle[17734] = 1'b0;  wr_cycle[17734] = 1'b0;  addr_rom[17734]='h00000000;  wr_data_rom[17734]='h00000000;
    rd_cycle[17735] = 1'b0;  wr_cycle[17735] = 1'b0;  addr_rom[17735]='h00000000;  wr_data_rom[17735]='h00000000;
    rd_cycle[17736] = 1'b0;  wr_cycle[17736] = 1'b0;  addr_rom[17736]='h00000000;  wr_data_rom[17736]='h00000000;
    rd_cycle[17737] = 1'b0;  wr_cycle[17737] = 1'b0;  addr_rom[17737]='h00000000;  wr_data_rom[17737]='h00000000;
    rd_cycle[17738] = 1'b0;  wr_cycle[17738] = 1'b0;  addr_rom[17738]='h00000000;  wr_data_rom[17738]='h00000000;
    rd_cycle[17739] = 1'b0;  wr_cycle[17739] = 1'b0;  addr_rom[17739]='h00000000;  wr_data_rom[17739]='h00000000;
    rd_cycle[17740] = 1'b0;  wr_cycle[17740] = 1'b0;  addr_rom[17740]='h00000000;  wr_data_rom[17740]='h00000000;
    rd_cycle[17741] = 1'b0;  wr_cycle[17741] = 1'b0;  addr_rom[17741]='h00000000;  wr_data_rom[17741]='h00000000;
    rd_cycle[17742] = 1'b0;  wr_cycle[17742] = 1'b0;  addr_rom[17742]='h00000000;  wr_data_rom[17742]='h00000000;
    rd_cycle[17743] = 1'b0;  wr_cycle[17743] = 1'b0;  addr_rom[17743]='h00000000;  wr_data_rom[17743]='h00000000;
    rd_cycle[17744] = 1'b0;  wr_cycle[17744] = 1'b0;  addr_rom[17744]='h00000000;  wr_data_rom[17744]='h00000000;
    rd_cycle[17745] = 1'b0;  wr_cycle[17745] = 1'b0;  addr_rom[17745]='h00000000;  wr_data_rom[17745]='h00000000;
    rd_cycle[17746] = 1'b0;  wr_cycle[17746] = 1'b0;  addr_rom[17746]='h00000000;  wr_data_rom[17746]='h00000000;
    rd_cycle[17747] = 1'b0;  wr_cycle[17747] = 1'b0;  addr_rom[17747]='h00000000;  wr_data_rom[17747]='h00000000;
    rd_cycle[17748] = 1'b0;  wr_cycle[17748] = 1'b0;  addr_rom[17748]='h00000000;  wr_data_rom[17748]='h00000000;
    rd_cycle[17749] = 1'b0;  wr_cycle[17749] = 1'b0;  addr_rom[17749]='h00000000;  wr_data_rom[17749]='h00000000;
    rd_cycle[17750] = 1'b0;  wr_cycle[17750] = 1'b0;  addr_rom[17750]='h00000000;  wr_data_rom[17750]='h00000000;
    rd_cycle[17751] = 1'b0;  wr_cycle[17751] = 1'b0;  addr_rom[17751]='h00000000;  wr_data_rom[17751]='h00000000;
    rd_cycle[17752] = 1'b0;  wr_cycle[17752] = 1'b0;  addr_rom[17752]='h00000000;  wr_data_rom[17752]='h00000000;
    rd_cycle[17753] = 1'b0;  wr_cycle[17753] = 1'b0;  addr_rom[17753]='h00000000;  wr_data_rom[17753]='h00000000;
    rd_cycle[17754] = 1'b0;  wr_cycle[17754] = 1'b0;  addr_rom[17754]='h00000000;  wr_data_rom[17754]='h00000000;
    rd_cycle[17755] = 1'b0;  wr_cycle[17755] = 1'b0;  addr_rom[17755]='h00000000;  wr_data_rom[17755]='h00000000;
    rd_cycle[17756] = 1'b0;  wr_cycle[17756] = 1'b0;  addr_rom[17756]='h00000000;  wr_data_rom[17756]='h00000000;
    rd_cycle[17757] = 1'b0;  wr_cycle[17757] = 1'b0;  addr_rom[17757]='h00000000;  wr_data_rom[17757]='h00000000;
    rd_cycle[17758] = 1'b0;  wr_cycle[17758] = 1'b0;  addr_rom[17758]='h00000000;  wr_data_rom[17758]='h00000000;
    rd_cycle[17759] = 1'b0;  wr_cycle[17759] = 1'b0;  addr_rom[17759]='h00000000;  wr_data_rom[17759]='h00000000;
    rd_cycle[17760] = 1'b0;  wr_cycle[17760] = 1'b0;  addr_rom[17760]='h00000000;  wr_data_rom[17760]='h00000000;
    rd_cycle[17761] = 1'b0;  wr_cycle[17761] = 1'b0;  addr_rom[17761]='h00000000;  wr_data_rom[17761]='h00000000;
    rd_cycle[17762] = 1'b0;  wr_cycle[17762] = 1'b0;  addr_rom[17762]='h00000000;  wr_data_rom[17762]='h00000000;
    rd_cycle[17763] = 1'b0;  wr_cycle[17763] = 1'b0;  addr_rom[17763]='h00000000;  wr_data_rom[17763]='h00000000;
    rd_cycle[17764] = 1'b0;  wr_cycle[17764] = 1'b0;  addr_rom[17764]='h00000000;  wr_data_rom[17764]='h00000000;
    rd_cycle[17765] = 1'b0;  wr_cycle[17765] = 1'b0;  addr_rom[17765]='h00000000;  wr_data_rom[17765]='h00000000;
    rd_cycle[17766] = 1'b0;  wr_cycle[17766] = 1'b0;  addr_rom[17766]='h00000000;  wr_data_rom[17766]='h00000000;
    rd_cycle[17767] = 1'b0;  wr_cycle[17767] = 1'b0;  addr_rom[17767]='h00000000;  wr_data_rom[17767]='h00000000;
    rd_cycle[17768] = 1'b0;  wr_cycle[17768] = 1'b0;  addr_rom[17768]='h00000000;  wr_data_rom[17768]='h00000000;
    rd_cycle[17769] = 1'b0;  wr_cycle[17769] = 1'b0;  addr_rom[17769]='h00000000;  wr_data_rom[17769]='h00000000;
    rd_cycle[17770] = 1'b0;  wr_cycle[17770] = 1'b0;  addr_rom[17770]='h00000000;  wr_data_rom[17770]='h00000000;
    rd_cycle[17771] = 1'b0;  wr_cycle[17771] = 1'b0;  addr_rom[17771]='h00000000;  wr_data_rom[17771]='h00000000;
    rd_cycle[17772] = 1'b0;  wr_cycle[17772] = 1'b0;  addr_rom[17772]='h00000000;  wr_data_rom[17772]='h00000000;
    rd_cycle[17773] = 1'b0;  wr_cycle[17773] = 1'b0;  addr_rom[17773]='h00000000;  wr_data_rom[17773]='h00000000;
    rd_cycle[17774] = 1'b0;  wr_cycle[17774] = 1'b0;  addr_rom[17774]='h00000000;  wr_data_rom[17774]='h00000000;
    rd_cycle[17775] = 1'b0;  wr_cycle[17775] = 1'b0;  addr_rom[17775]='h00000000;  wr_data_rom[17775]='h00000000;
    rd_cycle[17776] = 1'b0;  wr_cycle[17776] = 1'b0;  addr_rom[17776]='h00000000;  wr_data_rom[17776]='h00000000;
    rd_cycle[17777] = 1'b0;  wr_cycle[17777] = 1'b0;  addr_rom[17777]='h00000000;  wr_data_rom[17777]='h00000000;
    rd_cycle[17778] = 1'b0;  wr_cycle[17778] = 1'b0;  addr_rom[17778]='h00000000;  wr_data_rom[17778]='h00000000;
    rd_cycle[17779] = 1'b0;  wr_cycle[17779] = 1'b0;  addr_rom[17779]='h00000000;  wr_data_rom[17779]='h00000000;
    rd_cycle[17780] = 1'b0;  wr_cycle[17780] = 1'b0;  addr_rom[17780]='h00000000;  wr_data_rom[17780]='h00000000;
    rd_cycle[17781] = 1'b0;  wr_cycle[17781] = 1'b0;  addr_rom[17781]='h00000000;  wr_data_rom[17781]='h00000000;
    rd_cycle[17782] = 1'b0;  wr_cycle[17782] = 1'b0;  addr_rom[17782]='h00000000;  wr_data_rom[17782]='h00000000;
    rd_cycle[17783] = 1'b0;  wr_cycle[17783] = 1'b0;  addr_rom[17783]='h00000000;  wr_data_rom[17783]='h00000000;
    rd_cycle[17784] = 1'b0;  wr_cycle[17784] = 1'b0;  addr_rom[17784]='h00000000;  wr_data_rom[17784]='h00000000;
    rd_cycle[17785] = 1'b0;  wr_cycle[17785] = 1'b0;  addr_rom[17785]='h00000000;  wr_data_rom[17785]='h00000000;
    rd_cycle[17786] = 1'b0;  wr_cycle[17786] = 1'b0;  addr_rom[17786]='h00000000;  wr_data_rom[17786]='h00000000;
    rd_cycle[17787] = 1'b0;  wr_cycle[17787] = 1'b0;  addr_rom[17787]='h00000000;  wr_data_rom[17787]='h00000000;
    rd_cycle[17788] = 1'b0;  wr_cycle[17788] = 1'b0;  addr_rom[17788]='h00000000;  wr_data_rom[17788]='h00000000;
    rd_cycle[17789] = 1'b0;  wr_cycle[17789] = 1'b0;  addr_rom[17789]='h00000000;  wr_data_rom[17789]='h00000000;
    rd_cycle[17790] = 1'b0;  wr_cycle[17790] = 1'b0;  addr_rom[17790]='h00000000;  wr_data_rom[17790]='h00000000;
    rd_cycle[17791] = 1'b0;  wr_cycle[17791] = 1'b0;  addr_rom[17791]='h00000000;  wr_data_rom[17791]='h00000000;
    rd_cycle[17792] = 1'b0;  wr_cycle[17792] = 1'b0;  addr_rom[17792]='h00000000;  wr_data_rom[17792]='h00000000;
    rd_cycle[17793] = 1'b0;  wr_cycle[17793] = 1'b0;  addr_rom[17793]='h00000000;  wr_data_rom[17793]='h00000000;
    rd_cycle[17794] = 1'b0;  wr_cycle[17794] = 1'b0;  addr_rom[17794]='h00000000;  wr_data_rom[17794]='h00000000;
    rd_cycle[17795] = 1'b0;  wr_cycle[17795] = 1'b0;  addr_rom[17795]='h00000000;  wr_data_rom[17795]='h00000000;
    rd_cycle[17796] = 1'b0;  wr_cycle[17796] = 1'b0;  addr_rom[17796]='h00000000;  wr_data_rom[17796]='h00000000;
    rd_cycle[17797] = 1'b0;  wr_cycle[17797] = 1'b0;  addr_rom[17797]='h00000000;  wr_data_rom[17797]='h00000000;
    rd_cycle[17798] = 1'b0;  wr_cycle[17798] = 1'b0;  addr_rom[17798]='h00000000;  wr_data_rom[17798]='h00000000;
    rd_cycle[17799] = 1'b0;  wr_cycle[17799] = 1'b0;  addr_rom[17799]='h00000000;  wr_data_rom[17799]='h00000000;
    rd_cycle[17800] = 1'b0;  wr_cycle[17800] = 1'b0;  addr_rom[17800]='h00000000;  wr_data_rom[17800]='h00000000;
    rd_cycle[17801] = 1'b0;  wr_cycle[17801] = 1'b0;  addr_rom[17801]='h00000000;  wr_data_rom[17801]='h00000000;
    rd_cycle[17802] = 1'b0;  wr_cycle[17802] = 1'b0;  addr_rom[17802]='h00000000;  wr_data_rom[17802]='h00000000;
    rd_cycle[17803] = 1'b0;  wr_cycle[17803] = 1'b0;  addr_rom[17803]='h00000000;  wr_data_rom[17803]='h00000000;
    rd_cycle[17804] = 1'b0;  wr_cycle[17804] = 1'b0;  addr_rom[17804]='h00000000;  wr_data_rom[17804]='h00000000;
    rd_cycle[17805] = 1'b0;  wr_cycle[17805] = 1'b0;  addr_rom[17805]='h00000000;  wr_data_rom[17805]='h00000000;
    rd_cycle[17806] = 1'b0;  wr_cycle[17806] = 1'b0;  addr_rom[17806]='h00000000;  wr_data_rom[17806]='h00000000;
    rd_cycle[17807] = 1'b0;  wr_cycle[17807] = 1'b0;  addr_rom[17807]='h00000000;  wr_data_rom[17807]='h00000000;
    rd_cycle[17808] = 1'b0;  wr_cycle[17808] = 1'b0;  addr_rom[17808]='h00000000;  wr_data_rom[17808]='h00000000;
    rd_cycle[17809] = 1'b0;  wr_cycle[17809] = 1'b0;  addr_rom[17809]='h00000000;  wr_data_rom[17809]='h00000000;
    rd_cycle[17810] = 1'b0;  wr_cycle[17810] = 1'b0;  addr_rom[17810]='h00000000;  wr_data_rom[17810]='h00000000;
    rd_cycle[17811] = 1'b0;  wr_cycle[17811] = 1'b0;  addr_rom[17811]='h00000000;  wr_data_rom[17811]='h00000000;
    rd_cycle[17812] = 1'b0;  wr_cycle[17812] = 1'b0;  addr_rom[17812]='h00000000;  wr_data_rom[17812]='h00000000;
    rd_cycle[17813] = 1'b0;  wr_cycle[17813] = 1'b0;  addr_rom[17813]='h00000000;  wr_data_rom[17813]='h00000000;
    rd_cycle[17814] = 1'b0;  wr_cycle[17814] = 1'b0;  addr_rom[17814]='h00000000;  wr_data_rom[17814]='h00000000;
    rd_cycle[17815] = 1'b0;  wr_cycle[17815] = 1'b0;  addr_rom[17815]='h00000000;  wr_data_rom[17815]='h00000000;
    rd_cycle[17816] = 1'b0;  wr_cycle[17816] = 1'b0;  addr_rom[17816]='h00000000;  wr_data_rom[17816]='h00000000;
    rd_cycle[17817] = 1'b0;  wr_cycle[17817] = 1'b0;  addr_rom[17817]='h00000000;  wr_data_rom[17817]='h00000000;
    rd_cycle[17818] = 1'b0;  wr_cycle[17818] = 1'b0;  addr_rom[17818]='h00000000;  wr_data_rom[17818]='h00000000;
    rd_cycle[17819] = 1'b0;  wr_cycle[17819] = 1'b0;  addr_rom[17819]='h00000000;  wr_data_rom[17819]='h00000000;
    rd_cycle[17820] = 1'b0;  wr_cycle[17820] = 1'b0;  addr_rom[17820]='h00000000;  wr_data_rom[17820]='h00000000;
    rd_cycle[17821] = 1'b0;  wr_cycle[17821] = 1'b0;  addr_rom[17821]='h00000000;  wr_data_rom[17821]='h00000000;
    rd_cycle[17822] = 1'b0;  wr_cycle[17822] = 1'b0;  addr_rom[17822]='h00000000;  wr_data_rom[17822]='h00000000;
    rd_cycle[17823] = 1'b0;  wr_cycle[17823] = 1'b0;  addr_rom[17823]='h00000000;  wr_data_rom[17823]='h00000000;
    rd_cycle[17824] = 1'b0;  wr_cycle[17824] = 1'b0;  addr_rom[17824]='h00000000;  wr_data_rom[17824]='h00000000;
    rd_cycle[17825] = 1'b0;  wr_cycle[17825] = 1'b0;  addr_rom[17825]='h00000000;  wr_data_rom[17825]='h00000000;
    rd_cycle[17826] = 1'b0;  wr_cycle[17826] = 1'b0;  addr_rom[17826]='h00000000;  wr_data_rom[17826]='h00000000;
    rd_cycle[17827] = 1'b0;  wr_cycle[17827] = 1'b0;  addr_rom[17827]='h00000000;  wr_data_rom[17827]='h00000000;
    rd_cycle[17828] = 1'b0;  wr_cycle[17828] = 1'b0;  addr_rom[17828]='h00000000;  wr_data_rom[17828]='h00000000;
    rd_cycle[17829] = 1'b0;  wr_cycle[17829] = 1'b0;  addr_rom[17829]='h00000000;  wr_data_rom[17829]='h00000000;
    rd_cycle[17830] = 1'b0;  wr_cycle[17830] = 1'b0;  addr_rom[17830]='h00000000;  wr_data_rom[17830]='h00000000;
    rd_cycle[17831] = 1'b0;  wr_cycle[17831] = 1'b0;  addr_rom[17831]='h00000000;  wr_data_rom[17831]='h00000000;
    rd_cycle[17832] = 1'b0;  wr_cycle[17832] = 1'b0;  addr_rom[17832]='h00000000;  wr_data_rom[17832]='h00000000;
    rd_cycle[17833] = 1'b0;  wr_cycle[17833] = 1'b0;  addr_rom[17833]='h00000000;  wr_data_rom[17833]='h00000000;
    rd_cycle[17834] = 1'b0;  wr_cycle[17834] = 1'b0;  addr_rom[17834]='h00000000;  wr_data_rom[17834]='h00000000;
    rd_cycle[17835] = 1'b0;  wr_cycle[17835] = 1'b0;  addr_rom[17835]='h00000000;  wr_data_rom[17835]='h00000000;
    rd_cycle[17836] = 1'b0;  wr_cycle[17836] = 1'b0;  addr_rom[17836]='h00000000;  wr_data_rom[17836]='h00000000;
    rd_cycle[17837] = 1'b0;  wr_cycle[17837] = 1'b0;  addr_rom[17837]='h00000000;  wr_data_rom[17837]='h00000000;
    rd_cycle[17838] = 1'b0;  wr_cycle[17838] = 1'b0;  addr_rom[17838]='h00000000;  wr_data_rom[17838]='h00000000;
    rd_cycle[17839] = 1'b0;  wr_cycle[17839] = 1'b0;  addr_rom[17839]='h00000000;  wr_data_rom[17839]='h00000000;
    rd_cycle[17840] = 1'b0;  wr_cycle[17840] = 1'b0;  addr_rom[17840]='h00000000;  wr_data_rom[17840]='h00000000;
    rd_cycle[17841] = 1'b0;  wr_cycle[17841] = 1'b0;  addr_rom[17841]='h00000000;  wr_data_rom[17841]='h00000000;
    rd_cycle[17842] = 1'b0;  wr_cycle[17842] = 1'b0;  addr_rom[17842]='h00000000;  wr_data_rom[17842]='h00000000;
    rd_cycle[17843] = 1'b0;  wr_cycle[17843] = 1'b0;  addr_rom[17843]='h00000000;  wr_data_rom[17843]='h00000000;
    rd_cycle[17844] = 1'b0;  wr_cycle[17844] = 1'b0;  addr_rom[17844]='h00000000;  wr_data_rom[17844]='h00000000;
    rd_cycle[17845] = 1'b0;  wr_cycle[17845] = 1'b0;  addr_rom[17845]='h00000000;  wr_data_rom[17845]='h00000000;
    rd_cycle[17846] = 1'b0;  wr_cycle[17846] = 1'b0;  addr_rom[17846]='h00000000;  wr_data_rom[17846]='h00000000;
    rd_cycle[17847] = 1'b0;  wr_cycle[17847] = 1'b0;  addr_rom[17847]='h00000000;  wr_data_rom[17847]='h00000000;
    rd_cycle[17848] = 1'b0;  wr_cycle[17848] = 1'b0;  addr_rom[17848]='h00000000;  wr_data_rom[17848]='h00000000;
    rd_cycle[17849] = 1'b0;  wr_cycle[17849] = 1'b0;  addr_rom[17849]='h00000000;  wr_data_rom[17849]='h00000000;
    rd_cycle[17850] = 1'b0;  wr_cycle[17850] = 1'b0;  addr_rom[17850]='h00000000;  wr_data_rom[17850]='h00000000;
    rd_cycle[17851] = 1'b0;  wr_cycle[17851] = 1'b0;  addr_rom[17851]='h00000000;  wr_data_rom[17851]='h00000000;
    rd_cycle[17852] = 1'b0;  wr_cycle[17852] = 1'b0;  addr_rom[17852]='h00000000;  wr_data_rom[17852]='h00000000;
    rd_cycle[17853] = 1'b0;  wr_cycle[17853] = 1'b0;  addr_rom[17853]='h00000000;  wr_data_rom[17853]='h00000000;
    rd_cycle[17854] = 1'b0;  wr_cycle[17854] = 1'b0;  addr_rom[17854]='h00000000;  wr_data_rom[17854]='h00000000;
    rd_cycle[17855] = 1'b0;  wr_cycle[17855] = 1'b0;  addr_rom[17855]='h00000000;  wr_data_rom[17855]='h00000000;
    rd_cycle[17856] = 1'b0;  wr_cycle[17856] = 1'b0;  addr_rom[17856]='h00000000;  wr_data_rom[17856]='h00000000;
    rd_cycle[17857] = 1'b0;  wr_cycle[17857] = 1'b0;  addr_rom[17857]='h00000000;  wr_data_rom[17857]='h00000000;
    rd_cycle[17858] = 1'b0;  wr_cycle[17858] = 1'b0;  addr_rom[17858]='h00000000;  wr_data_rom[17858]='h00000000;
    rd_cycle[17859] = 1'b0;  wr_cycle[17859] = 1'b0;  addr_rom[17859]='h00000000;  wr_data_rom[17859]='h00000000;
    rd_cycle[17860] = 1'b0;  wr_cycle[17860] = 1'b0;  addr_rom[17860]='h00000000;  wr_data_rom[17860]='h00000000;
    rd_cycle[17861] = 1'b0;  wr_cycle[17861] = 1'b0;  addr_rom[17861]='h00000000;  wr_data_rom[17861]='h00000000;
    rd_cycle[17862] = 1'b0;  wr_cycle[17862] = 1'b0;  addr_rom[17862]='h00000000;  wr_data_rom[17862]='h00000000;
    rd_cycle[17863] = 1'b0;  wr_cycle[17863] = 1'b0;  addr_rom[17863]='h00000000;  wr_data_rom[17863]='h00000000;
    rd_cycle[17864] = 1'b0;  wr_cycle[17864] = 1'b0;  addr_rom[17864]='h00000000;  wr_data_rom[17864]='h00000000;
    rd_cycle[17865] = 1'b0;  wr_cycle[17865] = 1'b0;  addr_rom[17865]='h00000000;  wr_data_rom[17865]='h00000000;
    rd_cycle[17866] = 1'b0;  wr_cycle[17866] = 1'b0;  addr_rom[17866]='h00000000;  wr_data_rom[17866]='h00000000;
    rd_cycle[17867] = 1'b0;  wr_cycle[17867] = 1'b0;  addr_rom[17867]='h00000000;  wr_data_rom[17867]='h00000000;
    rd_cycle[17868] = 1'b0;  wr_cycle[17868] = 1'b0;  addr_rom[17868]='h00000000;  wr_data_rom[17868]='h00000000;
    rd_cycle[17869] = 1'b0;  wr_cycle[17869] = 1'b0;  addr_rom[17869]='h00000000;  wr_data_rom[17869]='h00000000;
    rd_cycle[17870] = 1'b0;  wr_cycle[17870] = 1'b0;  addr_rom[17870]='h00000000;  wr_data_rom[17870]='h00000000;
    rd_cycle[17871] = 1'b0;  wr_cycle[17871] = 1'b0;  addr_rom[17871]='h00000000;  wr_data_rom[17871]='h00000000;
    rd_cycle[17872] = 1'b0;  wr_cycle[17872] = 1'b0;  addr_rom[17872]='h00000000;  wr_data_rom[17872]='h00000000;
    rd_cycle[17873] = 1'b0;  wr_cycle[17873] = 1'b0;  addr_rom[17873]='h00000000;  wr_data_rom[17873]='h00000000;
    rd_cycle[17874] = 1'b0;  wr_cycle[17874] = 1'b0;  addr_rom[17874]='h00000000;  wr_data_rom[17874]='h00000000;
    rd_cycle[17875] = 1'b0;  wr_cycle[17875] = 1'b0;  addr_rom[17875]='h00000000;  wr_data_rom[17875]='h00000000;
    rd_cycle[17876] = 1'b0;  wr_cycle[17876] = 1'b0;  addr_rom[17876]='h00000000;  wr_data_rom[17876]='h00000000;
    rd_cycle[17877] = 1'b0;  wr_cycle[17877] = 1'b0;  addr_rom[17877]='h00000000;  wr_data_rom[17877]='h00000000;
    rd_cycle[17878] = 1'b0;  wr_cycle[17878] = 1'b0;  addr_rom[17878]='h00000000;  wr_data_rom[17878]='h00000000;
    rd_cycle[17879] = 1'b0;  wr_cycle[17879] = 1'b0;  addr_rom[17879]='h00000000;  wr_data_rom[17879]='h00000000;
    rd_cycle[17880] = 1'b0;  wr_cycle[17880] = 1'b0;  addr_rom[17880]='h00000000;  wr_data_rom[17880]='h00000000;
    rd_cycle[17881] = 1'b0;  wr_cycle[17881] = 1'b0;  addr_rom[17881]='h00000000;  wr_data_rom[17881]='h00000000;
    rd_cycle[17882] = 1'b0;  wr_cycle[17882] = 1'b0;  addr_rom[17882]='h00000000;  wr_data_rom[17882]='h00000000;
    rd_cycle[17883] = 1'b0;  wr_cycle[17883] = 1'b0;  addr_rom[17883]='h00000000;  wr_data_rom[17883]='h00000000;
    rd_cycle[17884] = 1'b0;  wr_cycle[17884] = 1'b0;  addr_rom[17884]='h00000000;  wr_data_rom[17884]='h00000000;
    rd_cycle[17885] = 1'b0;  wr_cycle[17885] = 1'b0;  addr_rom[17885]='h00000000;  wr_data_rom[17885]='h00000000;
    rd_cycle[17886] = 1'b0;  wr_cycle[17886] = 1'b0;  addr_rom[17886]='h00000000;  wr_data_rom[17886]='h00000000;
    rd_cycle[17887] = 1'b0;  wr_cycle[17887] = 1'b0;  addr_rom[17887]='h00000000;  wr_data_rom[17887]='h00000000;
    rd_cycle[17888] = 1'b0;  wr_cycle[17888] = 1'b0;  addr_rom[17888]='h00000000;  wr_data_rom[17888]='h00000000;
    rd_cycle[17889] = 1'b0;  wr_cycle[17889] = 1'b0;  addr_rom[17889]='h00000000;  wr_data_rom[17889]='h00000000;
    rd_cycle[17890] = 1'b0;  wr_cycle[17890] = 1'b0;  addr_rom[17890]='h00000000;  wr_data_rom[17890]='h00000000;
    rd_cycle[17891] = 1'b0;  wr_cycle[17891] = 1'b0;  addr_rom[17891]='h00000000;  wr_data_rom[17891]='h00000000;
    rd_cycle[17892] = 1'b0;  wr_cycle[17892] = 1'b0;  addr_rom[17892]='h00000000;  wr_data_rom[17892]='h00000000;
    rd_cycle[17893] = 1'b0;  wr_cycle[17893] = 1'b0;  addr_rom[17893]='h00000000;  wr_data_rom[17893]='h00000000;
    rd_cycle[17894] = 1'b0;  wr_cycle[17894] = 1'b0;  addr_rom[17894]='h00000000;  wr_data_rom[17894]='h00000000;
    rd_cycle[17895] = 1'b0;  wr_cycle[17895] = 1'b0;  addr_rom[17895]='h00000000;  wr_data_rom[17895]='h00000000;
    rd_cycle[17896] = 1'b0;  wr_cycle[17896] = 1'b0;  addr_rom[17896]='h00000000;  wr_data_rom[17896]='h00000000;
    rd_cycle[17897] = 1'b0;  wr_cycle[17897] = 1'b0;  addr_rom[17897]='h00000000;  wr_data_rom[17897]='h00000000;
    rd_cycle[17898] = 1'b0;  wr_cycle[17898] = 1'b0;  addr_rom[17898]='h00000000;  wr_data_rom[17898]='h00000000;
    rd_cycle[17899] = 1'b0;  wr_cycle[17899] = 1'b0;  addr_rom[17899]='h00000000;  wr_data_rom[17899]='h00000000;
    rd_cycle[17900] = 1'b0;  wr_cycle[17900] = 1'b0;  addr_rom[17900]='h00000000;  wr_data_rom[17900]='h00000000;
    rd_cycle[17901] = 1'b0;  wr_cycle[17901] = 1'b0;  addr_rom[17901]='h00000000;  wr_data_rom[17901]='h00000000;
    rd_cycle[17902] = 1'b0;  wr_cycle[17902] = 1'b0;  addr_rom[17902]='h00000000;  wr_data_rom[17902]='h00000000;
    rd_cycle[17903] = 1'b0;  wr_cycle[17903] = 1'b0;  addr_rom[17903]='h00000000;  wr_data_rom[17903]='h00000000;
    rd_cycle[17904] = 1'b0;  wr_cycle[17904] = 1'b0;  addr_rom[17904]='h00000000;  wr_data_rom[17904]='h00000000;
    rd_cycle[17905] = 1'b0;  wr_cycle[17905] = 1'b0;  addr_rom[17905]='h00000000;  wr_data_rom[17905]='h00000000;
    rd_cycle[17906] = 1'b0;  wr_cycle[17906] = 1'b0;  addr_rom[17906]='h00000000;  wr_data_rom[17906]='h00000000;
    rd_cycle[17907] = 1'b0;  wr_cycle[17907] = 1'b0;  addr_rom[17907]='h00000000;  wr_data_rom[17907]='h00000000;
    rd_cycle[17908] = 1'b0;  wr_cycle[17908] = 1'b0;  addr_rom[17908]='h00000000;  wr_data_rom[17908]='h00000000;
    rd_cycle[17909] = 1'b0;  wr_cycle[17909] = 1'b0;  addr_rom[17909]='h00000000;  wr_data_rom[17909]='h00000000;
    rd_cycle[17910] = 1'b0;  wr_cycle[17910] = 1'b0;  addr_rom[17910]='h00000000;  wr_data_rom[17910]='h00000000;
    rd_cycle[17911] = 1'b0;  wr_cycle[17911] = 1'b0;  addr_rom[17911]='h00000000;  wr_data_rom[17911]='h00000000;
    rd_cycle[17912] = 1'b0;  wr_cycle[17912] = 1'b0;  addr_rom[17912]='h00000000;  wr_data_rom[17912]='h00000000;
    rd_cycle[17913] = 1'b0;  wr_cycle[17913] = 1'b0;  addr_rom[17913]='h00000000;  wr_data_rom[17913]='h00000000;
    rd_cycle[17914] = 1'b0;  wr_cycle[17914] = 1'b0;  addr_rom[17914]='h00000000;  wr_data_rom[17914]='h00000000;
    rd_cycle[17915] = 1'b0;  wr_cycle[17915] = 1'b0;  addr_rom[17915]='h00000000;  wr_data_rom[17915]='h00000000;
    rd_cycle[17916] = 1'b0;  wr_cycle[17916] = 1'b0;  addr_rom[17916]='h00000000;  wr_data_rom[17916]='h00000000;
    rd_cycle[17917] = 1'b0;  wr_cycle[17917] = 1'b0;  addr_rom[17917]='h00000000;  wr_data_rom[17917]='h00000000;
    rd_cycle[17918] = 1'b0;  wr_cycle[17918] = 1'b0;  addr_rom[17918]='h00000000;  wr_data_rom[17918]='h00000000;
    rd_cycle[17919] = 1'b0;  wr_cycle[17919] = 1'b0;  addr_rom[17919]='h00000000;  wr_data_rom[17919]='h00000000;
    rd_cycle[17920] = 1'b0;  wr_cycle[17920] = 1'b0;  addr_rom[17920]='h00000000;  wr_data_rom[17920]='h00000000;
    rd_cycle[17921] = 1'b0;  wr_cycle[17921] = 1'b0;  addr_rom[17921]='h00000000;  wr_data_rom[17921]='h00000000;
    rd_cycle[17922] = 1'b0;  wr_cycle[17922] = 1'b0;  addr_rom[17922]='h00000000;  wr_data_rom[17922]='h00000000;
    rd_cycle[17923] = 1'b0;  wr_cycle[17923] = 1'b0;  addr_rom[17923]='h00000000;  wr_data_rom[17923]='h00000000;
    rd_cycle[17924] = 1'b0;  wr_cycle[17924] = 1'b0;  addr_rom[17924]='h00000000;  wr_data_rom[17924]='h00000000;
    rd_cycle[17925] = 1'b0;  wr_cycle[17925] = 1'b0;  addr_rom[17925]='h00000000;  wr_data_rom[17925]='h00000000;
    rd_cycle[17926] = 1'b0;  wr_cycle[17926] = 1'b0;  addr_rom[17926]='h00000000;  wr_data_rom[17926]='h00000000;
    rd_cycle[17927] = 1'b0;  wr_cycle[17927] = 1'b0;  addr_rom[17927]='h00000000;  wr_data_rom[17927]='h00000000;
    rd_cycle[17928] = 1'b0;  wr_cycle[17928] = 1'b0;  addr_rom[17928]='h00000000;  wr_data_rom[17928]='h00000000;
    rd_cycle[17929] = 1'b0;  wr_cycle[17929] = 1'b0;  addr_rom[17929]='h00000000;  wr_data_rom[17929]='h00000000;
    rd_cycle[17930] = 1'b0;  wr_cycle[17930] = 1'b0;  addr_rom[17930]='h00000000;  wr_data_rom[17930]='h00000000;
    rd_cycle[17931] = 1'b0;  wr_cycle[17931] = 1'b0;  addr_rom[17931]='h00000000;  wr_data_rom[17931]='h00000000;
    rd_cycle[17932] = 1'b0;  wr_cycle[17932] = 1'b0;  addr_rom[17932]='h00000000;  wr_data_rom[17932]='h00000000;
    rd_cycle[17933] = 1'b0;  wr_cycle[17933] = 1'b0;  addr_rom[17933]='h00000000;  wr_data_rom[17933]='h00000000;
    rd_cycle[17934] = 1'b0;  wr_cycle[17934] = 1'b0;  addr_rom[17934]='h00000000;  wr_data_rom[17934]='h00000000;
    rd_cycle[17935] = 1'b0;  wr_cycle[17935] = 1'b0;  addr_rom[17935]='h00000000;  wr_data_rom[17935]='h00000000;
    rd_cycle[17936] = 1'b0;  wr_cycle[17936] = 1'b0;  addr_rom[17936]='h00000000;  wr_data_rom[17936]='h00000000;
    rd_cycle[17937] = 1'b0;  wr_cycle[17937] = 1'b0;  addr_rom[17937]='h00000000;  wr_data_rom[17937]='h00000000;
    rd_cycle[17938] = 1'b0;  wr_cycle[17938] = 1'b0;  addr_rom[17938]='h00000000;  wr_data_rom[17938]='h00000000;
    rd_cycle[17939] = 1'b0;  wr_cycle[17939] = 1'b0;  addr_rom[17939]='h00000000;  wr_data_rom[17939]='h00000000;
    rd_cycle[17940] = 1'b0;  wr_cycle[17940] = 1'b0;  addr_rom[17940]='h00000000;  wr_data_rom[17940]='h00000000;
    rd_cycle[17941] = 1'b0;  wr_cycle[17941] = 1'b0;  addr_rom[17941]='h00000000;  wr_data_rom[17941]='h00000000;
    rd_cycle[17942] = 1'b0;  wr_cycle[17942] = 1'b0;  addr_rom[17942]='h00000000;  wr_data_rom[17942]='h00000000;
    rd_cycle[17943] = 1'b0;  wr_cycle[17943] = 1'b0;  addr_rom[17943]='h00000000;  wr_data_rom[17943]='h00000000;
    rd_cycle[17944] = 1'b0;  wr_cycle[17944] = 1'b0;  addr_rom[17944]='h00000000;  wr_data_rom[17944]='h00000000;
    rd_cycle[17945] = 1'b0;  wr_cycle[17945] = 1'b0;  addr_rom[17945]='h00000000;  wr_data_rom[17945]='h00000000;
    rd_cycle[17946] = 1'b0;  wr_cycle[17946] = 1'b0;  addr_rom[17946]='h00000000;  wr_data_rom[17946]='h00000000;
    rd_cycle[17947] = 1'b0;  wr_cycle[17947] = 1'b0;  addr_rom[17947]='h00000000;  wr_data_rom[17947]='h00000000;
    rd_cycle[17948] = 1'b0;  wr_cycle[17948] = 1'b0;  addr_rom[17948]='h00000000;  wr_data_rom[17948]='h00000000;
    rd_cycle[17949] = 1'b0;  wr_cycle[17949] = 1'b0;  addr_rom[17949]='h00000000;  wr_data_rom[17949]='h00000000;
    rd_cycle[17950] = 1'b0;  wr_cycle[17950] = 1'b0;  addr_rom[17950]='h00000000;  wr_data_rom[17950]='h00000000;
    rd_cycle[17951] = 1'b0;  wr_cycle[17951] = 1'b0;  addr_rom[17951]='h00000000;  wr_data_rom[17951]='h00000000;
    rd_cycle[17952] = 1'b0;  wr_cycle[17952] = 1'b0;  addr_rom[17952]='h00000000;  wr_data_rom[17952]='h00000000;
    rd_cycle[17953] = 1'b0;  wr_cycle[17953] = 1'b0;  addr_rom[17953]='h00000000;  wr_data_rom[17953]='h00000000;
    rd_cycle[17954] = 1'b0;  wr_cycle[17954] = 1'b0;  addr_rom[17954]='h00000000;  wr_data_rom[17954]='h00000000;
    rd_cycle[17955] = 1'b0;  wr_cycle[17955] = 1'b0;  addr_rom[17955]='h00000000;  wr_data_rom[17955]='h00000000;
    rd_cycle[17956] = 1'b0;  wr_cycle[17956] = 1'b0;  addr_rom[17956]='h00000000;  wr_data_rom[17956]='h00000000;
    rd_cycle[17957] = 1'b0;  wr_cycle[17957] = 1'b0;  addr_rom[17957]='h00000000;  wr_data_rom[17957]='h00000000;
    rd_cycle[17958] = 1'b0;  wr_cycle[17958] = 1'b0;  addr_rom[17958]='h00000000;  wr_data_rom[17958]='h00000000;
    rd_cycle[17959] = 1'b0;  wr_cycle[17959] = 1'b0;  addr_rom[17959]='h00000000;  wr_data_rom[17959]='h00000000;
    rd_cycle[17960] = 1'b0;  wr_cycle[17960] = 1'b0;  addr_rom[17960]='h00000000;  wr_data_rom[17960]='h00000000;
    rd_cycle[17961] = 1'b0;  wr_cycle[17961] = 1'b0;  addr_rom[17961]='h00000000;  wr_data_rom[17961]='h00000000;
    rd_cycle[17962] = 1'b0;  wr_cycle[17962] = 1'b0;  addr_rom[17962]='h00000000;  wr_data_rom[17962]='h00000000;
    rd_cycle[17963] = 1'b0;  wr_cycle[17963] = 1'b0;  addr_rom[17963]='h00000000;  wr_data_rom[17963]='h00000000;
    rd_cycle[17964] = 1'b0;  wr_cycle[17964] = 1'b0;  addr_rom[17964]='h00000000;  wr_data_rom[17964]='h00000000;
    rd_cycle[17965] = 1'b0;  wr_cycle[17965] = 1'b0;  addr_rom[17965]='h00000000;  wr_data_rom[17965]='h00000000;
    rd_cycle[17966] = 1'b0;  wr_cycle[17966] = 1'b0;  addr_rom[17966]='h00000000;  wr_data_rom[17966]='h00000000;
    rd_cycle[17967] = 1'b0;  wr_cycle[17967] = 1'b0;  addr_rom[17967]='h00000000;  wr_data_rom[17967]='h00000000;
    rd_cycle[17968] = 1'b0;  wr_cycle[17968] = 1'b0;  addr_rom[17968]='h00000000;  wr_data_rom[17968]='h00000000;
    rd_cycle[17969] = 1'b0;  wr_cycle[17969] = 1'b0;  addr_rom[17969]='h00000000;  wr_data_rom[17969]='h00000000;
    rd_cycle[17970] = 1'b0;  wr_cycle[17970] = 1'b0;  addr_rom[17970]='h00000000;  wr_data_rom[17970]='h00000000;
    rd_cycle[17971] = 1'b0;  wr_cycle[17971] = 1'b0;  addr_rom[17971]='h00000000;  wr_data_rom[17971]='h00000000;
    rd_cycle[17972] = 1'b0;  wr_cycle[17972] = 1'b0;  addr_rom[17972]='h00000000;  wr_data_rom[17972]='h00000000;
    rd_cycle[17973] = 1'b0;  wr_cycle[17973] = 1'b0;  addr_rom[17973]='h00000000;  wr_data_rom[17973]='h00000000;
    rd_cycle[17974] = 1'b0;  wr_cycle[17974] = 1'b0;  addr_rom[17974]='h00000000;  wr_data_rom[17974]='h00000000;
    rd_cycle[17975] = 1'b0;  wr_cycle[17975] = 1'b0;  addr_rom[17975]='h00000000;  wr_data_rom[17975]='h00000000;
    rd_cycle[17976] = 1'b0;  wr_cycle[17976] = 1'b0;  addr_rom[17976]='h00000000;  wr_data_rom[17976]='h00000000;
    rd_cycle[17977] = 1'b0;  wr_cycle[17977] = 1'b0;  addr_rom[17977]='h00000000;  wr_data_rom[17977]='h00000000;
    rd_cycle[17978] = 1'b0;  wr_cycle[17978] = 1'b0;  addr_rom[17978]='h00000000;  wr_data_rom[17978]='h00000000;
    rd_cycle[17979] = 1'b0;  wr_cycle[17979] = 1'b0;  addr_rom[17979]='h00000000;  wr_data_rom[17979]='h00000000;
    rd_cycle[17980] = 1'b0;  wr_cycle[17980] = 1'b0;  addr_rom[17980]='h00000000;  wr_data_rom[17980]='h00000000;
    rd_cycle[17981] = 1'b0;  wr_cycle[17981] = 1'b0;  addr_rom[17981]='h00000000;  wr_data_rom[17981]='h00000000;
    rd_cycle[17982] = 1'b0;  wr_cycle[17982] = 1'b0;  addr_rom[17982]='h00000000;  wr_data_rom[17982]='h00000000;
    rd_cycle[17983] = 1'b0;  wr_cycle[17983] = 1'b0;  addr_rom[17983]='h00000000;  wr_data_rom[17983]='h00000000;
    rd_cycle[17984] = 1'b0;  wr_cycle[17984] = 1'b0;  addr_rom[17984]='h00000000;  wr_data_rom[17984]='h00000000;
    rd_cycle[17985] = 1'b0;  wr_cycle[17985] = 1'b0;  addr_rom[17985]='h00000000;  wr_data_rom[17985]='h00000000;
    rd_cycle[17986] = 1'b0;  wr_cycle[17986] = 1'b0;  addr_rom[17986]='h00000000;  wr_data_rom[17986]='h00000000;
    rd_cycle[17987] = 1'b0;  wr_cycle[17987] = 1'b0;  addr_rom[17987]='h00000000;  wr_data_rom[17987]='h00000000;
    rd_cycle[17988] = 1'b0;  wr_cycle[17988] = 1'b0;  addr_rom[17988]='h00000000;  wr_data_rom[17988]='h00000000;
    rd_cycle[17989] = 1'b0;  wr_cycle[17989] = 1'b0;  addr_rom[17989]='h00000000;  wr_data_rom[17989]='h00000000;
    rd_cycle[17990] = 1'b0;  wr_cycle[17990] = 1'b0;  addr_rom[17990]='h00000000;  wr_data_rom[17990]='h00000000;
    rd_cycle[17991] = 1'b0;  wr_cycle[17991] = 1'b0;  addr_rom[17991]='h00000000;  wr_data_rom[17991]='h00000000;
    rd_cycle[17992] = 1'b0;  wr_cycle[17992] = 1'b0;  addr_rom[17992]='h00000000;  wr_data_rom[17992]='h00000000;
    rd_cycle[17993] = 1'b0;  wr_cycle[17993] = 1'b0;  addr_rom[17993]='h00000000;  wr_data_rom[17993]='h00000000;
    rd_cycle[17994] = 1'b0;  wr_cycle[17994] = 1'b0;  addr_rom[17994]='h00000000;  wr_data_rom[17994]='h00000000;
    rd_cycle[17995] = 1'b0;  wr_cycle[17995] = 1'b0;  addr_rom[17995]='h00000000;  wr_data_rom[17995]='h00000000;
    rd_cycle[17996] = 1'b0;  wr_cycle[17996] = 1'b0;  addr_rom[17996]='h00000000;  wr_data_rom[17996]='h00000000;
    rd_cycle[17997] = 1'b0;  wr_cycle[17997] = 1'b0;  addr_rom[17997]='h00000000;  wr_data_rom[17997]='h00000000;
    rd_cycle[17998] = 1'b0;  wr_cycle[17998] = 1'b0;  addr_rom[17998]='h00000000;  wr_data_rom[17998]='h00000000;
    rd_cycle[17999] = 1'b0;  wr_cycle[17999] = 1'b0;  addr_rom[17999]='h00000000;  wr_data_rom[17999]='h00000000;
    rd_cycle[18000] = 1'b0;  wr_cycle[18000] = 1'b0;  addr_rom[18000]='h00000000;  wr_data_rom[18000]='h00000000;
    rd_cycle[18001] = 1'b0;  wr_cycle[18001] = 1'b0;  addr_rom[18001]='h00000000;  wr_data_rom[18001]='h00000000;
    rd_cycle[18002] = 1'b0;  wr_cycle[18002] = 1'b0;  addr_rom[18002]='h00000000;  wr_data_rom[18002]='h00000000;
    rd_cycle[18003] = 1'b0;  wr_cycle[18003] = 1'b0;  addr_rom[18003]='h00000000;  wr_data_rom[18003]='h00000000;
    rd_cycle[18004] = 1'b0;  wr_cycle[18004] = 1'b0;  addr_rom[18004]='h00000000;  wr_data_rom[18004]='h00000000;
    rd_cycle[18005] = 1'b0;  wr_cycle[18005] = 1'b0;  addr_rom[18005]='h00000000;  wr_data_rom[18005]='h00000000;
    rd_cycle[18006] = 1'b0;  wr_cycle[18006] = 1'b0;  addr_rom[18006]='h00000000;  wr_data_rom[18006]='h00000000;
    rd_cycle[18007] = 1'b0;  wr_cycle[18007] = 1'b0;  addr_rom[18007]='h00000000;  wr_data_rom[18007]='h00000000;
    rd_cycle[18008] = 1'b0;  wr_cycle[18008] = 1'b0;  addr_rom[18008]='h00000000;  wr_data_rom[18008]='h00000000;
    rd_cycle[18009] = 1'b0;  wr_cycle[18009] = 1'b0;  addr_rom[18009]='h00000000;  wr_data_rom[18009]='h00000000;
    rd_cycle[18010] = 1'b0;  wr_cycle[18010] = 1'b0;  addr_rom[18010]='h00000000;  wr_data_rom[18010]='h00000000;
    rd_cycle[18011] = 1'b0;  wr_cycle[18011] = 1'b0;  addr_rom[18011]='h00000000;  wr_data_rom[18011]='h00000000;
    rd_cycle[18012] = 1'b0;  wr_cycle[18012] = 1'b0;  addr_rom[18012]='h00000000;  wr_data_rom[18012]='h00000000;
    rd_cycle[18013] = 1'b0;  wr_cycle[18013] = 1'b0;  addr_rom[18013]='h00000000;  wr_data_rom[18013]='h00000000;
    rd_cycle[18014] = 1'b0;  wr_cycle[18014] = 1'b0;  addr_rom[18014]='h00000000;  wr_data_rom[18014]='h00000000;
    rd_cycle[18015] = 1'b0;  wr_cycle[18015] = 1'b0;  addr_rom[18015]='h00000000;  wr_data_rom[18015]='h00000000;
    rd_cycle[18016] = 1'b0;  wr_cycle[18016] = 1'b0;  addr_rom[18016]='h00000000;  wr_data_rom[18016]='h00000000;
    rd_cycle[18017] = 1'b0;  wr_cycle[18017] = 1'b0;  addr_rom[18017]='h00000000;  wr_data_rom[18017]='h00000000;
    rd_cycle[18018] = 1'b0;  wr_cycle[18018] = 1'b0;  addr_rom[18018]='h00000000;  wr_data_rom[18018]='h00000000;
    rd_cycle[18019] = 1'b0;  wr_cycle[18019] = 1'b0;  addr_rom[18019]='h00000000;  wr_data_rom[18019]='h00000000;
    rd_cycle[18020] = 1'b0;  wr_cycle[18020] = 1'b0;  addr_rom[18020]='h00000000;  wr_data_rom[18020]='h00000000;
    rd_cycle[18021] = 1'b0;  wr_cycle[18021] = 1'b0;  addr_rom[18021]='h00000000;  wr_data_rom[18021]='h00000000;
    rd_cycle[18022] = 1'b0;  wr_cycle[18022] = 1'b0;  addr_rom[18022]='h00000000;  wr_data_rom[18022]='h00000000;
    rd_cycle[18023] = 1'b0;  wr_cycle[18023] = 1'b0;  addr_rom[18023]='h00000000;  wr_data_rom[18023]='h00000000;
    rd_cycle[18024] = 1'b0;  wr_cycle[18024] = 1'b0;  addr_rom[18024]='h00000000;  wr_data_rom[18024]='h00000000;
    rd_cycle[18025] = 1'b0;  wr_cycle[18025] = 1'b0;  addr_rom[18025]='h00000000;  wr_data_rom[18025]='h00000000;
    rd_cycle[18026] = 1'b0;  wr_cycle[18026] = 1'b0;  addr_rom[18026]='h00000000;  wr_data_rom[18026]='h00000000;
    rd_cycle[18027] = 1'b0;  wr_cycle[18027] = 1'b0;  addr_rom[18027]='h00000000;  wr_data_rom[18027]='h00000000;
    rd_cycle[18028] = 1'b0;  wr_cycle[18028] = 1'b0;  addr_rom[18028]='h00000000;  wr_data_rom[18028]='h00000000;
    rd_cycle[18029] = 1'b0;  wr_cycle[18029] = 1'b0;  addr_rom[18029]='h00000000;  wr_data_rom[18029]='h00000000;
    rd_cycle[18030] = 1'b0;  wr_cycle[18030] = 1'b0;  addr_rom[18030]='h00000000;  wr_data_rom[18030]='h00000000;
    rd_cycle[18031] = 1'b0;  wr_cycle[18031] = 1'b0;  addr_rom[18031]='h00000000;  wr_data_rom[18031]='h00000000;
    rd_cycle[18032] = 1'b0;  wr_cycle[18032] = 1'b0;  addr_rom[18032]='h00000000;  wr_data_rom[18032]='h00000000;
    rd_cycle[18033] = 1'b0;  wr_cycle[18033] = 1'b0;  addr_rom[18033]='h00000000;  wr_data_rom[18033]='h00000000;
    rd_cycle[18034] = 1'b0;  wr_cycle[18034] = 1'b0;  addr_rom[18034]='h00000000;  wr_data_rom[18034]='h00000000;
    rd_cycle[18035] = 1'b0;  wr_cycle[18035] = 1'b0;  addr_rom[18035]='h00000000;  wr_data_rom[18035]='h00000000;
    rd_cycle[18036] = 1'b0;  wr_cycle[18036] = 1'b0;  addr_rom[18036]='h00000000;  wr_data_rom[18036]='h00000000;
    rd_cycle[18037] = 1'b0;  wr_cycle[18037] = 1'b0;  addr_rom[18037]='h00000000;  wr_data_rom[18037]='h00000000;
    rd_cycle[18038] = 1'b0;  wr_cycle[18038] = 1'b0;  addr_rom[18038]='h00000000;  wr_data_rom[18038]='h00000000;
    rd_cycle[18039] = 1'b0;  wr_cycle[18039] = 1'b0;  addr_rom[18039]='h00000000;  wr_data_rom[18039]='h00000000;
    rd_cycle[18040] = 1'b0;  wr_cycle[18040] = 1'b0;  addr_rom[18040]='h00000000;  wr_data_rom[18040]='h00000000;
    rd_cycle[18041] = 1'b0;  wr_cycle[18041] = 1'b0;  addr_rom[18041]='h00000000;  wr_data_rom[18041]='h00000000;
    rd_cycle[18042] = 1'b0;  wr_cycle[18042] = 1'b0;  addr_rom[18042]='h00000000;  wr_data_rom[18042]='h00000000;
    rd_cycle[18043] = 1'b0;  wr_cycle[18043] = 1'b0;  addr_rom[18043]='h00000000;  wr_data_rom[18043]='h00000000;
    rd_cycle[18044] = 1'b0;  wr_cycle[18044] = 1'b0;  addr_rom[18044]='h00000000;  wr_data_rom[18044]='h00000000;
    rd_cycle[18045] = 1'b0;  wr_cycle[18045] = 1'b0;  addr_rom[18045]='h00000000;  wr_data_rom[18045]='h00000000;
    rd_cycle[18046] = 1'b0;  wr_cycle[18046] = 1'b0;  addr_rom[18046]='h00000000;  wr_data_rom[18046]='h00000000;
    rd_cycle[18047] = 1'b0;  wr_cycle[18047] = 1'b0;  addr_rom[18047]='h00000000;  wr_data_rom[18047]='h00000000;
    rd_cycle[18048] = 1'b0;  wr_cycle[18048] = 1'b0;  addr_rom[18048]='h00000000;  wr_data_rom[18048]='h00000000;
    rd_cycle[18049] = 1'b0;  wr_cycle[18049] = 1'b0;  addr_rom[18049]='h00000000;  wr_data_rom[18049]='h00000000;
    rd_cycle[18050] = 1'b0;  wr_cycle[18050] = 1'b0;  addr_rom[18050]='h00000000;  wr_data_rom[18050]='h00000000;
    rd_cycle[18051] = 1'b0;  wr_cycle[18051] = 1'b0;  addr_rom[18051]='h00000000;  wr_data_rom[18051]='h00000000;
    rd_cycle[18052] = 1'b0;  wr_cycle[18052] = 1'b0;  addr_rom[18052]='h00000000;  wr_data_rom[18052]='h00000000;
    rd_cycle[18053] = 1'b0;  wr_cycle[18053] = 1'b0;  addr_rom[18053]='h00000000;  wr_data_rom[18053]='h00000000;
    rd_cycle[18054] = 1'b0;  wr_cycle[18054] = 1'b0;  addr_rom[18054]='h00000000;  wr_data_rom[18054]='h00000000;
    rd_cycle[18055] = 1'b0;  wr_cycle[18055] = 1'b0;  addr_rom[18055]='h00000000;  wr_data_rom[18055]='h00000000;
    rd_cycle[18056] = 1'b0;  wr_cycle[18056] = 1'b0;  addr_rom[18056]='h00000000;  wr_data_rom[18056]='h00000000;
    rd_cycle[18057] = 1'b0;  wr_cycle[18057] = 1'b0;  addr_rom[18057]='h00000000;  wr_data_rom[18057]='h00000000;
    rd_cycle[18058] = 1'b0;  wr_cycle[18058] = 1'b0;  addr_rom[18058]='h00000000;  wr_data_rom[18058]='h00000000;
    rd_cycle[18059] = 1'b0;  wr_cycle[18059] = 1'b0;  addr_rom[18059]='h00000000;  wr_data_rom[18059]='h00000000;
    rd_cycle[18060] = 1'b0;  wr_cycle[18060] = 1'b0;  addr_rom[18060]='h00000000;  wr_data_rom[18060]='h00000000;
    rd_cycle[18061] = 1'b0;  wr_cycle[18061] = 1'b0;  addr_rom[18061]='h00000000;  wr_data_rom[18061]='h00000000;
    rd_cycle[18062] = 1'b0;  wr_cycle[18062] = 1'b0;  addr_rom[18062]='h00000000;  wr_data_rom[18062]='h00000000;
    rd_cycle[18063] = 1'b0;  wr_cycle[18063] = 1'b0;  addr_rom[18063]='h00000000;  wr_data_rom[18063]='h00000000;
    rd_cycle[18064] = 1'b0;  wr_cycle[18064] = 1'b0;  addr_rom[18064]='h00000000;  wr_data_rom[18064]='h00000000;
    rd_cycle[18065] = 1'b0;  wr_cycle[18065] = 1'b0;  addr_rom[18065]='h00000000;  wr_data_rom[18065]='h00000000;
    rd_cycle[18066] = 1'b0;  wr_cycle[18066] = 1'b0;  addr_rom[18066]='h00000000;  wr_data_rom[18066]='h00000000;
    rd_cycle[18067] = 1'b0;  wr_cycle[18067] = 1'b0;  addr_rom[18067]='h00000000;  wr_data_rom[18067]='h00000000;
    rd_cycle[18068] = 1'b0;  wr_cycle[18068] = 1'b0;  addr_rom[18068]='h00000000;  wr_data_rom[18068]='h00000000;
    rd_cycle[18069] = 1'b0;  wr_cycle[18069] = 1'b0;  addr_rom[18069]='h00000000;  wr_data_rom[18069]='h00000000;
    rd_cycle[18070] = 1'b0;  wr_cycle[18070] = 1'b0;  addr_rom[18070]='h00000000;  wr_data_rom[18070]='h00000000;
    rd_cycle[18071] = 1'b0;  wr_cycle[18071] = 1'b0;  addr_rom[18071]='h00000000;  wr_data_rom[18071]='h00000000;
    rd_cycle[18072] = 1'b0;  wr_cycle[18072] = 1'b0;  addr_rom[18072]='h00000000;  wr_data_rom[18072]='h00000000;
    rd_cycle[18073] = 1'b0;  wr_cycle[18073] = 1'b0;  addr_rom[18073]='h00000000;  wr_data_rom[18073]='h00000000;
    rd_cycle[18074] = 1'b0;  wr_cycle[18074] = 1'b0;  addr_rom[18074]='h00000000;  wr_data_rom[18074]='h00000000;
    rd_cycle[18075] = 1'b0;  wr_cycle[18075] = 1'b0;  addr_rom[18075]='h00000000;  wr_data_rom[18075]='h00000000;
    rd_cycle[18076] = 1'b0;  wr_cycle[18076] = 1'b0;  addr_rom[18076]='h00000000;  wr_data_rom[18076]='h00000000;
    rd_cycle[18077] = 1'b0;  wr_cycle[18077] = 1'b0;  addr_rom[18077]='h00000000;  wr_data_rom[18077]='h00000000;
    rd_cycle[18078] = 1'b0;  wr_cycle[18078] = 1'b0;  addr_rom[18078]='h00000000;  wr_data_rom[18078]='h00000000;
    rd_cycle[18079] = 1'b0;  wr_cycle[18079] = 1'b0;  addr_rom[18079]='h00000000;  wr_data_rom[18079]='h00000000;
    rd_cycle[18080] = 1'b0;  wr_cycle[18080] = 1'b0;  addr_rom[18080]='h00000000;  wr_data_rom[18080]='h00000000;
    rd_cycle[18081] = 1'b0;  wr_cycle[18081] = 1'b0;  addr_rom[18081]='h00000000;  wr_data_rom[18081]='h00000000;
    rd_cycle[18082] = 1'b0;  wr_cycle[18082] = 1'b0;  addr_rom[18082]='h00000000;  wr_data_rom[18082]='h00000000;
    rd_cycle[18083] = 1'b0;  wr_cycle[18083] = 1'b0;  addr_rom[18083]='h00000000;  wr_data_rom[18083]='h00000000;
    rd_cycle[18084] = 1'b0;  wr_cycle[18084] = 1'b0;  addr_rom[18084]='h00000000;  wr_data_rom[18084]='h00000000;
    rd_cycle[18085] = 1'b0;  wr_cycle[18085] = 1'b0;  addr_rom[18085]='h00000000;  wr_data_rom[18085]='h00000000;
    rd_cycle[18086] = 1'b0;  wr_cycle[18086] = 1'b0;  addr_rom[18086]='h00000000;  wr_data_rom[18086]='h00000000;
    rd_cycle[18087] = 1'b0;  wr_cycle[18087] = 1'b0;  addr_rom[18087]='h00000000;  wr_data_rom[18087]='h00000000;
    rd_cycle[18088] = 1'b0;  wr_cycle[18088] = 1'b0;  addr_rom[18088]='h00000000;  wr_data_rom[18088]='h00000000;
    rd_cycle[18089] = 1'b0;  wr_cycle[18089] = 1'b0;  addr_rom[18089]='h00000000;  wr_data_rom[18089]='h00000000;
    rd_cycle[18090] = 1'b0;  wr_cycle[18090] = 1'b0;  addr_rom[18090]='h00000000;  wr_data_rom[18090]='h00000000;
    rd_cycle[18091] = 1'b0;  wr_cycle[18091] = 1'b0;  addr_rom[18091]='h00000000;  wr_data_rom[18091]='h00000000;
    rd_cycle[18092] = 1'b0;  wr_cycle[18092] = 1'b0;  addr_rom[18092]='h00000000;  wr_data_rom[18092]='h00000000;
    rd_cycle[18093] = 1'b0;  wr_cycle[18093] = 1'b0;  addr_rom[18093]='h00000000;  wr_data_rom[18093]='h00000000;
    rd_cycle[18094] = 1'b0;  wr_cycle[18094] = 1'b0;  addr_rom[18094]='h00000000;  wr_data_rom[18094]='h00000000;
    rd_cycle[18095] = 1'b0;  wr_cycle[18095] = 1'b0;  addr_rom[18095]='h00000000;  wr_data_rom[18095]='h00000000;
    rd_cycle[18096] = 1'b0;  wr_cycle[18096] = 1'b0;  addr_rom[18096]='h00000000;  wr_data_rom[18096]='h00000000;
    rd_cycle[18097] = 1'b0;  wr_cycle[18097] = 1'b0;  addr_rom[18097]='h00000000;  wr_data_rom[18097]='h00000000;
    rd_cycle[18098] = 1'b0;  wr_cycle[18098] = 1'b0;  addr_rom[18098]='h00000000;  wr_data_rom[18098]='h00000000;
    rd_cycle[18099] = 1'b0;  wr_cycle[18099] = 1'b0;  addr_rom[18099]='h00000000;  wr_data_rom[18099]='h00000000;
    rd_cycle[18100] = 1'b0;  wr_cycle[18100] = 1'b0;  addr_rom[18100]='h00000000;  wr_data_rom[18100]='h00000000;
    rd_cycle[18101] = 1'b0;  wr_cycle[18101] = 1'b0;  addr_rom[18101]='h00000000;  wr_data_rom[18101]='h00000000;
    rd_cycle[18102] = 1'b0;  wr_cycle[18102] = 1'b0;  addr_rom[18102]='h00000000;  wr_data_rom[18102]='h00000000;
    rd_cycle[18103] = 1'b0;  wr_cycle[18103] = 1'b0;  addr_rom[18103]='h00000000;  wr_data_rom[18103]='h00000000;
    rd_cycle[18104] = 1'b0;  wr_cycle[18104] = 1'b0;  addr_rom[18104]='h00000000;  wr_data_rom[18104]='h00000000;
    rd_cycle[18105] = 1'b0;  wr_cycle[18105] = 1'b0;  addr_rom[18105]='h00000000;  wr_data_rom[18105]='h00000000;
    rd_cycle[18106] = 1'b0;  wr_cycle[18106] = 1'b0;  addr_rom[18106]='h00000000;  wr_data_rom[18106]='h00000000;
    rd_cycle[18107] = 1'b0;  wr_cycle[18107] = 1'b0;  addr_rom[18107]='h00000000;  wr_data_rom[18107]='h00000000;
    rd_cycle[18108] = 1'b0;  wr_cycle[18108] = 1'b0;  addr_rom[18108]='h00000000;  wr_data_rom[18108]='h00000000;
    rd_cycle[18109] = 1'b0;  wr_cycle[18109] = 1'b0;  addr_rom[18109]='h00000000;  wr_data_rom[18109]='h00000000;
    rd_cycle[18110] = 1'b0;  wr_cycle[18110] = 1'b0;  addr_rom[18110]='h00000000;  wr_data_rom[18110]='h00000000;
    rd_cycle[18111] = 1'b0;  wr_cycle[18111] = 1'b0;  addr_rom[18111]='h00000000;  wr_data_rom[18111]='h00000000;
    rd_cycle[18112] = 1'b0;  wr_cycle[18112] = 1'b0;  addr_rom[18112]='h00000000;  wr_data_rom[18112]='h00000000;
    rd_cycle[18113] = 1'b0;  wr_cycle[18113] = 1'b0;  addr_rom[18113]='h00000000;  wr_data_rom[18113]='h00000000;
    rd_cycle[18114] = 1'b0;  wr_cycle[18114] = 1'b0;  addr_rom[18114]='h00000000;  wr_data_rom[18114]='h00000000;
    rd_cycle[18115] = 1'b0;  wr_cycle[18115] = 1'b0;  addr_rom[18115]='h00000000;  wr_data_rom[18115]='h00000000;
    rd_cycle[18116] = 1'b0;  wr_cycle[18116] = 1'b0;  addr_rom[18116]='h00000000;  wr_data_rom[18116]='h00000000;
    rd_cycle[18117] = 1'b0;  wr_cycle[18117] = 1'b0;  addr_rom[18117]='h00000000;  wr_data_rom[18117]='h00000000;
    rd_cycle[18118] = 1'b0;  wr_cycle[18118] = 1'b0;  addr_rom[18118]='h00000000;  wr_data_rom[18118]='h00000000;
    rd_cycle[18119] = 1'b0;  wr_cycle[18119] = 1'b0;  addr_rom[18119]='h00000000;  wr_data_rom[18119]='h00000000;
    rd_cycle[18120] = 1'b0;  wr_cycle[18120] = 1'b0;  addr_rom[18120]='h00000000;  wr_data_rom[18120]='h00000000;
    rd_cycle[18121] = 1'b0;  wr_cycle[18121] = 1'b0;  addr_rom[18121]='h00000000;  wr_data_rom[18121]='h00000000;
    rd_cycle[18122] = 1'b0;  wr_cycle[18122] = 1'b0;  addr_rom[18122]='h00000000;  wr_data_rom[18122]='h00000000;
    rd_cycle[18123] = 1'b0;  wr_cycle[18123] = 1'b0;  addr_rom[18123]='h00000000;  wr_data_rom[18123]='h00000000;
    rd_cycle[18124] = 1'b0;  wr_cycle[18124] = 1'b0;  addr_rom[18124]='h00000000;  wr_data_rom[18124]='h00000000;
    rd_cycle[18125] = 1'b0;  wr_cycle[18125] = 1'b0;  addr_rom[18125]='h00000000;  wr_data_rom[18125]='h00000000;
    rd_cycle[18126] = 1'b0;  wr_cycle[18126] = 1'b0;  addr_rom[18126]='h00000000;  wr_data_rom[18126]='h00000000;
    rd_cycle[18127] = 1'b0;  wr_cycle[18127] = 1'b0;  addr_rom[18127]='h00000000;  wr_data_rom[18127]='h00000000;
    rd_cycle[18128] = 1'b0;  wr_cycle[18128] = 1'b0;  addr_rom[18128]='h00000000;  wr_data_rom[18128]='h00000000;
    rd_cycle[18129] = 1'b0;  wr_cycle[18129] = 1'b0;  addr_rom[18129]='h00000000;  wr_data_rom[18129]='h00000000;
    rd_cycle[18130] = 1'b0;  wr_cycle[18130] = 1'b0;  addr_rom[18130]='h00000000;  wr_data_rom[18130]='h00000000;
    rd_cycle[18131] = 1'b0;  wr_cycle[18131] = 1'b0;  addr_rom[18131]='h00000000;  wr_data_rom[18131]='h00000000;
    rd_cycle[18132] = 1'b0;  wr_cycle[18132] = 1'b0;  addr_rom[18132]='h00000000;  wr_data_rom[18132]='h00000000;
    rd_cycle[18133] = 1'b0;  wr_cycle[18133] = 1'b0;  addr_rom[18133]='h00000000;  wr_data_rom[18133]='h00000000;
    rd_cycle[18134] = 1'b0;  wr_cycle[18134] = 1'b0;  addr_rom[18134]='h00000000;  wr_data_rom[18134]='h00000000;
    rd_cycle[18135] = 1'b0;  wr_cycle[18135] = 1'b0;  addr_rom[18135]='h00000000;  wr_data_rom[18135]='h00000000;
    rd_cycle[18136] = 1'b0;  wr_cycle[18136] = 1'b0;  addr_rom[18136]='h00000000;  wr_data_rom[18136]='h00000000;
    rd_cycle[18137] = 1'b0;  wr_cycle[18137] = 1'b0;  addr_rom[18137]='h00000000;  wr_data_rom[18137]='h00000000;
    rd_cycle[18138] = 1'b0;  wr_cycle[18138] = 1'b0;  addr_rom[18138]='h00000000;  wr_data_rom[18138]='h00000000;
    rd_cycle[18139] = 1'b0;  wr_cycle[18139] = 1'b0;  addr_rom[18139]='h00000000;  wr_data_rom[18139]='h00000000;
    rd_cycle[18140] = 1'b0;  wr_cycle[18140] = 1'b0;  addr_rom[18140]='h00000000;  wr_data_rom[18140]='h00000000;
    rd_cycle[18141] = 1'b0;  wr_cycle[18141] = 1'b0;  addr_rom[18141]='h00000000;  wr_data_rom[18141]='h00000000;
    rd_cycle[18142] = 1'b0;  wr_cycle[18142] = 1'b0;  addr_rom[18142]='h00000000;  wr_data_rom[18142]='h00000000;
    rd_cycle[18143] = 1'b0;  wr_cycle[18143] = 1'b0;  addr_rom[18143]='h00000000;  wr_data_rom[18143]='h00000000;
    rd_cycle[18144] = 1'b0;  wr_cycle[18144] = 1'b0;  addr_rom[18144]='h00000000;  wr_data_rom[18144]='h00000000;
    rd_cycle[18145] = 1'b0;  wr_cycle[18145] = 1'b0;  addr_rom[18145]='h00000000;  wr_data_rom[18145]='h00000000;
    rd_cycle[18146] = 1'b0;  wr_cycle[18146] = 1'b0;  addr_rom[18146]='h00000000;  wr_data_rom[18146]='h00000000;
    rd_cycle[18147] = 1'b0;  wr_cycle[18147] = 1'b0;  addr_rom[18147]='h00000000;  wr_data_rom[18147]='h00000000;
    rd_cycle[18148] = 1'b0;  wr_cycle[18148] = 1'b0;  addr_rom[18148]='h00000000;  wr_data_rom[18148]='h00000000;
    rd_cycle[18149] = 1'b0;  wr_cycle[18149] = 1'b0;  addr_rom[18149]='h00000000;  wr_data_rom[18149]='h00000000;
    rd_cycle[18150] = 1'b0;  wr_cycle[18150] = 1'b0;  addr_rom[18150]='h00000000;  wr_data_rom[18150]='h00000000;
    rd_cycle[18151] = 1'b0;  wr_cycle[18151] = 1'b0;  addr_rom[18151]='h00000000;  wr_data_rom[18151]='h00000000;
    rd_cycle[18152] = 1'b0;  wr_cycle[18152] = 1'b0;  addr_rom[18152]='h00000000;  wr_data_rom[18152]='h00000000;
    rd_cycle[18153] = 1'b0;  wr_cycle[18153] = 1'b0;  addr_rom[18153]='h00000000;  wr_data_rom[18153]='h00000000;
    rd_cycle[18154] = 1'b0;  wr_cycle[18154] = 1'b0;  addr_rom[18154]='h00000000;  wr_data_rom[18154]='h00000000;
    rd_cycle[18155] = 1'b0;  wr_cycle[18155] = 1'b0;  addr_rom[18155]='h00000000;  wr_data_rom[18155]='h00000000;
    rd_cycle[18156] = 1'b0;  wr_cycle[18156] = 1'b0;  addr_rom[18156]='h00000000;  wr_data_rom[18156]='h00000000;
    rd_cycle[18157] = 1'b0;  wr_cycle[18157] = 1'b0;  addr_rom[18157]='h00000000;  wr_data_rom[18157]='h00000000;
    rd_cycle[18158] = 1'b0;  wr_cycle[18158] = 1'b0;  addr_rom[18158]='h00000000;  wr_data_rom[18158]='h00000000;
    rd_cycle[18159] = 1'b0;  wr_cycle[18159] = 1'b0;  addr_rom[18159]='h00000000;  wr_data_rom[18159]='h00000000;
    rd_cycle[18160] = 1'b0;  wr_cycle[18160] = 1'b0;  addr_rom[18160]='h00000000;  wr_data_rom[18160]='h00000000;
    rd_cycle[18161] = 1'b0;  wr_cycle[18161] = 1'b0;  addr_rom[18161]='h00000000;  wr_data_rom[18161]='h00000000;
    rd_cycle[18162] = 1'b0;  wr_cycle[18162] = 1'b0;  addr_rom[18162]='h00000000;  wr_data_rom[18162]='h00000000;
    rd_cycle[18163] = 1'b0;  wr_cycle[18163] = 1'b0;  addr_rom[18163]='h00000000;  wr_data_rom[18163]='h00000000;
    rd_cycle[18164] = 1'b0;  wr_cycle[18164] = 1'b0;  addr_rom[18164]='h00000000;  wr_data_rom[18164]='h00000000;
    rd_cycle[18165] = 1'b0;  wr_cycle[18165] = 1'b0;  addr_rom[18165]='h00000000;  wr_data_rom[18165]='h00000000;
    rd_cycle[18166] = 1'b0;  wr_cycle[18166] = 1'b0;  addr_rom[18166]='h00000000;  wr_data_rom[18166]='h00000000;
    rd_cycle[18167] = 1'b0;  wr_cycle[18167] = 1'b0;  addr_rom[18167]='h00000000;  wr_data_rom[18167]='h00000000;
    rd_cycle[18168] = 1'b0;  wr_cycle[18168] = 1'b0;  addr_rom[18168]='h00000000;  wr_data_rom[18168]='h00000000;
    rd_cycle[18169] = 1'b0;  wr_cycle[18169] = 1'b0;  addr_rom[18169]='h00000000;  wr_data_rom[18169]='h00000000;
    rd_cycle[18170] = 1'b0;  wr_cycle[18170] = 1'b0;  addr_rom[18170]='h00000000;  wr_data_rom[18170]='h00000000;
    rd_cycle[18171] = 1'b0;  wr_cycle[18171] = 1'b0;  addr_rom[18171]='h00000000;  wr_data_rom[18171]='h00000000;
    rd_cycle[18172] = 1'b0;  wr_cycle[18172] = 1'b0;  addr_rom[18172]='h00000000;  wr_data_rom[18172]='h00000000;
    rd_cycle[18173] = 1'b0;  wr_cycle[18173] = 1'b0;  addr_rom[18173]='h00000000;  wr_data_rom[18173]='h00000000;
    rd_cycle[18174] = 1'b0;  wr_cycle[18174] = 1'b0;  addr_rom[18174]='h00000000;  wr_data_rom[18174]='h00000000;
    rd_cycle[18175] = 1'b0;  wr_cycle[18175] = 1'b0;  addr_rom[18175]='h00000000;  wr_data_rom[18175]='h00000000;
    rd_cycle[18176] = 1'b0;  wr_cycle[18176] = 1'b0;  addr_rom[18176]='h00000000;  wr_data_rom[18176]='h00000000;
    rd_cycle[18177] = 1'b0;  wr_cycle[18177] = 1'b0;  addr_rom[18177]='h00000000;  wr_data_rom[18177]='h00000000;
    rd_cycle[18178] = 1'b0;  wr_cycle[18178] = 1'b0;  addr_rom[18178]='h00000000;  wr_data_rom[18178]='h00000000;
    rd_cycle[18179] = 1'b0;  wr_cycle[18179] = 1'b0;  addr_rom[18179]='h00000000;  wr_data_rom[18179]='h00000000;
    rd_cycle[18180] = 1'b0;  wr_cycle[18180] = 1'b0;  addr_rom[18180]='h00000000;  wr_data_rom[18180]='h00000000;
    rd_cycle[18181] = 1'b0;  wr_cycle[18181] = 1'b0;  addr_rom[18181]='h00000000;  wr_data_rom[18181]='h00000000;
    rd_cycle[18182] = 1'b0;  wr_cycle[18182] = 1'b0;  addr_rom[18182]='h00000000;  wr_data_rom[18182]='h00000000;
    rd_cycle[18183] = 1'b0;  wr_cycle[18183] = 1'b0;  addr_rom[18183]='h00000000;  wr_data_rom[18183]='h00000000;
    rd_cycle[18184] = 1'b0;  wr_cycle[18184] = 1'b0;  addr_rom[18184]='h00000000;  wr_data_rom[18184]='h00000000;
    rd_cycle[18185] = 1'b0;  wr_cycle[18185] = 1'b0;  addr_rom[18185]='h00000000;  wr_data_rom[18185]='h00000000;
    rd_cycle[18186] = 1'b0;  wr_cycle[18186] = 1'b0;  addr_rom[18186]='h00000000;  wr_data_rom[18186]='h00000000;
    rd_cycle[18187] = 1'b0;  wr_cycle[18187] = 1'b0;  addr_rom[18187]='h00000000;  wr_data_rom[18187]='h00000000;
    rd_cycle[18188] = 1'b0;  wr_cycle[18188] = 1'b0;  addr_rom[18188]='h00000000;  wr_data_rom[18188]='h00000000;
    rd_cycle[18189] = 1'b0;  wr_cycle[18189] = 1'b0;  addr_rom[18189]='h00000000;  wr_data_rom[18189]='h00000000;
    rd_cycle[18190] = 1'b0;  wr_cycle[18190] = 1'b0;  addr_rom[18190]='h00000000;  wr_data_rom[18190]='h00000000;
    rd_cycle[18191] = 1'b0;  wr_cycle[18191] = 1'b0;  addr_rom[18191]='h00000000;  wr_data_rom[18191]='h00000000;
    rd_cycle[18192] = 1'b0;  wr_cycle[18192] = 1'b0;  addr_rom[18192]='h00000000;  wr_data_rom[18192]='h00000000;
    rd_cycle[18193] = 1'b0;  wr_cycle[18193] = 1'b0;  addr_rom[18193]='h00000000;  wr_data_rom[18193]='h00000000;
    rd_cycle[18194] = 1'b0;  wr_cycle[18194] = 1'b0;  addr_rom[18194]='h00000000;  wr_data_rom[18194]='h00000000;
    rd_cycle[18195] = 1'b0;  wr_cycle[18195] = 1'b0;  addr_rom[18195]='h00000000;  wr_data_rom[18195]='h00000000;
    rd_cycle[18196] = 1'b0;  wr_cycle[18196] = 1'b0;  addr_rom[18196]='h00000000;  wr_data_rom[18196]='h00000000;
    rd_cycle[18197] = 1'b0;  wr_cycle[18197] = 1'b0;  addr_rom[18197]='h00000000;  wr_data_rom[18197]='h00000000;
    rd_cycle[18198] = 1'b0;  wr_cycle[18198] = 1'b0;  addr_rom[18198]='h00000000;  wr_data_rom[18198]='h00000000;
    rd_cycle[18199] = 1'b0;  wr_cycle[18199] = 1'b0;  addr_rom[18199]='h00000000;  wr_data_rom[18199]='h00000000;
    rd_cycle[18200] = 1'b0;  wr_cycle[18200] = 1'b0;  addr_rom[18200]='h00000000;  wr_data_rom[18200]='h00000000;
    rd_cycle[18201] = 1'b0;  wr_cycle[18201] = 1'b0;  addr_rom[18201]='h00000000;  wr_data_rom[18201]='h00000000;
    rd_cycle[18202] = 1'b0;  wr_cycle[18202] = 1'b0;  addr_rom[18202]='h00000000;  wr_data_rom[18202]='h00000000;
    rd_cycle[18203] = 1'b0;  wr_cycle[18203] = 1'b0;  addr_rom[18203]='h00000000;  wr_data_rom[18203]='h00000000;
    rd_cycle[18204] = 1'b0;  wr_cycle[18204] = 1'b0;  addr_rom[18204]='h00000000;  wr_data_rom[18204]='h00000000;
    rd_cycle[18205] = 1'b0;  wr_cycle[18205] = 1'b0;  addr_rom[18205]='h00000000;  wr_data_rom[18205]='h00000000;
    rd_cycle[18206] = 1'b0;  wr_cycle[18206] = 1'b0;  addr_rom[18206]='h00000000;  wr_data_rom[18206]='h00000000;
    rd_cycle[18207] = 1'b0;  wr_cycle[18207] = 1'b0;  addr_rom[18207]='h00000000;  wr_data_rom[18207]='h00000000;
    rd_cycle[18208] = 1'b0;  wr_cycle[18208] = 1'b0;  addr_rom[18208]='h00000000;  wr_data_rom[18208]='h00000000;
    rd_cycle[18209] = 1'b0;  wr_cycle[18209] = 1'b0;  addr_rom[18209]='h00000000;  wr_data_rom[18209]='h00000000;
    rd_cycle[18210] = 1'b0;  wr_cycle[18210] = 1'b0;  addr_rom[18210]='h00000000;  wr_data_rom[18210]='h00000000;
    rd_cycle[18211] = 1'b0;  wr_cycle[18211] = 1'b0;  addr_rom[18211]='h00000000;  wr_data_rom[18211]='h00000000;
    rd_cycle[18212] = 1'b0;  wr_cycle[18212] = 1'b0;  addr_rom[18212]='h00000000;  wr_data_rom[18212]='h00000000;
    rd_cycle[18213] = 1'b0;  wr_cycle[18213] = 1'b0;  addr_rom[18213]='h00000000;  wr_data_rom[18213]='h00000000;
    rd_cycle[18214] = 1'b0;  wr_cycle[18214] = 1'b0;  addr_rom[18214]='h00000000;  wr_data_rom[18214]='h00000000;
    rd_cycle[18215] = 1'b0;  wr_cycle[18215] = 1'b0;  addr_rom[18215]='h00000000;  wr_data_rom[18215]='h00000000;
    rd_cycle[18216] = 1'b0;  wr_cycle[18216] = 1'b0;  addr_rom[18216]='h00000000;  wr_data_rom[18216]='h00000000;
    rd_cycle[18217] = 1'b0;  wr_cycle[18217] = 1'b0;  addr_rom[18217]='h00000000;  wr_data_rom[18217]='h00000000;
    rd_cycle[18218] = 1'b0;  wr_cycle[18218] = 1'b0;  addr_rom[18218]='h00000000;  wr_data_rom[18218]='h00000000;
    rd_cycle[18219] = 1'b0;  wr_cycle[18219] = 1'b0;  addr_rom[18219]='h00000000;  wr_data_rom[18219]='h00000000;
    rd_cycle[18220] = 1'b0;  wr_cycle[18220] = 1'b0;  addr_rom[18220]='h00000000;  wr_data_rom[18220]='h00000000;
    rd_cycle[18221] = 1'b0;  wr_cycle[18221] = 1'b0;  addr_rom[18221]='h00000000;  wr_data_rom[18221]='h00000000;
    rd_cycle[18222] = 1'b0;  wr_cycle[18222] = 1'b0;  addr_rom[18222]='h00000000;  wr_data_rom[18222]='h00000000;
    rd_cycle[18223] = 1'b0;  wr_cycle[18223] = 1'b0;  addr_rom[18223]='h00000000;  wr_data_rom[18223]='h00000000;
    rd_cycle[18224] = 1'b0;  wr_cycle[18224] = 1'b0;  addr_rom[18224]='h00000000;  wr_data_rom[18224]='h00000000;
    rd_cycle[18225] = 1'b0;  wr_cycle[18225] = 1'b0;  addr_rom[18225]='h00000000;  wr_data_rom[18225]='h00000000;
    rd_cycle[18226] = 1'b0;  wr_cycle[18226] = 1'b0;  addr_rom[18226]='h00000000;  wr_data_rom[18226]='h00000000;
    rd_cycle[18227] = 1'b0;  wr_cycle[18227] = 1'b0;  addr_rom[18227]='h00000000;  wr_data_rom[18227]='h00000000;
    rd_cycle[18228] = 1'b0;  wr_cycle[18228] = 1'b0;  addr_rom[18228]='h00000000;  wr_data_rom[18228]='h00000000;
    rd_cycle[18229] = 1'b0;  wr_cycle[18229] = 1'b0;  addr_rom[18229]='h00000000;  wr_data_rom[18229]='h00000000;
    rd_cycle[18230] = 1'b0;  wr_cycle[18230] = 1'b0;  addr_rom[18230]='h00000000;  wr_data_rom[18230]='h00000000;
    rd_cycle[18231] = 1'b0;  wr_cycle[18231] = 1'b0;  addr_rom[18231]='h00000000;  wr_data_rom[18231]='h00000000;
    rd_cycle[18232] = 1'b0;  wr_cycle[18232] = 1'b0;  addr_rom[18232]='h00000000;  wr_data_rom[18232]='h00000000;
    rd_cycle[18233] = 1'b0;  wr_cycle[18233] = 1'b0;  addr_rom[18233]='h00000000;  wr_data_rom[18233]='h00000000;
    rd_cycle[18234] = 1'b0;  wr_cycle[18234] = 1'b0;  addr_rom[18234]='h00000000;  wr_data_rom[18234]='h00000000;
    rd_cycle[18235] = 1'b0;  wr_cycle[18235] = 1'b0;  addr_rom[18235]='h00000000;  wr_data_rom[18235]='h00000000;
    rd_cycle[18236] = 1'b0;  wr_cycle[18236] = 1'b0;  addr_rom[18236]='h00000000;  wr_data_rom[18236]='h00000000;
    rd_cycle[18237] = 1'b0;  wr_cycle[18237] = 1'b0;  addr_rom[18237]='h00000000;  wr_data_rom[18237]='h00000000;
    rd_cycle[18238] = 1'b0;  wr_cycle[18238] = 1'b0;  addr_rom[18238]='h00000000;  wr_data_rom[18238]='h00000000;
    rd_cycle[18239] = 1'b0;  wr_cycle[18239] = 1'b0;  addr_rom[18239]='h00000000;  wr_data_rom[18239]='h00000000;
    rd_cycle[18240] = 1'b0;  wr_cycle[18240] = 1'b0;  addr_rom[18240]='h00000000;  wr_data_rom[18240]='h00000000;
    rd_cycle[18241] = 1'b0;  wr_cycle[18241] = 1'b0;  addr_rom[18241]='h00000000;  wr_data_rom[18241]='h00000000;
    rd_cycle[18242] = 1'b0;  wr_cycle[18242] = 1'b0;  addr_rom[18242]='h00000000;  wr_data_rom[18242]='h00000000;
    rd_cycle[18243] = 1'b0;  wr_cycle[18243] = 1'b0;  addr_rom[18243]='h00000000;  wr_data_rom[18243]='h00000000;
    rd_cycle[18244] = 1'b0;  wr_cycle[18244] = 1'b0;  addr_rom[18244]='h00000000;  wr_data_rom[18244]='h00000000;
    rd_cycle[18245] = 1'b0;  wr_cycle[18245] = 1'b0;  addr_rom[18245]='h00000000;  wr_data_rom[18245]='h00000000;
    rd_cycle[18246] = 1'b0;  wr_cycle[18246] = 1'b0;  addr_rom[18246]='h00000000;  wr_data_rom[18246]='h00000000;
    rd_cycle[18247] = 1'b0;  wr_cycle[18247] = 1'b0;  addr_rom[18247]='h00000000;  wr_data_rom[18247]='h00000000;
    rd_cycle[18248] = 1'b0;  wr_cycle[18248] = 1'b0;  addr_rom[18248]='h00000000;  wr_data_rom[18248]='h00000000;
    rd_cycle[18249] = 1'b0;  wr_cycle[18249] = 1'b0;  addr_rom[18249]='h00000000;  wr_data_rom[18249]='h00000000;
    rd_cycle[18250] = 1'b0;  wr_cycle[18250] = 1'b0;  addr_rom[18250]='h00000000;  wr_data_rom[18250]='h00000000;
    rd_cycle[18251] = 1'b0;  wr_cycle[18251] = 1'b0;  addr_rom[18251]='h00000000;  wr_data_rom[18251]='h00000000;
    rd_cycle[18252] = 1'b0;  wr_cycle[18252] = 1'b0;  addr_rom[18252]='h00000000;  wr_data_rom[18252]='h00000000;
    rd_cycle[18253] = 1'b0;  wr_cycle[18253] = 1'b0;  addr_rom[18253]='h00000000;  wr_data_rom[18253]='h00000000;
    rd_cycle[18254] = 1'b0;  wr_cycle[18254] = 1'b0;  addr_rom[18254]='h00000000;  wr_data_rom[18254]='h00000000;
    rd_cycle[18255] = 1'b0;  wr_cycle[18255] = 1'b0;  addr_rom[18255]='h00000000;  wr_data_rom[18255]='h00000000;
    rd_cycle[18256] = 1'b0;  wr_cycle[18256] = 1'b0;  addr_rom[18256]='h00000000;  wr_data_rom[18256]='h00000000;
    rd_cycle[18257] = 1'b0;  wr_cycle[18257] = 1'b0;  addr_rom[18257]='h00000000;  wr_data_rom[18257]='h00000000;
    rd_cycle[18258] = 1'b0;  wr_cycle[18258] = 1'b0;  addr_rom[18258]='h00000000;  wr_data_rom[18258]='h00000000;
    rd_cycle[18259] = 1'b0;  wr_cycle[18259] = 1'b0;  addr_rom[18259]='h00000000;  wr_data_rom[18259]='h00000000;
    rd_cycle[18260] = 1'b0;  wr_cycle[18260] = 1'b0;  addr_rom[18260]='h00000000;  wr_data_rom[18260]='h00000000;
    rd_cycle[18261] = 1'b0;  wr_cycle[18261] = 1'b0;  addr_rom[18261]='h00000000;  wr_data_rom[18261]='h00000000;
    rd_cycle[18262] = 1'b0;  wr_cycle[18262] = 1'b0;  addr_rom[18262]='h00000000;  wr_data_rom[18262]='h00000000;
    rd_cycle[18263] = 1'b0;  wr_cycle[18263] = 1'b0;  addr_rom[18263]='h00000000;  wr_data_rom[18263]='h00000000;
    rd_cycle[18264] = 1'b0;  wr_cycle[18264] = 1'b0;  addr_rom[18264]='h00000000;  wr_data_rom[18264]='h00000000;
    rd_cycle[18265] = 1'b0;  wr_cycle[18265] = 1'b0;  addr_rom[18265]='h00000000;  wr_data_rom[18265]='h00000000;
    rd_cycle[18266] = 1'b0;  wr_cycle[18266] = 1'b0;  addr_rom[18266]='h00000000;  wr_data_rom[18266]='h00000000;
    rd_cycle[18267] = 1'b0;  wr_cycle[18267] = 1'b0;  addr_rom[18267]='h00000000;  wr_data_rom[18267]='h00000000;
    rd_cycle[18268] = 1'b0;  wr_cycle[18268] = 1'b0;  addr_rom[18268]='h00000000;  wr_data_rom[18268]='h00000000;
    rd_cycle[18269] = 1'b0;  wr_cycle[18269] = 1'b0;  addr_rom[18269]='h00000000;  wr_data_rom[18269]='h00000000;
    rd_cycle[18270] = 1'b0;  wr_cycle[18270] = 1'b0;  addr_rom[18270]='h00000000;  wr_data_rom[18270]='h00000000;
    rd_cycle[18271] = 1'b0;  wr_cycle[18271] = 1'b0;  addr_rom[18271]='h00000000;  wr_data_rom[18271]='h00000000;
    rd_cycle[18272] = 1'b0;  wr_cycle[18272] = 1'b0;  addr_rom[18272]='h00000000;  wr_data_rom[18272]='h00000000;
    rd_cycle[18273] = 1'b0;  wr_cycle[18273] = 1'b0;  addr_rom[18273]='h00000000;  wr_data_rom[18273]='h00000000;
    rd_cycle[18274] = 1'b0;  wr_cycle[18274] = 1'b0;  addr_rom[18274]='h00000000;  wr_data_rom[18274]='h00000000;
    rd_cycle[18275] = 1'b0;  wr_cycle[18275] = 1'b0;  addr_rom[18275]='h00000000;  wr_data_rom[18275]='h00000000;
    rd_cycle[18276] = 1'b0;  wr_cycle[18276] = 1'b0;  addr_rom[18276]='h00000000;  wr_data_rom[18276]='h00000000;
    rd_cycle[18277] = 1'b0;  wr_cycle[18277] = 1'b0;  addr_rom[18277]='h00000000;  wr_data_rom[18277]='h00000000;
    rd_cycle[18278] = 1'b0;  wr_cycle[18278] = 1'b0;  addr_rom[18278]='h00000000;  wr_data_rom[18278]='h00000000;
    rd_cycle[18279] = 1'b0;  wr_cycle[18279] = 1'b0;  addr_rom[18279]='h00000000;  wr_data_rom[18279]='h00000000;
    rd_cycle[18280] = 1'b0;  wr_cycle[18280] = 1'b0;  addr_rom[18280]='h00000000;  wr_data_rom[18280]='h00000000;
    rd_cycle[18281] = 1'b0;  wr_cycle[18281] = 1'b0;  addr_rom[18281]='h00000000;  wr_data_rom[18281]='h00000000;
    rd_cycle[18282] = 1'b0;  wr_cycle[18282] = 1'b0;  addr_rom[18282]='h00000000;  wr_data_rom[18282]='h00000000;
    rd_cycle[18283] = 1'b0;  wr_cycle[18283] = 1'b0;  addr_rom[18283]='h00000000;  wr_data_rom[18283]='h00000000;
    rd_cycle[18284] = 1'b0;  wr_cycle[18284] = 1'b0;  addr_rom[18284]='h00000000;  wr_data_rom[18284]='h00000000;
    rd_cycle[18285] = 1'b0;  wr_cycle[18285] = 1'b0;  addr_rom[18285]='h00000000;  wr_data_rom[18285]='h00000000;
    rd_cycle[18286] = 1'b0;  wr_cycle[18286] = 1'b0;  addr_rom[18286]='h00000000;  wr_data_rom[18286]='h00000000;
    rd_cycle[18287] = 1'b0;  wr_cycle[18287] = 1'b0;  addr_rom[18287]='h00000000;  wr_data_rom[18287]='h00000000;
    rd_cycle[18288] = 1'b0;  wr_cycle[18288] = 1'b0;  addr_rom[18288]='h00000000;  wr_data_rom[18288]='h00000000;
    rd_cycle[18289] = 1'b0;  wr_cycle[18289] = 1'b0;  addr_rom[18289]='h00000000;  wr_data_rom[18289]='h00000000;
    rd_cycle[18290] = 1'b0;  wr_cycle[18290] = 1'b0;  addr_rom[18290]='h00000000;  wr_data_rom[18290]='h00000000;
    rd_cycle[18291] = 1'b0;  wr_cycle[18291] = 1'b0;  addr_rom[18291]='h00000000;  wr_data_rom[18291]='h00000000;
    rd_cycle[18292] = 1'b0;  wr_cycle[18292] = 1'b0;  addr_rom[18292]='h00000000;  wr_data_rom[18292]='h00000000;
    rd_cycle[18293] = 1'b0;  wr_cycle[18293] = 1'b0;  addr_rom[18293]='h00000000;  wr_data_rom[18293]='h00000000;
    rd_cycle[18294] = 1'b0;  wr_cycle[18294] = 1'b0;  addr_rom[18294]='h00000000;  wr_data_rom[18294]='h00000000;
    rd_cycle[18295] = 1'b0;  wr_cycle[18295] = 1'b0;  addr_rom[18295]='h00000000;  wr_data_rom[18295]='h00000000;
    rd_cycle[18296] = 1'b0;  wr_cycle[18296] = 1'b0;  addr_rom[18296]='h00000000;  wr_data_rom[18296]='h00000000;
    rd_cycle[18297] = 1'b0;  wr_cycle[18297] = 1'b0;  addr_rom[18297]='h00000000;  wr_data_rom[18297]='h00000000;
    rd_cycle[18298] = 1'b0;  wr_cycle[18298] = 1'b0;  addr_rom[18298]='h00000000;  wr_data_rom[18298]='h00000000;
    rd_cycle[18299] = 1'b0;  wr_cycle[18299] = 1'b0;  addr_rom[18299]='h00000000;  wr_data_rom[18299]='h00000000;
    rd_cycle[18300] = 1'b0;  wr_cycle[18300] = 1'b0;  addr_rom[18300]='h00000000;  wr_data_rom[18300]='h00000000;
    rd_cycle[18301] = 1'b0;  wr_cycle[18301] = 1'b0;  addr_rom[18301]='h00000000;  wr_data_rom[18301]='h00000000;
    rd_cycle[18302] = 1'b0;  wr_cycle[18302] = 1'b0;  addr_rom[18302]='h00000000;  wr_data_rom[18302]='h00000000;
    rd_cycle[18303] = 1'b0;  wr_cycle[18303] = 1'b0;  addr_rom[18303]='h00000000;  wr_data_rom[18303]='h00000000;
    rd_cycle[18304] = 1'b0;  wr_cycle[18304] = 1'b0;  addr_rom[18304]='h00000000;  wr_data_rom[18304]='h00000000;
    rd_cycle[18305] = 1'b0;  wr_cycle[18305] = 1'b0;  addr_rom[18305]='h00000000;  wr_data_rom[18305]='h00000000;
    rd_cycle[18306] = 1'b0;  wr_cycle[18306] = 1'b0;  addr_rom[18306]='h00000000;  wr_data_rom[18306]='h00000000;
    rd_cycle[18307] = 1'b0;  wr_cycle[18307] = 1'b0;  addr_rom[18307]='h00000000;  wr_data_rom[18307]='h00000000;
    rd_cycle[18308] = 1'b0;  wr_cycle[18308] = 1'b0;  addr_rom[18308]='h00000000;  wr_data_rom[18308]='h00000000;
    rd_cycle[18309] = 1'b0;  wr_cycle[18309] = 1'b0;  addr_rom[18309]='h00000000;  wr_data_rom[18309]='h00000000;
    rd_cycle[18310] = 1'b0;  wr_cycle[18310] = 1'b0;  addr_rom[18310]='h00000000;  wr_data_rom[18310]='h00000000;
    rd_cycle[18311] = 1'b0;  wr_cycle[18311] = 1'b0;  addr_rom[18311]='h00000000;  wr_data_rom[18311]='h00000000;
    rd_cycle[18312] = 1'b0;  wr_cycle[18312] = 1'b0;  addr_rom[18312]='h00000000;  wr_data_rom[18312]='h00000000;
    rd_cycle[18313] = 1'b0;  wr_cycle[18313] = 1'b0;  addr_rom[18313]='h00000000;  wr_data_rom[18313]='h00000000;
    rd_cycle[18314] = 1'b0;  wr_cycle[18314] = 1'b0;  addr_rom[18314]='h00000000;  wr_data_rom[18314]='h00000000;
    rd_cycle[18315] = 1'b0;  wr_cycle[18315] = 1'b0;  addr_rom[18315]='h00000000;  wr_data_rom[18315]='h00000000;
    rd_cycle[18316] = 1'b0;  wr_cycle[18316] = 1'b0;  addr_rom[18316]='h00000000;  wr_data_rom[18316]='h00000000;
    rd_cycle[18317] = 1'b0;  wr_cycle[18317] = 1'b0;  addr_rom[18317]='h00000000;  wr_data_rom[18317]='h00000000;
    rd_cycle[18318] = 1'b0;  wr_cycle[18318] = 1'b0;  addr_rom[18318]='h00000000;  wr_data_rom[18318]='h00000000;
    rd_cycle[18319] = 1'b0;  wr_cycle[18319] = 1'b0;  addr_rom[18319]='h00000000;  wr_data_rom[18319]='h00000000;
    rd_cycle[18320] = 1'b0;  wr_cycle[18320] = 1'b0;  addr_rom[18320]='h00000000;  wr_data_rom[18320]='h00000000;
    rd_cycle[18321] = 1'b0;  wr_cycle[18321] = 1'b0;  addr_rom[18321]='h00000000;  wr_data_rom[18321]='h00000000;
    rd_cycle[18322] = 1'b0;  wr_cycle[18322] = 1'b0;  addr_rom[18322]='h00000000;  wr_data_rom[18322]='h00000000;
    rd_cycle[18323] = 1'b0;  wr_cycle[18323] = 1'b0;  addr_rom[18323]='h00000000;  wr_data_rom[18323]='h00000000;
    rd_cycle[18324] = 1'b0;  wr_cycle[18324] = 1'b0;  addr_rom[18324]='h00000000;  wr_data_rom[18324]='h00000000;
    rd_cycle[18325] = 1'b0;  wr_cycle[18325] = 1'b0;  addr_rom[18325]='h00000000;  wr_data_rom[18325]='h00000000;
    rd_cycle[18326] = 1'b0;  wr_cycle[18326] = 1'b0;  addr_rom[18326]='h00000000;  wr_data_rom[18326]='h00000000;
    rd_cycle[18327] = 1'b0;  wr_cycle[18327] = 1'b0;  addr_rom[18327]='h00000000;  wr_data_rom[18327]='h00000000;
    rd_cycle[18328] = 1'b0;  wr_cycle[18328] = 1'b0;  addr_rom[18328]='h00000000;  wr_data_rom[18328]='h00000000;
    rd_cycle[18329] = 1'b0;  wr_cycle[18329] = 1'b0;  addr_rom[18329]='h00000000;  wr_data_rom[18329]='h00000000;
    rd_cycle[18330] = 1'b0;  wr_cycle[18330] = 1'b0;  addr_rom[18330]='h00000000;  wr_data_rom[18330]='h00000000;
    rd_cycle[18331] = 1'b0;  wr_cycle[18331] = 1'b0;  addr_rom[18331]='h00000000;  wr_data_rom[18331]='h00000000;
    rd_cycle[18332] = 1'b0;  wr_cycle[18332] = 1'b0;  addr_rom[18332]='h00000000;  wr_data_rom[18332]='h00000000;
    rd_cycle[18333] = 1'b0;  wr_cycle[18333] = 1'b0;  addr_rom[18333]='h00000000;  wr_data_rom[18333]='h00000000;
    rd_cycle[18334] = 1'b0;  wr_cycle[18334] = 1'b0;  addr_rom[18334]='h00000000;  wr_data_rom[18334]='h00000000;
    rd_cycle[18335] = 1'b0;  wr_cycle[18335] = 1'b0;  addr_rom[18335]='h00000000;  wr_data_rom[18335]='h00000000;
    rd_cycle[18336] = 1'b0;  wr_cycle[18336] = 1'b0;  addr_rom[18336]='h00000000;  wr_data_rom[18336]='h00000000;
    rd_cycle[18337] = 1'b0;  wr_cycle[18337] = 1'b0;  addr_rom[18337]='h00000000;  wr_data_rom[18337]='h00000000;
    rd_cycle[18338] = 1'b0;  wr_cycle[18338] = 1'b0;  addr_rom[18338]='h00000000;  wr_data_rom[18338]='h00000000;
    rd_cycle[18339] = 1'b0;  wr_cycle[18339] = 1'b0;  addr_rom[18339]='h00000000;  wr_data_rom[18339]='h00000000;
    rd_cycle[18340] = 1'b0;  wr_cycle[18340] = 1'b0;  addr_rom[18340]='h00000000;  wr_data_rom[18340]='h00000000;
    rd_cycle[18341] = 1'b0;  wr_cycle[18341] = 1'b0;  addr_rom[18341]='h00000000;  wr_data_rom[18341]='h00000000;
    rd_cycle[18342] = 1'b0;  wr_cycle[18342] = 1'b0;  addr_rom[18342]='h00000000;  wr_data_rom[18342]='h00000000;
    rd_cycle[18343] = 1'b0;  wr_cycle[18343] = 1'b0;  addr_rom[18343]='h00000000;  wr_data_rom[18343]='h00000000;
    rd_cycle[18344] = 1'b0;  wr_cycle[18344] = 1'b0;  addr_rom[18344]='h00000000;  wr_data_rom[18344]='h00000000;
    rd_cycle[18345] = 1'b0;  wr_cycle[18345] = 1'b0;  addr_rom[18345]='h00000000;  wr_data_rom[18345]='h00000000;
    rd_cycle[18346] = 1'b0;  wr_cycle[18346] = 1'b0;  addr_rom[18346]='h00000000;  wr_data_rom[18346]='h00000000;
    rd_cycle[18347] = 1'b0;  wr_cycle[18347] = 1'b0;  addr_rom[18347]='h00000000;  wr_data_rom[18347]='h00000000;
    rd_cycle[18348] = 1'b0;  wr_cycle[18348] = 1'b0;  addr_rom[18348]='h00000000;  wr_data_rom[18348]='h00000000;
    rd_cycle[18349] = 1'b0;  wr_cycle[18349] = 1'b0;  addr_rom[18349]='h00000000;  wr_data_rom[18349]='h00000000;
    rd_cycle[18350] = 1'b0;  wr_cycle[18350] = 1'b0;  addr_rom[18350]='h00000000;  wr_data_rom[18350]='h00000000;
    rd_cycle[18351] = 1'b0;  wr_cycle[18351] = 1'b0;  addr_rom[18351]='h00000000;  wr_data_rom[18351]='h00000000;
    rd_cycle[18352] = 1'b0;  wr_cycle[18352] = 1'b0;  addr_rom[18352]='h00000000;  wr_data_rom[18352]='h00000000;
    rd_cycle[18353] = 1'b0;  wr_cycle[18353] = 1'b0;  addr_rom[18353]='h00000000;  wr_data_rom[18353]='h00000000;
    rd_cycle[18354] = 1'b0;  wr_cycle[18354] = 1'b0;  addr_rom[18354]='h00000000;  wr_data_rom[18354]='h00000000;
    rd_cycle[18355] = 1'b0;  wr_cycle[18355] = 1'b0;  addr_rom[18355]='h00000000;  wr_data_rom[18355]='h00000000;
    rd_cycle[18356] = 1'b0;  wr_cycle[18356] = 1'b0;  addr_rom[18356]='h00000000;  wr_data_rom[18356]='h00000000;
    rd_cycle[18357] = 1'b0;  wr_cycle[18357] = 1'b0;  addr_rom[18357]='h00000000;  wr_data_rom[18357]='h00000000;
    rd_cycle[18358] = 1'b0;  wr_cycle[18358] = 1'b0;  addr_rom[18358]='h00000000;  wr_data_rom[18358]='h00000000;
    rd_cycle[18359] = 1'b0;  wr_cycle[18359] = 1'b0;  addr_rom[18359]='h00000000;  wr_data_rom[18359]='h00000000;
    rd_cycle[18360] = 1'b0;  wr_cycle[18360] = 1'b0;  addr_rom[18360]='h00000000;  wr_data_rom[18360]='h00000000;
    rd_cycle[18361] = 1'b0;  wr_cycle[18361] = 1'b0;  addr_rom[18361]='h00000000;  wr_data_rom[18361]='h00000000;
    rd_cycle[18362] = 1'b0;  wr_cycle[18362] = 1'b0;  addr_rom[18362]='h00000000;  wr_data_rom[18362]='h00000000;
    rd_cycle[18363] = 1'b0;  wr_cycle[18363] = 1'b0;  addr_rom[18363]='h00000000;  wr_data_rom[18363]='h00000000;
    rd_cycle[18364] = 1'b0;  wr_cycle[18364] = 1'b0;  addr_rom[18364]='h00000000;  wr_data_rom[18364]='h00000000;
    rd_cycle[18365] = 1'b0;  wr_cycle[18365] = 1'b0;  addr_rom[18365]='h00000000;  wr_data_rom[18365]='h00000000;
    rd_cycle[18366] = 1'b0;  wr_cycle[18366] = 1'b0;  addr_rom[18366]='h00000000;  wr_data_rom[18366]='h00000000;
    rd_cycle[18367] = 1'b0;  wr_cycle[18367] = 1'b0;  addr_rom[18367]='h00000000;  wr_data_rom[18367]='h00000000;
    rd_cycle[18368] = 1'b0;  wr_cycle[18368] = 1'b0;  addr_rom[18368]='h00000000;  wr_data_rom[18368]='h00000000;
    rd_cycle[18369] = 1'b0;  wr_cycle[18369] = 1'b0;  addr_rom[18369]='h00000000;  wr_data_rom[18369]='h00000000;
    rd_cycle[18370] = 1'b0;  wr_cycle[18370] = 1'b0;  addr_rom[18370]='h00000000;  wr_data_rom[18370]='h00000000;
    rd_cycle[18371] = 1'b0;  wr_cycle[18371] = 1'b0;  addr_rom[18371]='h00000000;  wr_data_rom[18371]='h00000000;
    rd_cycle[18372] = 1'b0;  wr_cycle[18372] = 1'b0;  addr_rom[18372]='h00000000;  wr_data_rom[18372]='h00000000;
    rd_cycle[18373] = 1'b0;  wr_cycle[18373] = 1'b0;  addr_rom[18373]='h00000000;  wr_data_rom[18373]='h00000000;
    rd_cycle[18374] = 1'b0;  wr_cycle[18374] = 1'b0;  addr_rom[18374]='h00000000;  wr_data_rom[18374]='h00000000;
    rd_cycle[18375] = 1'b0;  wr_cycle[18375] = 1'b0;  addr_rom[18375]='h00000000;  wr_data_rom[18375]='h00000000;
    rd_cycle[18376] = 1'b0;  wr_cycle[18376] = 1'b0;  addr_rom[18376]='h00000000;  wr_data_rom[18376]='h00000000;
    rd_cycle[18377] = 1'b0;  wr_cycle[18377] = 1'b0;  addr_rom[18377]='h00000000;  wr_data_rom[18377]='h00000000;
    rd_cycle[18378] = 1'b0;  wr_cycle[18378] = 1'b0;  addr_rom[18378]='h00000000;  wr_data_rom[18378]='h00000000;
    rd_cycle[18379] = 1'b0;  wr_cycle[18379] = 1'b0;  addr_rom[18379]='h00000000;  wr_data_rom[18379]='h00000000;
    rd_cycle[18380] = 1'b0;  wr_cycle[18380] = 1'b0;  addr_rom[18380]='h00000000;  wr_data_rom[18380]='h00000000;
    rd_cycle[18381] = 1'b0;  wr_cycle[18381] = 1'b0;  addr_rom[18381]='h00000000;  wr_data_rom[18381]='h00000000;
    rd_cycle[18382] = 1'b0;  wr_cycle[18382] = 1'b0;  addr_rom[18382]='h00000000;  wr_data_rom[18382]='h00000000;
    rd_cycle[18383] = 1'b0;  wr_cycle[18383] = 1'b0;  addr_rom[18383]='h00000000;  wr_data_rom[18383]='h00000000;
    rd_cycle[18384] = 1'b0;  wr_cycle[18384] = 1'b0;  addr_rom[18384]='h00000000;  wr_data_rom[18384]='h00000000;
    rd_cycle[18385] = 1'b0;  wr_cycle[18385] = 1'b0;  addr_rom[18385]='h00000000;  wr_data_rom[18385]='h00000000;
    rd_cycle[18386] = 1'b0;  wr_cycle[18386] = 1'b0;  addr_rom[18386]='h00000000;  wr_data_rom[18386]='h00000000;
    rd_cycle[18387] = 1'b0;  wr_cycle[18387] = 1'b0;  addr_rom[18387]='h00000000;  wr_data_rom[18387]='h00000000;
    rd_cycle[18388] = 1'b0;  wr_cycle[18388] = 1'b0;  addr_rom[18388]='h00000000;  wr_data_rom[18388]='h00000000;
    rd_cycle[18389] = 1'b0;  wr_cycle[18389] = 1'b0;  addr_rom[18389]='h00000000;  wr_data_rom[18389]='h00000000;
    rd_cycle[18390] = 1'b0;  wr_cycle[18390] = 1'b0;  addr_rom[18390]='h00000000;  wr_data_rom[18390]='h00000000;
    rd_cycle[18391] = 1'b0;  wr_cycle[18391] = 1'b0;  addr_rom[18391]='h00000000;  wr_data_rom[18391]='h00000000;
    rd_cycle[18392] = 1'b0;  wr_cycle[18392] = 1'b0;  addr_rom[18392]='h00000000;  wr_data_rom[18392]='h00000000;
    rd_cycle[18393] = 1'b0;  wr_cycle[18393] = 1'b0;  addr_rom[18393]='h00000000;  wr_data_rom[18393]='h00000000;
    rd_cycle[18394] = 1'b0;  wr_cycle[18394] = 1'b0;  addr_rom[18394]='h00000000;  wr_data_rom[18394]='h00000000;
    rd_cycle[18395] = 1'b0;  wr_cycle[18395] = 1'b0;  addr_rom[18395]='h00000000;  wr_data_rom[18395]='h00000000;
    rd_cycle[18396] = 1'b0;  wr_cycle[18396] = 1'b0;  addr_rom[18396]='h00000000;  wr_data_rom[18396]='h00000000;
    rd_cycle[18397] = 1'b0;  wr_cycle[18397] = 1'b0;  addr_rom[18397]='h00000000;  wr_data_rom[18397]='h00000000;
    rd_cycle[18398] = 1'b0;  wr_cycle[18398] = 1'b0;  addr_rom[18398]='h00000000;  wr_data_rom[18398]='h00000000;
    rd_cycle[18399] = 1'b0;  wr_cycle[18399] = 1'b0;  addr_rom[18399]='h00000000;  wr_data_rom[18399]='h00000000;
    rd_cycle[18400] = 1'b0;  wr_cycle[18400] = 1'b0;  addr_rom[18400]='h00000000;  wr_data_rom[18400]='h00000000;
    rd_cycle[18401] = 1'b0;  wr_cycle[18401] = 1'b0;  addr_rom[18401]='h00000000;  wr_data_rom[18401]='h00000000;
    rd_cycle[18402] = 1'b0;  wr_cycle[18402] = 1'b0;  addr_rom[18402]='h00000000;  wr_data_rom[18402]='h00000000;
    rd_cycle[18403] = 1'b0;  wr_cycle[18403] = 1'b0;  addr_rom[18403]='h00000000;  wr_data_rom[18403]='h00000000;
    rd_cycle[18404] = 1'b0;  wr_cycle[18404] = 1'b0;  addr_rom[18404]='h00000000;  wr_data_rom[18404]='h00000000;
    rd_cycle[18405] = 1'b0;  wr_cycle[18405] = 1'b0;  addr_rom[18405]='h00000000;  wr_data_rom[18405]='h00000000;
    rd_cycle[18406] = 1'b0;  wr_cycle[18406] = 1'b0;  addr_rom[18406]='h00000000;  wr_data_rom[18406]='h00000000;
    rd_cycle[18407] = 1'b0;  wr_cycle[18407] = 1'b0;  addr_rom[18407]='h00000000;  wr_data_rom[18407]='h00000000;
    rd_cycle[18408] = 1'b0;  wr_cycle[18408] = 1'b0;  addr_rom[18408]='h00000000;  wr_data_rom[18408]='h00000000;
    rd_cycle[18409] = 1'b0;  wr_cycle[18409] = 1'b0;  addr_rom[18409]='h00000000;  wr_data_rom[18409]='h00000000;
    rd_cycle[18410] = 1'b0;  wr_cycle[18410] = 1'b0;  addr_rom[18410]='h00000000;  wr_data_rom[18410]='h00000000;
    rd_cycle[18411] = 1'b0;  wr_cycle[18411] = 1'b0;  addr_rom[18411]='h00000000;  wr_data_rom[18411]='h00000000;
    rd_cycle[18412] = 1'b0;  wr_cycle[18412] = 1'b0;  addr_rom[18412]='h00000000;  wr_data_rom[18412]='h00000000;
    rd_cycle[18413] = 1'b0;  wr_cycle[18413] = 1'b0;  addr_rom[18413]='h00000000;  wr_data_rom[18413]='h00000000;
    rd_cycle[18414] = 1'b0;  wr_cycle[18414] = 1'b0;  addr_rom[18414]='h00000000;  wr_data_rom[18414]='h00000000;
    rd_cycle[18415] = 1'b0;  wr_cycle[18415] = 1'b0;  addr_rom[18415]='h00000000;  wr_data_rom[18415]='h00000000;
    rd_cycle[18416] = 1'b0;  wr_cycle[18416] = 1'b0;  addr_rom[18416]='h00000000;  wr_data_rom[18416]='h00000000;
    rd_cycle[18417] = 1'b0;  wr_cycle[18417] = 1'b0;  addr_rom[18417]='h00000000;  wr_data_rom[18417]='h00000000;
    rd_cycle[18418] = 1'b0;  wr_cycle[18418] = 1'b0;  addr_rom[18418]='h00000000;  wr_data_rom[18418]='h00000000;
    rd_cycle[18419] = 1'b0;  wr_cycle[18419] = 1'b0;  addr_rom[18419]='h00000000;  wr_data_rom[18419]='h00000000;
    rd_cycle[18420] = 1'b0;  wr_cycle[18420] = 1'b0;  addr_rom[18420]='h00000000;  wr_data_rom[18420]='h00000000;
    rd_cycle[18421] = 1'b0;  wr_cycle[18421] = 1'b0;  addr_rom[18421]='h00000000;  wr_data_rom[18421]='h00000000;
    rd_cycle[18422] = 1'b0;  wr_cycle[18422] = 1'b0;  addr_rom[18422]='h00000000;  wr_data_rom[18422]='h00000000;
    rd_cycle[18423] = 1'b0;  wr_cycle[18423] = 1'b0;  addr_rom[18423]='h00000000;  wr_data_rom[18423]='h00000000;
    rd_cycle[18424] = 1'b0;  wr_cycle[18424] = 1'b0;  addr_rom[18424]='h00000000;  wr_data_rom[18424]='h00000000;
    rd_cycle[18425] = 1'b0;  wr_cycle[18425] = 1'b0;  addr_rom[18425]='h00000000;  wr_data_rom[18425]='h00000000;
    rd_cycle[18426] = 1'b0;  wr_cycle[18426] = 1'b0;  addr_rom[18426]='h00000000;  wr_data_rom[18426]='h00000000;
    rd_cycle[18427] = 1'b0;  wr_cycle[18427] = 1'b0;  addr_rom[18427]='h00000000;  wr_data_rom[18427]='h00000000;
    rd_cycle[18428] = 1'b0;  wr_cycle[18428] = 1'b0;  addr_rom[18428]='h00000000;  wr_data_rom[18428]='h00000000;
    rd_cycle[18429] = 1'b0;  wr_cycle[18429] = 1'b0;  addr_rom[18429]='h00000000;  wr_data_rom[18429]='h00000000;
    rd_cycle[18430] = 1'b0;  wr_cycle[18430] = 1'b0;  addr_rom[18430]='h00000000;  wr_data_rom[18430]='h00000000;
    rd_cycle[18431] = 1'b0;  wr_cycle[18431] = 1'b0;  addr_rom[18431]='h00000000;  wr_data_rom[18431]='h00000000;
    rd_cycle[18432] = 1'b0;  wr_cycle[18432] = 1'b0;  addr_rom[18432]='h00000000;  wr_data_rom[18432]='h00000000;
    rd_cycle[18433] = 1'b0;  wr_cycle[18433] = 1'b0;  addr_rom[18433]='h00000000;  wr_data_rom[18433]='h00000000;
    rd_cycle[18434] = 1'b0;  wr_cycle[18434] = 1'b0;  addr_rom[18434]='h00000000;  wr_data_rom[18434]='h00000000;
    rd_cycle[18435] = 1'b0;  wr_cycle[18435] = 1'b0;  addr_rom[18435]='h00000000;  wr_data_rom[18435]='h00000000;
    rd_cycle[18436] = 1'b0;  wr_cycle[18436] = 1'b0;  addr_rom[18436]='h00000000;  wr_data_rom[18436]='h00000000;
    rd_cycle[18437] = 1'b0;  wr_cycle[18437] = 1'b0;  addr_rom[18437]='h00000000;  wr_data_rom[18437]='h00000000;
    rd_cycle[18438] = 1'b0;  wr_cycle[18438] = 1'b0;  addr_rom[18438]='h00000000;  wr_data_rom[18438]='h00000000;
    rd_cycle[18439] = 1'b0;  wr_cycle[18439] = 1'b0;  addr_rom[18439]='h00000000;  wr_data_rom[18439]='h00000000;
    rd_cycle[18440] = 1'b0;  wr_cycle[18440] = 1'b0;  addr_rom[18440]='h00000000;  wr_data_rom[18440]='h00000000;
    rd_cycle[18441] = 1'b0;  wr_cycle[18441] = 1'b0;  addr_rom[18441]='h00000000;  wr_data_rom[18441]='h00000000;
    rd_cycle[18442] = 1'b0;  wr_cycle[18442] = 1'b0;  addr_rom[18442]='h00000000;  wr_data_rom[18442]='h00000000;
    rd_cycle[18443] = 1'b0;  wr_cycle[18443] = 1'b0;  addr_rom[18443]='h00000000;  wr_data_rom[18443]='h00000000;
    rd_cycle[18444] = 1'b0;  wr_cycle[18444] = 1'b0;  addr_rom[18444]='h00000000;  wr_data_rom[18444]='h00000000;
    rd_cycle[18445] = 1'b0;  wr_cycle[18445] = 1'b0;  addr_rom[18445]='h00000000;  wr_data_rom[18445]='h00000000;
    rd_cycle[18446] = 1'b0;  wr_cycle[18446] = 1'b0;  addr_rom[18446]='h00000000;  wr_data_rom[18446]='h00000000;
    rd_cycle[18447] = 1'b0;  wr_cycle[18447] = 1'b0;  addr_rom[18447]='h00000000;  wr_data_rom[18447]='h00000000;
    rd_cycle[18448] = 1'b0;  wr_cycle[18448] = 1'b0;  addr_rom[18448]='h00000000;  wr_data_rom[18448]='h00000000;
    rd_cycle[18449] = 1'b0;  wr_cycle[18449] = 1'b0;  addr_rom[18449]='h00000000;  wr_data_rom[18449]='h00000000;
    rd_cycle[18450] = 1'b0;  wr_cycle[18450] = 1'b0;  addr_rom[18450]='h00000000;  wr_data_rom[18450]='h00000000;
    rd_cycle[18451] = 1'b0;  wr_cycle[18451] = 1'b0;  addr_rom[18451]='h00000000;  wr_data_rom[18451]='h00000000;
    rd_cycle[18452] = 1'b0;  wr_cycle[18452] = 1'b0;  addr_rom[18452]='h00000000;  wr_data_rom[18452]='h00000000;
    rd_cycle[18453] = 1'b0;  wr_cycle[18453] = 1'b0;  addr_rom[18453]='h00000000;  wr_data_rom[18453]='h00000000;
    rd_cycle[18454] = 1'b0;  wr_cycle[18454] = 1'b0;  addr_rom[18454]='h00000000;  wr_data_rom[18454]='h00000000;
    rd_cycle[18455] = 1'b0;  wr_cycle[18455] = 1'b0;  addr_rom[18455]='h00000000;  wr_data_rom[18455]='h00000000;
    rd_cycle[18456] = 1'b0;  wr_cycle[18456] = 1'b0;  addr_rom[18456]='h00000000;  wr_data_rom[18456]='h00000000;
    rd_cycle[18457] = 1'b0;  wr_cycle[18457] = 1'b0;  addr_rom[18457]='h00000000;  wr_data_rom[18457]='h00000000;
    rd_cycle[18458] = 1'b0;  wr_cycle[18458] = 1'b0;  addr_rom[18458]='h00000000;  wr_data_rom[18458]='h00000000;
    rd_cycle[18459] = 1'b0;  wr_cycle[18459] = 1'b0;  addr_rom[18459]='h00000000;  wr_data_rom[18459]='h00000000;
    rd_cycle[18460] = 1'b0;  wr_cycle[18460] = 1'b0;  addr_rom[18460]='h00000000;  wr_data_rom[18460]='h00000000;
    rd_cycle[18461] = 1'b0;  wr_cycle[18461] = 1'b0;  addr_rom[18461]='h00000000;  wr_data_rom[18461]='h00000000;
    rd_cycle[18462] = 1'b0;  wr_cycle[18462] = 1'b0;  addr_rom[18462]='h00000000;  wr_data_rom[18462]='h00000000;
    rd_cycle[18463] = 1'b0;  wr_cycle[18463] = 1'b0;  addr_rom[18463]='h00000000;  wr_data_rom[18463]='h00000000;
    rd_cycle[18464] = 1'b0;  wr_cycle[18464] = 1'b0;  addr_rom[18464]='h00000000;  wr_data_rom[18464]='h00000000;
    rd_cycle[18465] = 1'b0;  wr_cycle[18465] = 1'b0;  addr_rom[18465]='h00000000;  wr_data_rom[18465]='h00000000;
    rd_cycle[18466] = 1'b0;  wr_cycle[18466] = 1'b0;  addr_rom[18466]='h00000000;  wr_data_rom[18466]='h00000000;
    rd_cycle[18467] = 1'b0;  wr_cycle[18467] = 1'b0;  addr_rom[18467]='h00000000;  wr_data_rom[18467]='h00000000;
    rd_cycle[18468] = 1'b0;  wr_cycle[18468] = 1'b0;  addr_rom[18468]='h00000000;  wr_data_rom[18468]='h00000000;
    rd_cycle[18469] = 1'b0;  wr_cycle[18469] = 1'b0;  addr_rom[18469]='h00000000;  wr_data_rom[18469]='h00000000;
    rd_cycle[18470] = 1'b0;  wr_cycle[18470] = 1'b0;  addr_rom[18470]='h00000000;  wr_data_rom[18470]='h00000000;
    rd_cycle[18471] = 1'b0;  wr_cycle[18471] = 1'b0;  addr_rom[18471]='h00000000;  wr_data_rom[18471]='h00000000;
    rd_cycle[18472] = 1'b0;  wr_cycle[18472] = 1'b0;  addr_rom[18472]='h00000000;  wr_data_rom[18472]='h00000000;
    rd_cycle[18473] = 1'b0;  wr_cycle[18473] = 1'b0;  addr_rom[18473]='h00000000;  wr_data_rom[18473]='h00000000;
    rd_cycle[18474] = 1'b0;  wr_cycle[18474] = 1'b0;  addr_rom[18474]='h00000000;  wr_data_rom[18474]='h00000000;
    rd_cycle[18475] = 1'b0;  wr_cycle[18475] = 1'b0;  addr_rom[18475]='h00000000;  wr_data_rom[18475]='h00000000;
    rd_cycle[18476] = 1'b0;  wr_cycle[18476] = 1'b0;  addr_rom[18476]='h00000000;  wr_data_rom[18476]='h00000000;
    rd_cycle[18477] = 1'b0;  wr_cycle[18477] = 1'b0;  addr_rom[18477]='h00000000;  wr_data_rom[18477]='h00000000;
    rd_cycle[18478] = 1'b0;  wr_cycle[18478] = 1'b0;  addr_rom[18478]='h00000000;  wr_data_rom[18478]='h00000000;
    rd_cycle[18479] = 1'b0;  wr_cycle[18479] = 1'b0;  addr_rom[18479]='h00000000;  wr_data_rom[18479]='h00000000;
    rd_cycle[18480] = 1'b0;  wr_cycle[18480] = 1'b0;  addr_rom[18480]='h00000000;  wr_data_rom[18480]='h00000000;
    rd_cycle[18481] = 1'b0;  wr_cycle[18481] = 1'b0;  addr_rom[18481]='h00000000;  wr_data_rom[18481]='h00000000;
    rd_cycle[18482] = 1'b0;  wr_cycle[18482] = 1'b0;  addr_rom[18482]='h00000000;  wr_data_rom[18482]='h00000000;
    rd_cycle[18483] = 1'b0;  wr_cycle[18483] = 1'b0;  addr_rom[18483]='h00000000;  wr_data_rom[18483]='h00000000;
    rd_cycle[18484] = 1'b0;  wr_cycle[18484] = 1'b0;  addr_rom[18484]='h00000000;  wr_data_rom[18484]='h00000000;
    rd_cycle[18485] = 1'b0;  wr_cycle[18485] = 1'b0;  addr_rom[18485]='h00000000;  wr_data_rom[18485]='h00000000;
    rd_cycle[18486] = 1'b0;  wr_cycle[18486] = 1'b0;  addr_rom[18486]='h00000000;  wr_data_rom[18486]='h00000000;
    rd_cycle[18487] = 1'b0;  wr_cycle[18487] = 1'b0;  addr_rom[18487]='h00000000;  wr_data_rom[18487]='h00000000;
    rd_cycle[18488] = 1'b0;  wr_cycle[18488] = 1'b0;  addr_rom[18488]='h00000000;  wr_data_rom[18488]='h00000000;
    rd_cycle[18489] = 1'b0;  wr_cycle[18489] = 1'b0;  addr_rom[18489]='h00000000;  wr_data_rom[18489]='h00000000;
    rd_cycle[18490] = 1'b0;  wr_cycle[18490] = 1'b0;  addr_rom[18490]='h00000000;  wr_data_rom[18490]='h00000000;
    rd_cycle[18491] = 1'b0;  wr_cycle[18491] = 1'b0;  addr_rom[18491]='h00000000;  wr_data_rom[18491]='h00000000;
    rd_cycle[18492] = 1'b0;  wr_cycle[18492] = 1'b0;  addr_rom[18492]='h00000000;  wr_data_rom[18492]='h00000000;
    rd_cycle[18493] = 1'b0;  wr_cycle[18493] = 1'b0;  addr_rom[18493]='h00000000;  wr_data_rom[18493]='h00000000;
    rd_cycle[18494] = 1'b0;  wr_cycle[18494] = 1'b0;  addr_rom[18494]='h00000000;  wr_data_rom[18494]='h00000000;
    rd_cycle[18495] = 1'b0;  wr_cycle[18495] = 1'b0;  addr_rom[18495]='h00000000;  wr_data_rom[18495]='h00000000;
    rd_cycle[18496] = 1'b0;  wr_cycle[18496] = 1'b0;  addr_rom[18496]='h00000000;  wr_data_rom[18496]='h00000000;
    rd_cycle[18497] = 1'b0;  wr_cycle[18497] = 1'b0;  addr_rom[18497]='h00000000;  wr_data_rom[18497]='h00000000;
    rd_cycle[18498] = 1'b0;  wr_cycle[18498] = 1'b0;  addr_rom[18498]='h00000000;  wr_data_rom[18498]='h00000000;
    rd_cycle[18499] = 1'b0;  wr_cycle[18499] = 1'b0;  addr_rom[18499]='h00000000;  wr_data_rom[18499]='h00000000;
    rd_cycle[18500] = 1'b0;  wr_cycle[18500] = 1'b0;  addr_rom[18500]='h00000000;  wr_data_rom[18500]='h00000000;
    rd_cycle[18501] = 1'b0;  wr_cycle[18501] = 1'b0;  addr_rom[18501]='h00000000;  wr_data_rom[18501]='h00000000;
    rd_cycle[18502] = 1'b0;  wr_cycle[18502] = 1'b0;  addr_rom[18502]='h00000000;  wr_data_rom[18502]='h00000000;
    rd_cycle[18503] = 1'b0;  wr_cycle[18503] = 1'b0;  addr_rom[18503]='h00000000;  wr_data_rom[18503]='h00000000;
    rd_cycle[18504] = 1'b0;  wr_cycle[18504] = 1'b0;  addr_rom[18504]='h00000000;  wr_data_rom[18504]='h00000000;
    rd_cycle[18505] = 1'b0;  wr_cycle[18505] = 1'b0;  addr_rom[18505]='h00000000;  wr_data_rom[18505]='h00000000;
    rd_cycle[18506] = 1'b0;  wr_cycle[18506] = 1'b0;  addr_rom[18506]='h00000000;  wr_data_rom[18506]='h00000000;
    rd_cycle[18507] = 1'b0;  wr_cycle[18507] = 1'b0;  addr_rom[18507]='h00000000;  wr_data_rom[18507]='h00000000;
    rd_cycle[18508] = 1'b0;  wr_cycle[18508] = 1'b0;  addr_rom[18508]='h00000000;  wr_data_rom[18508]='h00000000;
    rd_cycle[18509] = 1'b0;  wr_cycle[18509] = 1'b0;  addr_rom[18509]='h00000000;  wr_data_rom[18509]='h00000000;
    rd_cycle[18510] = 1'b0;  wr_cycle[18510] = 1'b0;  addr_rom[18510]='h00000000;  wr_data_rom[18510]='h00000000;
    rd_cycle[18511] = 1'b0;  wr_cycle[18511] = 1'b0;  addr_rom[18511]='h00000000;  wr_data_rom[18511]='h00000000;
    rd_cycle[18512] = 1'b0;  wr_cycle[18512] = 1'b0;  addr_rom[18512]='h00000000;  wr_data_rom[18512]='h00000000;
    rd_cycle[18513] = 1'b0;  wr_cycle[18513] = 1'b0;  addr_rom[18513]='h00000000;  wr_data_rom[18513]='h00000000;
    rd_cycle[18514] = 1'b0;  wr_cycle[18514] = 1'b0;  addr_rom[18514]='h00000000;  wr_data_rom[18514]='h00000000;
    rd_cycle[18515] = 1'b0;  wr_cycle[18515] = 1'b0;  addr_rom[18515]='h00000000;  wr_data_rom[18515]='h00000000;
    rd_cycle[18516] = 1'b0;  wr_cycle[18516] = 1'b0;  addr_rom[18516]='h00000000;  wr_data_rom[18516]='h00000000;
    rd_cycle[18517] = 1'b0;  wr_cycle[18517] = 1'b0;  addr_rom[18517]='h00000000;  wr_data_rom[18517]='h00000000;
    rd_cycle[18518] = 1'b0;  wr_cycle[18518] = 1'b0;  addr_rom[18518]='h00000000;  wr_data_rom[18518]='h00000000;
    rd_cycle[18519] = 1'b0;  wr_cycle[18519] = 1'b0;  addr_rom[18519]='h00000000;  wr_data_rom[18519]='h00000000;
    rd_cycle[18520] = 1'b0;  wr_cycle[18520] = 1'b0;  addr_rom[18520]='h00000000;  wr_data_rom[18520]='h00000000;
    rd_cycle[18521] = 1'b0;  wr_cycle[18521] = 1'b0;  addr_rom[18521]='h00000000;  wr_data_rom[18521]='h00000000;
    rd_cycle[18522] = 1'b0;  wr_cycle[18522] = 1'b0;  addr_rom[18522]='h00000000;  wr_data_rom[18522]='h00000000;
    rd_cycle[18523] = 1'b0;  wr_cycle[18523] = 1'b0;  addr_rom[18523]='h00000000;  wr_data_rom[18523]='h00000000;
    rd_cycle[18524] = 1'b0;  wr_cycle[18524] = 1'b0;  addr_rom[18524]='h00000000;  wr_data_rom[18524]='h00000000;
    rd_cycle[18525] = 1'b0;  wr_cycle[18525] = 1'b0;  addr_rom[18525]='h00000000;  wr_data_rom[18525]='h00000000;
    rd_cycle[18526] = 1'b0;  wr_cycle[18526] = 1'b0;  addr_rom[18526]='h00000000;  wr_data_rom[18526]='h00000000;
    rd_cycle[18527] = 1'b0;  wr_cycle[18527] = 1'b0;  addr_rom[18527]='h00000000;  wr_data_rom[18527]='h00000000;
    rd_cycle[18528] = 1'b0;  wr_cycle[18528] = 1'b0;  addr_rom[18528]='h00000000;  wr_data_rom[18528]='h00000000;
    rd_cycle[18529] = 1'b0;  wr_cycle[18529] = 1'b0;  addr_rom[18529]='h00000000;  wr_data_rom[18529]='h00000000;
    rd_cycle[18530] = 1'b0;  wr_cycle[18530] = 1'b0;  addr_rom[18530]='h00000000;  wr_data_rom[18530]='h00000000;
    rd_cycle[18531] = 1'b0;  wr_cycle[18531] = 1'b0;  addr_rom[18531]='h00000000;  wr_data_rom[18531]='h00000000;
    rd_cycle[18532] = 1'b0;  wr_cycle[18532] = 1'b0;  addr_rom[18532]='h00000000;  wr_data_rom[18532]='h00000000;
    rd_cycle[18533] = 1'b0;  wr_cycle[18533] = 1'b0;  addr_rom[18533]='h00000000;  wr_data_rom[18533]='h00000000;
    rd_cycle[18534] = 1'b0;  wr_cycle[18534] = 1'b0;  addr_rom[18534]='h00000000;  wr_data_rom[18534]='h00000000;
    rd_cycle[18535] = 1'b0;  wr_cycle[18535] = 1'b0;  addr_rom[18535]='h00000000;  wr_data_rom[18535]='h00000000;
    rd_cycle[18536] = 1'b0;  wr_cycle[18536] = 1'b0;  addr_rom[18536]='h00000000;  wr_data_rom[18536]='h00000000;
    rd_cycle[18537] = 1'b0;  wr_cycle[18537] = 1'b0;  addr_rom[18537]='h00000000;  wr_data_rom[18537]='h00000000;
    rd_cycle[18538] = 1'b0;  wr_cycle[18538] = 1'b0;  addr_rom[18538]='h00000000;  wr_data_rom[18538]='h00000000;
    rd_cycle[18539] = 1'b0;  wr_cycle[18539] = 1'b0;  addr_rom[18539]='h00000000;  wr_data_rom[18539]='h00000000;
    rd_cycle[18540] = 1'b0;  wr_cycle[18540] = 1'b0;  addr_rom[18540]='h00000000;  wr_data_rom[18540]='h00000000;
    rd_cycle[18541] = 1'b0;  wr_cycle[18541] = 1'b0;  addr_rom[18541]='h00000000;  wr_data_rom[18541]='h00000000;
    rd_cycle[18542] = 1'b0;  wr_cycle[18542] = 1'b0;  addr_rom[18542]='h00000000;  wr_data_rom[18542]='h00000000;
    rd_cycle[18543] = 1'b0;  wr_cycle[18543] = 1'b0;  addr_rom[18543]='h00000000;  wr_data_rom[18543]='h00000000;
    rd_cycle[18544] = 1'b0;  wr_cycle[18544] = 1'b0;  addr_rom[18544]='h00000000;  wr_data_rom[18544]='h00000000;
    rd_cycle[18545] = 1'b0;  wr_cycle[18545] = 1'b0;  addr_rom[18545]='h00000000;  wr_data_rom[18545]='h00000000;
    rd_cycle[18546] = 1'b0;  wr_cycle[18546] = 1'b0;  addr_rom[18546]='h00000000;  wr_data_rom[18546]='h00000000;
    rd_cycle[18547] = 1'b0;  wr_cycle[18547] = 1'b0;  addr_rom[18547]='h00000000;  wr_data_rom[18547]='h00000000;
    rd_cycle[18548] = 1'b0;  wr_cycle[18548] = 1'b0;  addr_rom[18548]='h00000000;  wr_data_rom[18548]='h00000000;
    rd_cycle[18549] = 1'b0;  wr_cycle[18549] = 1'b0;  addr_rom[18549]='h00000000;  wr_data_rom[18549]='h00000000;
    rd_cycle[18550] = 1'b0;  wr_cycle[18550] = 1'b0;  addr_rom[18550]='h00000000;  wr_data_rom[18550]='h00000000;
    rd_cycle[18551] = 1'b0;  wr_cycle[18551] = 1'b0;  addr_rom[18551]='h00000000;  wr_data_rom[18551]='h00000000;
    rd_cycle[18552] = 1'b0;  wr_cycle[18552] = 1'b0;  addr_rom[18552]='h00000000;  wr_data_rom[18552]='h00000000;
    rd_cycle[18553] = 1'b0;  wr_cycle[18553] = 1'b0;  addr_rom[18553]='h00000000;  wr_data_rom[18553]='h00000000;
    rd_cycle[18554] = 1'b0;  wr_cycle[18554] = 1'b0;  addr_rom[18554]='h00000000;  wr_data_rom[18554]='h00000000;
    rd_cycle[18555] = 1'b0;  wr_cycle[18555] = 1'b0;  addr_rom[18555]='h00000000;  wr_data_rom[18555]='h00000000;
    rd_cycle[18556] = 1'b0;  wr_cycle[18556] = 1'b0;  addr_rom[18556]='h00000000;  wr_data_rom[18556]='h00000000;
    rd_cycle[18557] = 1'b0;  wr_cycle[18557] = 1'b0;  addr_rom[18557]='h00000000;  wr_data_rom[18557]='h00000000;
    rd_cycle[18558] = 1'b0;  wr_cycle[18558] = 1'b0;  addr_rom[18558]='h00000000;  wr_data_rom[18558]='h00000000;
    rd_cycle[18559] = 1'b0;  wr_cycle[18559] = 1'b0;  addr_rom[18559]='h00000000;  wr_data_rom[18559]='h00000000;
    rd_cycle[18560] = 1'b0;  wr_cycle[18560] = 1'b0;  addr_rom[18560]='h00000000;  wr_data_rom[18560]='h00000000;
    rd_cycle[18561] = 1'b0;  wr_cycle[18561] = 1'b0;  addr_rom[18561]='h00000000;  wr_data_rom[18561]='h00000000;
    rd_cycle[18562] = 1'b0;  wr_cycle[18562] = 1'b0;  addr_rom[18562]='h00000000;  wr_data_rom[18562]='h00000000;
    rd_cycle[18563] = 1'b0;  wr_cycle[18563] = 1'b0;  addr_rom[18563]='h00000000;  wr_data_rom[18563]='h00000000;
    rd_cycle[18564] = 1'b0;  wr_cycle[18564] = 1'b0;  addr_rom[18564]='h00000000;  wr_data_rom[18564]='h00000000;
    rd_cycle[18565] = 1'b0;  wr_cycle[18565] = 1'b0;  addr_rom[18565]='h00000000;  wr_data_rom[18565]='h00000000;
    rd_cycle[18566] = 1'b0;  wr_cycle[18566] = 1'b0;  addr_rom[18566]='h00000000;  wr_data_rom[18566]='h00000000;
    rd_cycle[18567] = 1'b0;  wr_cycle[18567] = 1'b0;  addr_rom[18567]='h00000000;  wr_data_rom[18567]='h00000000;
    rd_cycle[18568] = 1'b0;  wr_cycle[18568] = 1'b0;  addr_rom[18568]='h00000000;  wr_data_rom[18568]='h00000000;
    rd_cycle[18569] = 1'b0;  wr_cycle[18569] = 1'b0;  addr_rom[18569]='h00000000;  wr_data_rom[18569]='h00000000;
    rd_cycle[18570] = 1'b0;  wr_cycle[18570] = 1'b0;  addr_rom[18570]='h00000000;  wr_data_rom[18570]='h00000000;
    rd_cycle[18571] = 1'b0;  wr_cycle[18571] = 1'b0;  addr_rom[18571]='h00000000;  wr_data_rom[18571]='h00000000;
    rd_cycle[18572] = 1'b0;  wr_cycle[18572] = 1'b0;  addr_rom[18572]='h00000000;  wr_data_rom[18572]='h00000000;
    rd_cycle[18573] = 1'b0;  wr_cycle[18573] = 1'b0;  addr_rom[18573]='h00000000;  wr_data_rom[18573]='h00000000;
    rd_cycle[18574] = 1'b0;  wr_cycle[18574] = 1'b0;  addr_rom[18574]='h00000000;  wr_data_rom[18574]='h00000000;
    rd_cycle[18575] = 1'b0;  wr_cycle[18575] = 1'b0;  addr_rom[18575]='h00000000;  wr_data_rom[18575]='h00000000;
    rd_cycle[18576] = 1'b0;  wr_cycle[18576] = 1'b0;  addr_rom[18576]='h00000000;  wr_data_rom[18576]='h00000000;
    rd_cycle[18577] = 1'b0;  wr_cycle[18577] = 1'b0;  addr_rom[18577]='h00000000;  wr_data_rom[18577]='h00000000;
    rd_cycle[18578] = 1'b0;  wr_cycle[18578] = 1'b0;  addr_rom[18578]='h00000000;  wr_data_rom[18578]='h00000000;
    rd_cycle[18579] = 1'b0;  wr_cycle[18579] = 1'b0;  addr_rom[18579]='h00000000;  wr_data_rom[18579]='h00000000;
    rd_cycle[18580] = 1'b0;  wr_cycle[18580] = 1'b0;  addr_rom[18580]='h00000000;  wr_data_rom[18580]='h00000000;
    rd_cycle[18581] = 1'b0;  wr_cycle[18581] = 1'b0;  addr_rom[18581]='h00000000;  wr_data_rom[18581]='h00000000;
    rd_cycle[18582] = 1'b0;  wr_cycle[18582] = 1'b0;  addr_rom[18582]='h00000000;  wr_data_rom[18582]='h00000000;
    rd_cycle[18583] = 1'b0;  wr_cycle[18583] = 1'b0;  addr_rom[18583]='h00000000;  wr_data_rom[18583]='h00000000;
    rd_cycle[18584] = 1'b0;  wr_cycle[18584] = 1'b0;  addr_rom[18584]='h00000000;  wr_data_rom[18584]='h00000000;
    rd_cycle[18585] = 1'b0;  wr_cycle[18585] = 1'b0;  addr_rom[18585]='h00000000;  wr_data_rom[18585]='h00000000;
    rd_cycle[18586] = 1'b0;  wr_cycle[18586] = 1'b0;  addr_rom[18586]='h00000000;  wr_data_rom[18586]='h00000000;
    rd_cycle[18587] = 1'b0;  wr_cycle[18587] = 1'b0;  addr_rom[18587]='h00000000;  wr_data_rom[18587]='h00000000;
    rd_cycle[18588] = 1'b0;  wr_cycle[18588] = 1'b0;  addr_rom[18588]='h00000000;  wr_data_rom[18588]='h00000000;
    rd_cycle[18589] = 1'b0;  wr_cycle[18589] = 1'b0;  addr_rom[18589]='h00000000;  wr_data_rom[18589]='h00000000;
    rd_cycle[18590] = 1'b0;  wr_cycle[18590] = 1'b0;  addr_rom[18590]='h00000000;  wr_data_rom[18590]='h00000000;
    rd_cycle[18591] = 1'b0;  wr_cycle[18591] = 1'b0;  addr_rom[18591]='h00000000;  wr_data_rom[18591]='h00000000;
    rd_cycle[18592] = 1'b0;  wr_cycle[18592] = 1'b0;  addr_rom[18592]='h00000000;  wr_data_rom[18592]='h00000000;
    rd_cycle[18593] = 1'b0;  wr_cycle[18593] = 1'b0;  addr_rom[18593]='h00000000;  wr_data_rom[18593]='h00000000;
    rd_cycle[18594] = 1'b0;  wr_cycle[18594] = 1'b0;  addr_rom[18594]='h00000000;  wr_data_rom[18594]='h00000000;
    rd_cycle[18595] = 1'b0;  wr_cycle[18595] = 1'b0;  addr_rom[18595]='h00000000;  wr_data_rom[18595]='h00000000;
    rd_cycle[18596] = 1'b0;  wr_cycle[18596] = 1'b0;  addr_rom[18596]='h00000000;  wr_data_rom[18596]='h00000000;
    rd_cycle[18597] = 1'b0;  wr_cycle[18597] = 1'b0;  addr_rom[18597]='h00000000;  wr_data_rom[18597]='h00000000;
    rd_cycle[18598] = 1'b0;  wr_cycle[18598] = 1'b0;  addr_rom[18598]='h00000000;  wr_data_rom[18598]='h00000000;
    rd_cycle[18599] = 1'b0;  wr_cycle[18599] = 1'b0;  addr_rom[18599]='h00000000;  wr_data_rom[18599]='h00000000;
    rd_cycle[18600] = 1'b0;  wr_cycle[18600] = 1'b0;  addr_rom[18600]='h00000000;  wr_data_rom[18600]='h00000000;
    rd_cycle[18601] = 1'b0;  wr_cycle[18601] = 1'b0;  addr_rom[18601]='h00000000;  wr_data_rom[18601]='h00000000;
    rd_cycle[18602] = 1'b0;  wr_cycle[18602] = 1'b0;  addr_rom[18602]='h00000000;  wr_data_rom[18602]='h00000000;
    rd_cycle[18603] = 1'b0;  wr_cycle[18603] = 1'b0;  addr_rom[18603]='h00000000;  wr_data_rom[18603]='h00000000;
    rd_cycle[18604] = 1'b0;  wr_cycle[18604] = 1'b0;  addr_rom[18604]='h00000000;  wr_data_rom[18604]='h00000000;
    rd_cycle[18605] = 1'b0;  wr_cycle[18605] = 1'b0;  addr_rom[18605]='h00000000;  wr_data_rom[18605]='h00000000;
    rd_cycle[18606] = 1'b0;  wr_cycle[18606] = 1'b0;  addr_rom[18606]='h00000000;  wr_data_rom[18606]='h00000000;
    rd_cycle[18607] = 1'b0;  wr_cycle[18607] = 1'b0;  addr_rom[18607]='h00000000;  wr_data_rom[18607]='h00000000;
    rd_cycle[18608] = 1'b0;  wr_cycle[18608] = 1'b0;  addr_rom[18608]='h00000000;  wr_data_rom[18608]='h00000000;
    rd_cycle[18609] = 1'b0;  wr_cycle[18609] = 1'b0;  addr_rom[18609]='h00000000;  wr_data_rom[18609]='h00000000;
    rd_cycle[18610] = 1'b0;  wr_cycle[18610] = 1'b0;  addr_rom[18610]='h00000000;  wr_data_rom[18610]='h00000000;
    rd_cycle[18611] = 1'b0;  wr_cycle[18611] = 1'b0;  addr_rom[18611]='h00000000;  wr_data_rom[18611]='h00000000;
    rd_cycle[18612] = 1'b0;  wr_cycle[18612] = 1'b0;  addr_rom[18612]='h00000000;  wr_data_rom[18612]='h00000000;
    rd_cycle[18613] = 1'b0;  wr_cycle[18613] = 1'b0;  addr_rom[18613]='h00000000;  wr_data_rom[18613]='h00000000;
    rd_cycle[18614] = 1'b0;  wr_cycle[18614] = 1'b0;  addr_rom[18614]='h00000000;  wr_data_rom[18614]='h00000000;
    rd_cycle[18615] = 1'b0;  wr_cycle[18615] = 1'b0;  addr_rom[18615]='h00000000;  wr_data_rom[18615]='h00000000;
    rd_cycle[18616] = 1'b0;  wr_cycle[18616] = 1'b0;  addr_rom[18616]='h00000000;  wr_data_rom[18616]='h00000000;
    rd_cycle[18617] = 1'b0;  wr_cycle[18617] = 1'b0;  addr_rom[18617]='h00000000;  wr_data_rom[18617]='h00000000;
    rd_cycle[18618] = 1'b0;  wr_cycle[18618] = 1'b0;  addr_rom[18618]='h00000000;  wr_data_rom[18618]='h00000000;
    rd_cycle[18619] = 1'b0;  wr_cycle[18619] = 1'b0;  addr_rom[18619]='h00000000;  wr_data_rom[18619]='h00000000;
    rd_cycle[18620] = 1'b0;  wr_cycle[18620] = 1'b0;  addr_rom[18620]='h00000000;  wr_data_rom[18620]='h00000000;
    rd_cycle[18621] = 1'b0;  wr_cycle[18621] = 1'b0;  addr_rom[18621]='h00000000;  wr_data_rom[18621]='h00000000;
    rd_cycle[18622] = 1'b0;  wr_cycle[18622] = 1'b0;  addr_rom[18622]='h00000000;  wr_data_rom[18622]='h00000000;
    rd_cycle[18623] = 1'b0;  wr_cycle[18623] = 1'b0;  addr_rom[18623]='h00000000;  wr_data_rom[18623]='h00000000;
    rd_cycle[18624] = 1'b0;  wr_cycle[18624] = 1'b0;  addr_rom[18624]='h00000000;  wr_data_rom[18624]='h00000000;
    rd_cycle[18625] = 1'b0;  wr_cycle[18625] = 1'b0;  addr_rom[18625]='h00000000;  wr_data_rom[18625]='h00000000;
    rd_cycle[18626] = 1'b0;  wr_cycle[18626] = 1'b0;  addr_rom[18626]='h00000000;  wr_data_rom[18626]='h00000000;
    rd_cycle[18627] = 1'b0;  wr_cycle[18627] = 1'b0;  addr_rom[18627]='h00000000;  wr_data_rom[18627]='h00000000;
    rd_cycle[18628] = 1'b0;  wr_cycle[18628] = 1'b0;  addr_rom[18628]='h00000000;  wr_data_rom[18628]='h00000000;
    rd_cycle[18629] = 1'b0;  wr_cycle[18629] = 1'b0;  addr_rom[18629]='h00000000;  wr_data_rom[18629]='h00000000;
    rd_cycle[18630] = 1'b0;  wr_cycle[18630] = 1'b0;  addr_rom[18630]='h00000000;  wr_data_rom[18630]='h00000000;
    rd_cycle[18631] = 1'b0;  wr_cycle[18631] = 1'b0;  addr_rom[18631]='h00000000;  wr_data_rom[18631]='h00000000;
    rd_cycle[18632] = 1'b0;  wr_cycle[18632] = 1'b0;  addr_rom[18632]='h00000000;  wr_data_rom[18632]='h00000000;
    rd_cycle[18633] = 1'b0;  wr_cycle[18633] = 1'b0;  addr_rom[18633]='h00000000;  wr_data_rom[18633]='h00000000;
    rd_cycle[18634] = 1'b0;  wr_cycle[18634] = 1'b0;  addr_rom[18634]='h00000000;  wr_data_rom[18634]='h00000000;
    rd_cycle[18635] = 1'b0;  wr_cycle[18635] = 1'b0;  addr_rom[18635]='h00000000;  wr_data_rom[18635]='h00000000;
    rd_cycle[18636] = 1'b0;  wr_cycle[18636] = 1'b0;  addr_rom[18636]='h00000000;  wr_data_rom[18636]='h00000000;
    rd_cycle[18637] = 1'b0;  wr_cycle[18637] = 1'b0;  addr_rom[18637]='h00000000;  wr_data_rom[18637]='h00000000;
    rd_cycle[18638] = 1'b0;  wr_cycle[18638] = 1'b0;  addr_rom[18638]='h00000000;  wr_data_rom[18638]='h00000000;
    rd_cycle[18639] = 1'b0;  wr_cycle[18639] = 1'b0;  addr_rom[18639]='h00000000;  wr_data_rom[18639]='h00000000;
    rd_cycle[18640] = 1'b0;  wr_cycle[18640] = 1'b0;  addr_rom[18640]='h00000000;  wr_data_rom[18640]='h00000000;
    rd_cycle[18641] = 1'b0;  wr_cycle[18641] = 1'b0;  addr_rom[18641]='h00000000;  wr_data_rom[18641]='h00000000;
    rd_cycle[18642] = 1'b0;  wr_cycle[18642] = 1'b0;  addr_rom[18642]='h00000000;  wr_data_rom[18642]='h00000000;
    rd_cycle[18643] = 1'b0;  wr_cycle[18643] = 1'b0;  addr_rom[18643]='h00000000;  wr_data_rom[18643]='h00000000;
    rd_cycle[18644] = 1'b0;  wr_cycle[18644] = 1'b0;  addr_rom[18644]='h00000000;  wr_data_rom[18644]='h00000000;
    rd_cycle[18645] = 1'b0;  wr_cycle[18645] = 1'b0;  addr_rom[18645]='h00000000;  wr_data_rom[18645]='h00000000;
    rd_cycle[18646] = 1'b0;  wr_cycle[18646] = 1'b0;  addr_rom[18646]='h00000000;  wr_data_rom[18646]='h00000000;
    rd_cycle[18647] = 1'b0;  wr_cycle[18647] = 1'b0;  addr_rom[18647]='h00000000;  wr_data_rom[18647]='h00000000;
    rd_cycle[18648] = 1'b0;  wr_cycle[18648] = 1'b0;  addr_rom[18648]='h00000000;  wr_data_rom[18648]='h00000000;
    rd_cycle[18649] = 1'b0;  wr_cycle[18649] = 1'b0;  addr_rom[18649]='h00000000;  wr_data_rom[18649]='h00000000;
    rd_cycle[18650] = 1'b0;  wr_cycle[18650] = 1'b0;  addr_rom[18650]='h00000000;  wr_data_rom[18650]='h00000000;
    rd_cycle[18651] = 1'b0;  wr_cycle[18651] = 1'b0;  addr_rom[18651]='h00000000;  wr_data_rom[18651]='h00000000;
    rd_cycle[18652] = 1'b0;  wr_cycle[18652] = 1'b0;  addr_rom[18652]='h00000000;  wr_data_rom[18652]='h00000000;
    rd_cycle[18653] = 1'b0;  wr_cycle[18653] = 1'b0;  addr_rom[18653]='h00000000;  wr_data_rom[18653]='h00000000;
    rd_cycle[18654] = 1'b0;  wr_cycle[18654] = 1'b0;  addr_rom[18654]='h00000000;  wr_data_rom[18654]='h00000000;
    rd_cycle[18655] = 1'b0;  wr_cycle[18655] = 1'b0;  addr_rom[18655]='h00000000;  wr_data_rom[18655]='h00000000;
    rd_cycle[18656] = 1'b0;  wr_cycle[18656] = 1'b0;  addr_rom[18656]='h00000000;  wr_data_rom[18656]='h00000000;
    rd_cycle[18657] = 1'b0;  wr_cycle[18657] = 1'b0;  addr_rom[18657]='h00000000;  wr_data_rom[18657]='h00000000;
    rd_cycle[18658] = 1'b0;  wr_cycle[18658] = 1'b0;  addr_rom[18658]='h00000000;  wr_data_rom[18658]='h00000000;
    rd_cycle[18659] = 1'b0;  wr_cycle[18659] = 1'b0;  addr_rom[18659]='h00000000;  wr_data_rom[18659]='h00000000;
    rd_cycle[18660] = 1'b0;  wr_cycle[18660] = 1'b0;  addr_rom[18660]='h00000000;  wr_data_rom[18660]='h00000000;
    rd_cycle[18661] = 1'b0;  wr_cycle[18661] = 1'b0;  addr_rom[18661]='h00000000;  wr_data_rom[18661]='h00000000;
    rd_cycle[18662] = 1'b0;  wr_cycle[18662] = 1'b0;  addr_rom[18662]='h00000000;  wr_data_rom[18662]='h00000000;
    rd_cycle[18663] = 1'b0;  wr_cycle[18663] = 1'b0;  addr_rom[18663]='h00000000;  wr_data_rom[18663]='h00000000;
    rd_cycle[18664] = 1'b0;  wr_cycle[18664] = 1'b0;  addr_rom[18664]='h00000000;  wr_data_rom[18664]='h00000000;
    rd_cycle[18665] = 1'b0;  wr_cycle[18665] = 1'b0;  addr_rom[18665]='h00000000;  wr_data_rom[18665]='h00000000;
    rd_cycle[18666] = 1'b0;  wr_cycle[18666] = 1'b0;  addr_rom[18666]='h00000000;  wr_data_rom[18666]='h00000000;
    rd_cycle[18667] = 1'b0;  wr_cycle[18667] = 1'b0;  addr_rom[18667]='h00000000;  wr_data_rom[18667]='h00000000;
    rd_cycle[18668] = 1'b0;  wr_cycle[18668] = 1'b0;  addr_rom[18668]='h00000000;  wr_data_rom[18668]='h00000000;
    rd_cycle[18669] = 1'b0;  wr_cycle[18669] = 1'b0;  addr_rom[18669]='h00000000;  wr_data_rom[18669]='h00000000;
    rd_cycle[18670] = 1'b0;  wr_cycle[18670] = 1'b0;  addr_rom[18670]='h00000000;  wr_data_rom[18670]='h00000000;
    rd_cycle[18671] = 1'b0;  wr_cycle[18671] = 1'b0;  addr_rom[18671]='h00000000;  wr_data_rom[18671]='h00000000;
    rd_cycle[18672] = 1'b0;  wr_cycle[18672] = 1'b0;  addr_rom[18672]='h00000000;  wr_data_rom[18672]='h00000000;
    rd_cycle[18673] = 1'b0;  wr_cycle[18673] = 1'b0;  addr_rom[18673]='h00000000;  wr_data_rom[18673]='h00000000;
    rd_cycle[18674] = 1'b0;  wr_cycle[18674] = 1'b0;  addr_rom[18674]='h00000000;  wr_data_rom[18674]='h00000000;
    rd_cycle[18675] = 1'b0;  wr_cycle[18675] = 1'b0;  addr_rom[18675]='h00000000;  wr_data_rom[18675]='h00000000;
    rd_cycle[18676] = 1'b0;  wr_cycle[18676] = 1'b0;  addr_rom[18676]='h00000000;  wr_data_rom[18676]='h00000000;
    rd_cycle[18677] = 1'b0;  wr_cycle[18677] = 1'b0;  addr_rom[18677]='h00000000;  wr_data_rom[18677]='h00000000;
    rd_cycle[18678] = 1'b0;  wr_cycle[18678] = 1'b0;  addr_rom[18678]='h00000000;  wr_data_rom[18678]='h00000000;
    rd_cycle[18679] = 1'b0;  wr_cycle[18679] = 1'b0;  addr_rom[18679]='h00000000;  wr_data_rom[18679]='h00000000;
    rd_cycle[18680] = 1'b0;  wr_cycle[18680] = 1'b0;  addr_rom[18680]='h00000000;  wr_data_rom[18680]='h00000000;
    rd_cycle[18681] = 1'b0;  wr_cycle[18681] = 1'b0;  addr_rom[18681]='h00000000;  wr_data_rom[18681]='h00000000;
    rd_cycle[18682] = 1'b0;  wr_cycle[18682] = 1'b0;  addr_rom[18682]='h00000000;  wr_data_rom[18682]='h00000000;
    rd_cycle[18683] = 1'b0;  wr_cycle[18683] = 1'b0;  addr_rom[18683]='h00000000;  wr_data_rom[18683]='h00000000;
    rd_cycle[18684] = 1'b0;  wr_cycle[18684] = 1'b0;  addr_rom[18684]='h00000000;  wr_data_rom[18684]='h00000000;
    rd_cycle[18685] = 1'b0;  wr_cycle[18685] = 1'b0;  addr_rom[18685]='h00000000;  wr_data_rom[18685]='h00000000;
    rd_cycle[18686] = 1'b0;  wr_cycle[18686] = 1'b0;  addr_rom[18686]='h00000000;  wr_data_rom[18686]='h00000000;
    rd_cycle[18687] = 1'b0;  wr_cycle[18687] = 1'b0;  addr_rom[18687]='h00000000;  wr_data_rom[18687]='h00000000;
    rd_cycle[18688] = 1'b0;  wr_cycle[18688] = 1'b0;  addr_rom[18688]='h00000000;  wr_data_rom[18688]='h00000000;
    rd_cycle[18689] = 1'b0;  wr_cycle[18689] = 1'b0;  addr_rom[18689]='h00000000;  wr_data_rom[18689]='h00000000;
    rd_cycle[18690] = 1'b0;  wr_cycle[18690] = 1'b0;  addr_rom[18690]='h00000000;  wr_data_rom[18690]='h00000000;
    rd_cycle[18691] = 1'b0;  wr_cycle[18691] = 1'b0;  addr_rom[18691]='h00000000;  wr_data_rom[18691]='h00000000;
    rd_cycle[18692] = 1'b0;  wr_cycle[18692] = 1'b0;  addr_rom[18692]='h00000000;  wr_data_rom[18692]='h00000000;
    rd_cycle[18693] = 1'b0;  wr_cycle[18693] = 1'b0;  addr_rom[18693]='h00000000;  wr_data_rom[18693]='h00000000;
    rd_cycle[18694] = 1'b0;  wr_cycle[18694] = 1'b0;  addr_rom[18694]='h00000000;  wr_data_rom[18694]='h00000000;
    rd_cycle[18695] = 1'b0;  wr_cycle[18695] = 1'b0;  addr_rom[18695]='h00000000;  wr_data_rom[18695]='h00000000;
    rd_cycle[18696] = 1'b0;  wr_cycle[18696] = 1'b0;  addr_rom[18696]='h00000000;  wr_data_rom[18696]='h00000000;
    rd_cycle[18697] = 1'b0;  wr_cycle[18697] = 1'b0;  addr_rom[18697]='h00000000;  wr_data_rom[18697]='h00000000;
    rd_cycle[18698] = 1'b0;  wr_cycle[18698] = 1'b0;  addr_rom[18698]='h00000000;  wr_data_rom[18698]='h00000000;
    rd_cycle[18699] = 1'b0;  wr_cycle[18699] = 1'b0;  addr_rom[18699]='h00000000;  wr_data_rom[18699]='h00000000;
    rd_cycle[18700] = 1'b0;  wr_cycle[18700] = 1'b0;  addr_rom[18700]='h00000000;  wr_data_rom[18700]='h00000000;
    rd_cycle[18701] = 1'b0;  wr_cycle[18701] = 1'b0;  addr_rom[18701]='h00000000;  wr_data_rom[18701]='h00000000;
    rd_cycle[18702] = 1'b0;  wr_cycle[18702] = 1'b0;  addr_rom[18702]='h00000000;  wr_data_rom[18702]='h00000000;
    rd_cycle[18703] = 1'b0;  wr_cycle[18703] = 1'b0;  addr_rom[18703]='h00000000;  wr_data_rom[18703]='h00000000;
    rd_cycle[18704] = 1'b0;  wr_cycle[18704] = 1'b0;  addr_rom[18704]='h00000000;  wr_data_rom[18704]='h00000000;
    rd_cycle[18705] = 1'b0;  wr_cycle[18705] = 1'b0;  addr_rom[18705]='h00000000;  wr_data_rom[18705]='h00000000;
    rd_cycle[18706] = 1'b0;  wr_cycle[18706] = 1'b0;  addr_rom[18706]='h00000000;  wr_data_rom[18706]='h00000000;
    rd_cycle[18707] = 1'b0;  wr_cycle[18707] = 1'b0;  addr_rom[18707]='h00000000;  wr_data_rom[18707]='h00000000;
    rd_cycle[18708] = 1'b0;  wr_cycle[18708] = 1'b0;  addr_rom[18708]='h00000000;  wr_data_rom[18708]='h00000000;
    rd_cycle[18709] = 1'b0;  wr_cycle[18709] = 1'b0;  addr_rom[18709]='h00000000;  wr_data_rom[18709]='h00000000;
    rd_cycle[18710] = 1'b0;  wr_cycle[18710] = 1'b0;  addr_rom[18710]='h00000000;  wr_data_rom[18710]='h00000000;
    rd_cycle[18711] = 1'b0;  wr_cycle[18711] = 1'b0;  addr_rom[18711]='h00000000;  wr_data_rom[18711]='h00000000;
    rd_cycle[18712] = 1'b0;  wr_cycle[18712] = 1'b0;  addr_rom[18712]='h00000000;  wr_data_rom[18712]='h00000000;
    rd_cycle[18713] = 1'b0;  wr_cycle[18713] = 1'b0;  addr_rom[18713]='h00000000;  wr_data_rom[18713]='h00000000;
    rd_cycle[18714] = 1'b0;  wr_cycle[18714] = 1'b0;  addr_rom[18714]='h00000000;  wr_data_rom[18714]='h00000000;
    rd_cycle[18715] = 1'b0;  wr_cycle[18715] = 1'b0;  addr_rom[18715]='h00000000;  wr_data_rom[18715]='h00000000;
    rd_cycle[18716] = 1'b0;  wr_cycle[18716] = 1'b0;  addr_rom[18716]='h00000000;  wr_data_rom[18716]='h00000000;
    rd_cycle[18717] = 1'b0;  wr_cycle[18717] = 1'b0;  addr_rom[18717]='h00000000;  wr_data_rom[18717]='h00000000;
    rd_cycle[18718] = 1'b0;  wr_cycle[18718] = 1'b0;  addr_rom[18718]='h00000000;  wr_data_rom[18718]='h00000000;
    rd_cycle[18719] = 1'b0;  wr_cycle[18719] = 1'b0;  addr_rom[18719]='h00000000;  wr_data_rom[18719]='h00000000;
    rd_cycle[18720] = 1'b0;  wr_cycle[18720] = 1'b0;  addr_rom[18720]='h00000000;  wr_data_rom[18720]='h00000000;
    rd_cycle[18721] = 1'b0;  wr_cycle[18721] = 1'b0;  addr_rom[18721]='h00000000;  wr_data_rom[18721]='h00000000;
    rd_cycle[18722] = 1'b0;  wr_cycle[18722] = 1'b0;  addr_rom[18722]='h00000000;  wr_data_rom[18722]='h00000000;
    rd_cycle[18723] = 1'b0;  wr_cycle[18723] = 1'b0;  addr_rom[18723]='h00000000;  wr_data_rom[18723]='h00000000;
    rd_cycle[18724] = 1'b0;  wr_cycle[18724] = 1'b0;  addr_rom[18724]='h00000000;  wr_data_rom[18724]='h00000000;
    rd_cycle[18725] = 1'b0;  wr_cycle[18725] = 1'b0;  addr_rom[18725]='h00000000;  wr_data_rom[18725]='h00000000;
    rd_cycle[18726] = 1'b0;  wr_cycle[18726] = 1'b0;  addr_rom[18726]='h00000000;  wr_data_rom[18726]='h00000000;
    rd_cycle[18727] = 1'b0;  wr_cycle[18727] = 1'b0;  addr_rom[18727]='h00000000;  wr_data_rom[18727]='h00000000;
    rd_cycle[18728] = 1'b0;  wr_cycle[18728] = 1'b0;  addr_rom[18728]='h00000000;  wr_data_rom[18728]='h00000000;
    rd_cycle[18729] = 1'b0;  wr_cycle[18729] = 1'b0;  addr_rom[18729]='h00000000;  wr_data_rom[18729]='h00000000;
    rd_cycle[18730] = 1'b0;  wr_cycle[18730] = 1'b0;  addr_rom[18730]='h00000000;  wr_data_rom[18730]='h00000000;
    rd_cycle[18731] = 1'b0;  wr_cycle[18731] = 1'b0;  addr_rom[18731]='h00000000;  wr_data_rom[18731]='h00000000;
    rd_cycle[18732] = 1'b0;  wr_cycle[18732] = 1'b0;  addr_rom[18732]='h00000000;  wr_data_rom[18732]='h00000000;
    rd_cycle[18733] = 1'b0;  wr_cycle[18733] = 1'b0;  addr_rom[18733]='h00000000;  wr_data_rom[18733]='h00000000;
    rd_cycle[18734] = 1'b0;  wr_cycle[18734] = 1'b0;  addr_rom[18734]='h00000000;  wr_data_rom[18734]='h00000000;
    rd_cycle[18735] = 1'b0;  wr_cycle[18735] = 1'b0;  addr_rom[18735]='h00000000;  wr_data_rom[18735]='h00000000;
    rd_cycle[18736] = 1'b0;  wr_cycle[18736] = 1'b0;  addr_rom[18736]='h00000000;  wr_data_rom[18736]='h00000000;
    rd_cycle[18737] = 1'b0;  wr_cycle[18737] = 1'b0;  addr_rom[18737]='h00000000;  wr_data_rom[18737]='h00000000;
    rd_cycle[18738] = 1'b0;  wr_cycle[18738] = 1'b0;  addr_rom[18738]='h00000000;  wr_data_rom[18738]='h00000000;
    rd_cycle[18739] = 1'b0;  wr_cycle[18739] = 1'b0;  addr_rom[18739]='h00000000;  wr_data_rom[18739]='h00000000;
    rd_cycle[18740] = 1'b0;  wr_cycle[18740] = 1'b0;  addr_rom[18740]='h00000000;  wr_data_rom[18740]='h00000000;
    rd_cycle[18741] = 1'b0;  wr_cycle[18741] = 1'b0;  addr_rom[18741]='h00000000;  wr_data_rom[18741]='h00000000;
    rd_cycle[18742] = 1'b0;  wr_cycle[18742] = 1'b0;  addr_rom[18742]='h00000000;  wr_data_rom[18742]='h00000000;
    rd_cycle[18743] = 1'b0;  wr_cycle[18743] = 1'b0;  addr_rom[18743]='h00000000;  wr_data_rom[18743]='h00000000;
    rd_cycle[18744] = 1'b0;  wr_cycle[18744] = 1'b0;  addr_rom[18744]='h00000000;  wr_data_rom[18744]='h00000000;
    rd_cycle[18745] = 1'b0;  wr_cycle[18745] = 1'b0;  addr_rom[18745]='h00000000;  wr_data_rom[18745]='h00000000;
    rd_cycle[18746] = 1'b0;  wr_cycle[18746] = 1'b0;  addr_rom[18746]='h00000000;  wr_data_rom[18746]='h00000000;
    rd_cycle[18747] = 1'b0;  wr_cycle[18747] = 1'b0;  addr_rom[18747]='h00000000;  wr_data_rom[18747]='h00000000;
    rd_cycle[18748] = 1'b0;  wr_cycle[18748] = 1'b0;  addr_rom[18748]='h00000000;  wr_data_rom[18748]='h00000000;
    rd_cycle[18749] = 1'b0;  wr_cycle[18749] = 1'b0;  addr_rom[18749]='h00000000;  wr_data_rom[18749]='h00000000;
    rd_cycle[18750] = 1'b0;  wr_cycle[18750] = 1'b0;  addr_rom[18750]='h00000000;  wr_data_rom[18750]='h00000000;
    rd_cycle[18751] = 1'b0;  wr_cycle[18751] = 1'b0;  addr_rom[18751]='h00000000;  wr_data_rom[18751]='h00000000;
    rd_cycle[18752] = 1'b0;  wr_cycle[18752] = 1'b0;  addr_rom[18752]='h00000000;  wr_data_rom[18752]='h00000000;
    rd_cycle[18753] = 1'b0;  wr_cycle[18753] = 1'b0;  addr_rom[18753]='h00000000;  wr_data_rom[18753]='h00000000;
    rd_cycle[18754] = 1'b0;  wr_cycle[18754] = 1'b0;  addr_rom[18754]='h00000000;  wr_data_rom[18754]='h00000000;
    rd_cycle[18755] = 1'b0;  wr_cycle[18755] = 1'b0;  addr_rom[18755]='h00000000;  wr_data_rom[18755]='h00000000;
    rd_cycle[18756] = 1'b0;  wr_cycle[18756] = 1'b0;  addr_rom[18756]='h00000000;  wr_data_rom[18756]='h00000000;
    rd_cycle[18757] = 1'b0;  wr_cycle[18757] = 1'b0;  addr_rom[18757]='h00000000;  wr_data_rom[18757]='h00000000;
    rd_cycle[18758] = 1'b0;  wr_cycle[18758] = 1'b0;  addr_rom[18758]='h00000000;  wr_data_rom[18758]='h00000000;
    rd_cycle[18759] = 1'b0;  wr_cycle[18759] = 1'b0;  addr_rom[18759]='h00000000;  wr_data_rom[18759]='h00000000;
    rd_cycle[18760] = 1'b0;  wr_cycle[18760] = 1'b0;  addr_rom[18760]='h00000000;  wr_data_rom[18760]='h00000000;
    rd_cycle[18761] = 1'b0;  wr_cycle[18761] = 1'b0;  addr_rom[18761]='h00000000;  wr_data_rom[18761]='h00000000;
    rd_cycle[18762] = 1'b0;  wr_cycle[18762] = 1'b0;  addr_rom[18762]='h00000000;  wr_data_rom[18762]='h00000000;
    rd_cycle[18763] = 1'b0;  wr_cycle[18763] = 1'b0;  addr_rom[18763]='h00000000;  wr_data_rom[18763]='h00000000;
    rd_cycle[18764] = 1'b0;  wr_cycle[18764] = 1'b0;  addr_rom[18764]='h00000000;  wr_data_rom[18764]='h00000000;
    rd_cycle[18765] = 1'b0;  wr_cycle[18765] = 1'b0;  addr_rom[18765]='h00000000;  wr_data_rom[18765]='h00000000;
    rd_cycle[18766] = 1'b0;  wr_cycle[18766] = 1'b0;  addr_rom[18766]='h00000000;  wr_data_rom[18766]='h00000000;
    rd_cycle[18767] = 1'b0;  wr_cycle[18767] = 1'b0;  addr_rom[18767]='h00000000;  wr_data_rom[18767]='h00000000;
    rd_cycle[18768] = 1'b0;  wr_cycle[18768] = 1'b0;  addr_rom[18768]='h00000000;  wr_data_rom[18768]='h00000000;
    rd_cycle[18769] = 1'b0;  wr_cycle[18769] = 1'b0;  addr_rom[18769]='h00000000;  wr_data_rom[18769]='h00000000;
    rd_cycle[18770] = 1'b0;  wr_cycle[18770] = 1'b0;  addr_rom[18770]='h00000000;  wr_data_rom[18770]='h00000000;
    rd_cycle[18771] = 1'b0;  wr_cycle[18771] = 1'b0;  addr_rom[18771]='h00000000;  wr_data_rom[18771]='h00000000;
    rd_cycle[18772] = 1'b0;  wr_cycle[18772] = 1'b0;  addr_rom[18772]='h00000000;  wr_data_rom[18772]='h00000000;
    rd_cycle[18773] = 1'b0;  wr_cycle[18773] = 1'b0;  addr_rom[18773]='h00000000;  wr_data_rom[18773]='h00000000;
    rd_cycle[18774] = 1'b0;  wr_cycle[18774] = 1'b0;  addr_rom[18774]='h00000000;  wr_data_rom[18774]='h00000000;
    rd_cycle[18775] = 1'b0;  wr_cycle[18775] = 1'b0;  addr_rom[18775]='h00000000;  wr_data_rom[18775]='h00000000;
    rd_cycle[18776] = 1'b0;  wr_cycle[18776] = 1'b0;  addr_rom[18776]='h00000000;  wr_data_rom[18776]='h00000000;
    rd_cycle[18777] = 1'b0;  wr_cycle[18777] = 1'b0;  addr_rom[18777]='h00000000;  wr_data_rom[18777]='h00000000;
    rd_cycle[18778] = 1'b0;  wr_cycle[18778] = 1'b0;  addr_rom[18778]='h00000000;  wr_data_rom[18778]='h00000000;
    rd_cycle[18779] = 1'b0;  wr_cycle[18779] = 1'b0;  addr_rom[18779]='h00000000;  wr_data_rom[18779]='h00000000;
    rd_cycle[18780] = 1'b0;  wr_cycle[18780] = 1'b0;  addr_rom[18780]='h00000000;  wr_data_rom[18780]='h00000000;
    rd_cycle[18781] = 1'b0;  wr_cycle[18781] = 1'b0;  addr_rom[18781]='h00000000;  wr_data_rom[18781]='h00000000;
    rd_cycle[18782] = 1'b0;  wr_cycle[18782] = 1'b0;  addr_rom[18782]='h00000000;  wr_data_rom[18782]='h00000000;
    rd_cycle[18783] = 1'b0;  wr_cycle[18783] = 1'b0;  addr_rom[18783]='h00000000;  wr_data_rom[18783]='h00000000;
    rd_cycle[18784] = 1'b0;  wr_cycle[18784] = 1'b0;  addr_rom[18784]='h00000000;  wr_data_rom[18784]='h00000000;
    rd_cycle[18785] = 1'b0;  wr_cycle[18785] = 1'b0;  addr_rom[18785]='h00000000;  wr_data_rom[18785]='h00000000;
    rd_cycle[18786] = 1'b0;  wr_cycle[18786] = 1'b0;  addr_rom[18786]='h00000000;  wr_data_rom[18786]='h00000000;
    rd_cycle[18787] = 1'b0;  wr_cycle[18787] = 1'b0;  addr_rom[18787]='h00000000;  wr_data_rom[18787]='h00000000;
    rd_cycle[18788] = 1'b0;  wr_cycle[18788] = 1'b0;  addr_rom[18788]='h00000000;  wr_data_rom[18788]='h00000000;
    rd_cycle[18789] = 1'b0;  wr_cycle[18789] = 1'b0;  addr_rom[18789]='h00000000;  wr_data_rom[18789]='h00000000;
    rd_cycle[18790] = 1'b0;  wr_cycle[18790] = 1'b0;  addr_rom[18790]='h00000000;  wr_data_rom[18790]='h00000000;
    rd_cycle[18791] = 1'b0;  wr_cycle[18791] = 1'b0;  addr_rom[18791]='h00000000;  wr_data_rom[18791]='h00000000;
    rd_cycle[18792] = 1'b0;  wr_cycle[18792] = 1'b0;  addr_rom[18792]='h00000000;  wr_data_rom[18792]='h00000000;
    rd_cycle[18793] = 1'b0;  wr_cycle[18793] = 1'b0;  addr_rom[18793]='h00000000;  wr_data_rom[18793]='h00000000;
    rd_cycle[18794] = 1'b0;  wr_cycle[18794] = 1'b0;  addr_rom[18794]='h00000000;  wr_data_rom[18794]='h00000000;
    rd_cycle[18795] = 1'b0;  wr_cycle[18795] = 1'b0;  addr_rom[18795]='h00000000;  wr_data_rom[18795]='h00000000;
    rd_cycle[18796] = 1'b0;  wr_cycle[18796] = 1'b0;  addr_rom[18796]='h00000000;  wr_data_rom[18796]='h00000000;
    rd_cycle[18797] = 1'b0;  wr_cycle[18797] = 1'b0;  addr_rom[18797]='h00000000;  wr_data_rom[18797]='h00000000;
    rd_cycle[18798] = 1'b0;  wr_cycle[18798] = 1'b0;  addr_rom[18798]='h00000000;  wr_data_rom[18798]='h00000000;
    rd_cycle[18799] = 1'b0;  wr_cycle[18799] = 1'b0;  addr_rom[18799]='h00000000;  wr_data_rom[18799]='h00000000;
    rd_cycle[18800] = 1'b0;  wr_cycle[18800] = 1'b0;  addr_rom[18800]='h00000000;  wr_data_rom[18800]='h00000000;
    rd_cycle[18801] = 1'b0;  wr_cycle[18801] = 1'b0;  addr_rom[18801]='h00000000;  wr_data_rom[18801]='h00000000;
    rd_cycle[18802] = 1'b0;  wr_cycle[18802] = 1'b0;  addr_rom[18802]='h00000000;  wr_data_rom[18802]='h00000000;
    rd_cycle[18803] = 1'b0;  wr_cycle[18803] = 1'b0;  addr_rom[18803]='h00000000;  wr_data_rom[18803]='h00000000;
    rd_cycle[18804] = 1'b0;  wr_cycle[18804] = 1'b0;  addr_rom[18804]='h00000000;  wr_data_rom[18804]='h00000000;
    rd_cycle[18805] = 1'b0;  wr_cycle[18805] = 1'b0;  addr_rom[18805]='h00000000;  wr_data_rom[18805]='h00000000;
    rd_cycle[18806] = 1'b0;  wr_cycle[18806] = 1'b0;  addr_rom[18806]='h00000000;  wr_data_rom[18806]='h00000000;
    rd_cycle[18807] = 1'b0;  wr_cycle[18807] = 1'b0;  addr_rom[18807]='h00000000;  wr_data_rom[18807]='h00000000;
    rd_cycle[18808] = 1'b0;  wr_cycle[18808] = 1'b0;  addr_rom[18808]='h00000000;  wr_data_rom[18808]='h00000000;
    rd_cycle[18809] = 1'b0;  wr_cycle[18809] = 1'b0;  addr_rom[18809]='h00000000;  wr_data_rom[18809]='h00000000;
    rd_cycle[18810] = 1'b0;  wr_cycle[18810] = 1'b0;  addr_rom[18810]='h00000000;  wr_data_rom[18810]='h00000000;
    rd_cycle[18811] = 1'b0;  wr_cycle[18811] = 1'b0;  addr_rom[18811]='h00000000;  wr_data_rom[18811]='h00000000;
    rd_cycle[18812] = 1'b0;  wr_cycle[18812] = 1'b0;  addr_rom[18812]='h00000000;  wr_data_rom[18812]='h00000000;
    rd_cycle[18813] = 1'b0;  wr_cycle[18813] = 1'b0;  addr_rom[18813]='h00000000;  wr_data_rom[18813]='h00000000;
    rd_cycle[18814] = 1'b0;  wr_cycle[18814] = 1'b0;  addr_rom[18814]='h00000000;  wr_data_rom[18814]='h00000000;
    rd_cycle[18815] = 1'b0;  wr_cycle[18815] = 1'b0;  addr_rom[18815]='h00000000;  wr_data_rom[18815]='h00000000;
    rd_cycle[18816] = 1'b0;  wr_cycle[18816] = 1'b0;  addr_rom[18816]='h00000000;  wr_data_rom[18816]='h00000000;
    rd_cycle[18817] = 1'b0;  wr_cycle[18817] = 1'b0;  addr_rom[18817]='h00000000;  wr_data_rom[18817]='h00000000;
    rd_cycle[18818] = 1'b0;  wr_cycle[18818] = 1'b0;  addr_rom[18818]='h00000000;  wr_data_rom[18818]='h00000000;
    rd_cycle[18819] = 1'b0;  wr_cycle[18819] = 1'b0;  addr_rom[18819]='h00000000;  wr_data_rom[18819]='h00000000;
    rd_cycle[18820] = 1'b0;  wr_cycle[18820] = 1'b0;  addr_rom[18820]='h00000000;  wr_data_rom[18820]='h00000000;
    rd_cycle[18821] = 1'b0;  wr_cycle[18821] = 1'b0;  addr_rom[18821]='h00000000;  wr_data_rom[18821]='h00000000;
    rd_cycle[18822] = 1'b0;  wr_cycle[18822] = 1'b0;  addr_rom[18822]='h00000000;  wr_data_rom[18822]='h00000000;
    rd_cycle[18823] = 1'b0;  wr_cycle[18823] = 1'b0;  addr_rom[18823]='h00000000;  wr_data_rom[18823]='h00000000;
    rd_cycle[18824] = 1'b0;  wr_cycle[18824] = 1'b0;  addr_rom[18824]='h00000000;  wr_data_rom[18824]='h00000000;
    rd_cycle[18825] = 1'b0;  wr_cycle[18825] = 1'b0;  addr_rom[18825]='h00000000;  wr_data_rom[18825]='h00000000;
    rd_cycle[18826] = 1'b0;  wr_cycle[18826] = 1'b0;  addr_rom[18826]='h00000000;  wr_data_rom[18826]='h00000000;
    rd_cycle[18827] = 1'b0;  wr_cycle[18827] = 1'b0;  addr_rom[18827]='h00000000;  wr_data_rom[18827]='h00000000;
    rd_cycle[18828] = 1'b0;  wr_cycle[18828] = 1'b0;  addr_rom[18828]='h00000000;  wr_data_rom[18828]='h00000000;
    rd_cycle[18829] = 1'b0;  wr_cycle[18829] = 1'b0;  addr_rom[18829]='h00000000;  wr_data_rom[18829]='h00000000;
    rd_cycle[18830] = 1'b0;  wr_cycle[18830] = 1'b0;  addr_rom[18830]='h00000000;  wr_data_rom[18830]='h00000000;
    rd_cycle[18831] = 1'b0;  wr_cycle[18831] = 1'b0;  addr_rom[18831]='h00000000;  wr_data_rom[18831]='h00000000;
    rd_cycle[18832] = 1'b0;  wr_cycle[18832] = 1'b0;  addr_rom[18832]='h00000000;  wr_data_rom[18832]='h00000000;
    rd_cycle[18833] = 1'b0;  wr_cycle[18833] = 1'b0;  addr_rom[18833]='h00000000;  wr_data_rom[18833]='h00000000;
    rd_cycle[18834] = 1'b0;  wr_cycle[18834] = 1'b0;  addr_rom[18834]='h00000000;  wr_data_rom[18834]='h00000000;
    rd_cycle[18835] = 1'b0;  wr_cycle[18835] = 1'b0;  addr_rom[18835]='h00000000;  wr_data_rom[18835]='h00000000;
    rd_cycle[18836] = 1'b0;  wr_cycle[18836] = 1'b0;  addr_rom[18836]='h00000000;  wr_data_rom[18836]='h00000000;
    rd_cycle[18837] = 1'b0;  wr_cycle[18837] = 1'b0;  addr_rom[18837]='h00000000;  wr_data_rom[18837]='h00000000;
    rd_cycle[18838] = 1'b0;  wr_cycle[18838] = 1'b0;  addr_rom[18838]='h00000000;  wr_data_rom[18838]='h00000000;
    rd_cycle[18839] = 1'b0;  wr_cycle[18839] = 1'b0;  addr_rom[18839]='h00000000;  wr_data_rom[18839]='h00000000;
    rd_cycle[18840] = 1'b0;  wr_cycle[18840] = 1'b0;  addr_rom[18840]='h00000000;  wr_data_rom[18840]='h00000000;
    rd_cycle[18841] = 1'b0;  wr_cycle[18841] = 1'b0;  addr_rom[18841]='h00000000;  wr_data_rom[18841]='h00000000;
    rd_cycle[18842] = 1'b0;  wr_cycle[18842] = 1'b0;  addr_rom[18842]='h00000000;  wr_data_rom[18842]='h00000000;
    rd_cycle[18843] = 1'b0;  wr_cycle[18843] = 1'b0;  addr_rom[18843]='h00000000;  wr_data_rom[18843]='h00000000;
    rd_cycle[18844] = 1'b0;  wr_cycle[18844] = 1'b0;  addr_rom[18844]='h00000000;  wr_data_rom[18844]='h00000000;
    rd_cycle[18845] = 1'b0;  wr_cycle[18845] = 1'b0;  addr_rom[18845]='h00000000;  wr_data_rom[18845]='h00000000;
    rd_cycle[18846] = 1'b0;  wr_cycle[18846] = 1'b0;  addr_rom[18846]='h00000000;  wr_data_rom[18846]='h00000000;
    rd_cycle[18847] = 1'b0;  wr_cycle[18847] = 1'b0;  addr_rom[18847]='h00000000;  wr_data_rom[18847]='h00000000;
    rd_cycle[18848] = 1'b0;  wr_cycle[18848] = 1'b0;  addr_rom[18848]='h00000000;  wr_data_rom[18848]='h00000000;
    rd_cycle[18849] = 1'b0;  wr_cycle[18849] = 1'b0;  addr_rom[18849]='h00000000;  wr_data_rom[18849]='h00000000;
    rd_cycle[18850] = 1'b0;  wr_cycle[18850] = 1'b0;  addr_rom[18850]='h00000000;  wr_data_rom[18850]='h00000000;
    rd_cycle[18851] = 1'b0;  wr_cycle[18851] = 1'b0;  addr_rom[18851]='h00000000;  wr_data_rom[18851]='h00000000;
    rd_cycle[18852] = 1'b0;  wr_cycle[18852] = 1'b0;  addr_rom[18852]='h00000000;  wr_data_rom[18852]='h00000000;
    rd_cycle[18853] = 1'b0;  wr_cycle[18853] = 1'b0;  addr_rom[18853]='h00000000;  wr_data_rom[18853]='h00000000;
    rd_cycle[18854] = 1'b0;  wr_cycle[18854] = 1'b0;  addr_rom[18854]='h00000000;  wr_data_rom[18854]='h00000000;
    rd_cycle[18855] = 1'b0;  wr_cycle[18855] = 1'b0;  addr_rom[18855]='h00000000;  wr_data_rom[18855]='h00000000;
    rd_cycle[18856] = 1'b0;  wr_cycle[18856] = 1'b0;  addr_rom[18856]='h00000000;  wr_data_rom[18856]='h00000000;
    rd_cycle[18857] = 1'b0;  wr_cycle[18857] = 1'b0;  addr_rom[18857]='h00000000;  wr_data_rom[18857]='h00000000;
    rd_cycle[18858] = 1'b0;  wr_cycle[18858] = 1'b0;  addr_rom[18858]='h00000000;  wr_data_rom[18858]='h00000000;
    rd_cycle[18859] = 1'b0;  wr_cycle[18859] = 1'b0;  addr_rom[18859]='h00000000;  wr_data_rom[18859]='h00000000;
    rd_cycle[18860] = 1'b0;  wr_cycle[18860] = 1'b0;  addr_rom[18860]='h00000000;  wr_data_rom[18860]='h00000000;
    rd_cycle[18861] = 1'b0;  wr_cycle[18861] = 1'b0;  addr_rom[18861]='h00000000;  wr_data_rom[18861]='h00000000;
    rd_cycle[18862] = 1'b0;  wr_cycle[18862] = 1'b0;  addr_rom[18862]='h00000000;  wr_data_rom[18862]='h00000000;
    rd_cycle[18863] = 1'b0;  wr_cycle[18863] = 1'b0;  addr_rom[18863]='h00000000;  wr_data_rom[18863]='h00000000;
    rd_cycle[18864] = 1'b0;  wr_cycle[18864] = 1'b0;  addr_rom[18864]='h00000000;  wr_data_rom[18864]='h00000000;
    rd_cycle[18865] = 1'b0;  wr_cycle[18865] = 1'b0;  addr_rom[18865]='h00000000;  wr_data_rom[18865]='h00000000;
    rd_cycle[18866] = 1'b0;  wr_cycle[18866] = 1'b0;  addr_rom[18866]='h00000000;  wr_data_rom[18866]='h00000000;
    rd_cycle[18867] = 1'b0;  wr_cycle[18867] = 1'b0;  addr_rom[18867]='h00000000;  wr_data_rom[18867]='h00000000;
    rd_cycle[18868] = 1'b0;  wr_cycle[18868] = 1'b0;  addr_rom[18868]='h00000000;  wr_data_rom[18868]='h00000000;
    rd_cycle[18869] = 1'b0;  wr_cycle[18869] = 1'b0;  addr_rom[18869]='h00000000;  wr_data_rom[18869]='h00000000;
    rd_cycle[18870] = 1'b0;  wr_cycle[18870] = 1'b0;  addr_rom[18870]='h00000000;  wr_data_rom[18870]='h00000000;
    rd_cycle[18871] = 1'b0;  wr_cycle[18871] = 1'b0;  addr_rom[18871]='h00000000;  wr_data_rom[18871]='h00000000;
    rd_cycle[18872] = 1'b0;  wr_cycle[18872] = 1'b0;  addr_rom[18872]='h00000000;  wr_data_rom[18872]='h00000000;
    rd_cycle[18873] = 1'b0;  wr_cycle[18873] = 1'b0;  addr_rom[18873]='h00000000;  wr_data_rom[18873]='h00000000;
    rd_cycle[18874] = 1'b0;  wr_cycle[18874] = 1'b0;  addr_rom[18874]='h00000000;  wr_data_rom[18874]='h00000000;
    rd_cycle[18875] = 1'b0;  wr_cycle[18875] = 1'b0;  addr_rom[18875]='h00000000;  wr_data_rom[18875]='h00000000;
    rd_cycle[18876] = 1'b0;  wr_cycle[18876] = 1'b0;  addr_rom[18876]='h00000000;  wr_data_rom[18876]='h00000000;
    rd_cycle[18877] = 1'b0;  wr_cycle[18877] = 1'b0;  addr_rom[18877]='h00000000;  wr_data_rom[18877]='h00000000;
    rd_cycle[18878] = 1'b0;  wr_cycle[18878] = 1'b0;  addr_rom[18878]='h00000000;  wr_data_rom[18878]='h00000000;
    rd_cycle[18879] = 1'b0;  wr_cycle[18879] = 1'b0;  addr_rom[18879]='h00000000;  wr_data_rom[18879]='h00000000;
    rd_cycle[18880] = 1'b0;  wr_cycle[18880] = 1'b0;  addr_rom[18880]='h00000000;  wr_data_rom[18880]='h00000000;
    rd_cycle[18881] = 1'b0;  wr_cycle[18881] = 1'b0;  addr_rom[18881]='h00000000;  wr_data_rom[18881]='h00000000;
    rd_cycle[18882] = 1'b0;  wr_cycle[18882] = 1'b0;  addr_rom[18882]='h00000000;  wr_data_rom[18882]='h00000000;
    rd_cycle[18883] = 1'b0;  wr_cycle[18883] = 1'b0;  addr_rom[18883]='h00000000;  wr_data_rom[18883]='h00000000;
    rd_cycle[18884] = 1'b0;  wr_cycle[18884] = 1'b0;  addr_rom[18884]='h00000000;  wr_data_rom[18884]='h00000000;
    rd_cycle[18885] = 1'b0;  wr_cycle[18885] = 1'b0;  addr_rom[18885]='h00000000;  wr_data_rom[18885]='h00000000;
    rd_cycle[18886] = 1'b0;  wr_cycle[18886] = 1'b0;  addr_rom[18886]='h00000000;  wr_data_rom[18886]='h00000000;
    rd_cycle[18887] = 1'b0;  wr_cycle[18887] = 1'b0;  addr_rom[18887]='h00000000;  wr_data_rom[18887]='h00000000;
    rd_cycle[18888] = 1'b0;  wr_cycle[18888] = 1'b0;  addr_rom[18888]='h00000000;  wr_data_rom[18888]='h00000000;
    rd_cycle[18889] = 1'b0;  wr_cycle[18889] = 1'b0;  addr_rom[18889]='h00000000;  wr_data_rom[18889]='h00000000;
    rd_cycle[18890] = 1'b0;  wr_cycle[18890] = 1'b0;  addr_rom[18890]='h00000000;  wr_data_rom[18890]='h00000000;
    rd_cycle[18891] = 1'b0;  wr_cycle[18891] = 1'b0;  addr_rom[18891]='h00000000;  wr_data_rom[18891]='h00000000;
    rd_cycle[18892] = 1'b0;  wr_cycle[18892] = 1'b0;  addr_rom[18892]='h00000000;  wr_data_rom[18892]='h00000000;
    rd_cycle[18893] = 1'b0;  wr_cycle[18893] = 1'b0;  addr_rom[18893]='h00000000;  wr_data_rom[18893]='h00000000;
    rd_cycle[18894] = 1'b0;  wr_cycle[18894] = 1'b0;  addr_rom[18894]='h00000000;  wr_data_rom[18894]='h00000000;
    rd_cycle[18895] = 1'b0;  wr_cycle[18895] = 1'b0;  addr_rom[18895]='h00000000;  wr_data_rom[18895]='h00000000;
    rd_cycle[18896] = 1'b0;  wr_cycle[18896] = 1'b0;  addr_rom[18896]='h00000000;  wr_data_rom[18896]='h00000000;
    rd_cycle[18897] = 1'b0;  wr_cycle[18897] = 1'b0;  addr_rom[18897]='h00000000;  wr_data_rom[18897]='h00000000;
    rd_cycle[18898] = 1'b0;  wr_cycle[18898] = 1'b0;  addr_rom[18898]='h00000000;  wr_data_rom[18898]='h00000000;
    rd_cycle[18899] = 1'b0;  wr_cycle[18899] = 1'b0;  addr_rom[18899]='h00000000;  wr_data_rom[18899]='h00000000;
    rd_cycle[18900] = 1'b0;  wr_cycle[18900] = 1'b0;  addr_rom[18900]='h00000000;  wr_data_rom[18900]='h00000000;
    rd_cycle[18901] = 1'b0;  wr_cycle[18901] = 1'b0;  addr_rom[18901]='h00000000;  wr_data_rom[18901]='h00000000;
    rd_cycle[18902] = 1'b0;  wr_cycle[18902] = 1'b0;  addr_rom[18902]='h00000000;  wr_data_rom[18902]='h00000000;
    rd_cycle[18903] = 1'b0;  wr_cycle[18903] = 1'b0;  addr_rom[18903]='h00000000;  wr_data_rom[18903]='h00000000;
    rd_cycle[18904] = 1'b0;  wr_cycle[18904] = 1'b0;  addr_rom[18904]='h00000000;  wr_data_rom[18904]='h00000000;
    rd_cycle[18905] = 1'b0;  wr_cycle[18905] = 1'b0;  addr_rom[18905]='h00000000;  wr_data_rom[18905]='h00000000;
    rd_cycle[18906] = 1'b0;  wr_cycle[18906] = 1'b0;  addr_rom[18906]='h00000000;  wr_data_rom[18906]='h00000000;
    rd_cycle[18907] = 1'b0;  wr_cycle[18907] = 1'b0;  addr_rom[18907]='h00000000;  wr_data_rom[18907]='h00000000;
    rd_cycle[18908] = 1'b0;  wr_cycle[18908] = 1'b0;  addr_rom[18908]='h00000000;  wr_data_rom[18908]='h00000000;
    rd_cycle[18909] = 1'b0;  wr_cycle[18909] = 1'b0;  addr_rom[18909]='h00000000;  wr_data_rom[18909]='h00000000;
    rd_cycle[18910] = 1'b0;  wr_cycle[18910] = 1'b0;  addr_rom[18910]='h00000000;  wr_data_rom[18910]='h00000000;
    rd_cycle[18911] = 1'b0;  wr_cycle[18911] = 1'b0;  addr_rom[18911]='h00000000;  wr_data_rom[18911]='h00000000;
    rd_cycle[18912] = 1'b0;  wr_cycle[18912] = 1'b0;  addr_rom[18912]='h00000000;  wr_data_rom[18912]='h00000000;
    rd_cycle[18913] = 1'b0;  wr_cycle[18913] = 1'b0;  addr_rom[18913]='h00000000;  wr_data_rom[18913]='h00000000;
    rd_cycle[18914] = 1'b0;  wr_cycle[18914] = 1'b0;  addr_rom[18914]='h00000000;  wr_data_rom[18914]='h00000000;
    rd_cycle[18915] = 1'b0;  wr_cycle[18915] = 1'b0;  addr_rom[18915]='h00000000;  wr_data_rom[18915]='h00000000;
    rd_cycle[18916] = 1'b0;  wr_cycle[18916] = 1'b0;  addr_rom[18916]='h00000000;  wr_data_rom[18916]='h00000000;
    rd_cycle[18917] = 1'b0;  wr_cycle[18917] = 1'b0;  addr_rom[18917]='h00000000;  wr_data_rom[18917]='h00000000;
    rd_cycle[18918] = 1'b0;  wr_cycle[18918] = 1'b0;  addr_rom[18918]='h00000000;  wr_data_rom[18918]='h00000000;
    rd_cycle[18919] = 1'b0;  wr_cycle[18919] = 1'b0;  addr_rom[18919]='h00000000;  wr_data_rom[18919]='h00000000;
    rd_cycle[18920] = 1'b0;  wr_cycle[18920] = 1'b0;  addr_rom[18920]='h00000000;  wr_data_rom[18920]='h00000000;
    rd_cycle[18921] = 1'b0;  wr_cycle[18921] = 1'b0;  addr_rom[18921]='h00000000;  wr_data_rom[18921]='h00000000;
    rd_cycle[18922] = 1'b0;  wr_cycle[18922] = 1'b0;  addr_rom[18922]='h00000000;  wr_data_rom[18922]='h00000000;
    rd_cycle[18923] = 1'b0;  wr_cycle[18923] = 1'b0;  addr_rom[18923]='h00000000;  wr_data_rom[18923]='h00000000;
    rd_cycle[18924] = 1'b0;  wr_cycle[18924] = 1'b0;  addr_rom[18924]='h00000000;  wr_data_rom[18924]='h00000000;
    rd_cycle[18925] = 1'b0;  wr_cycle[18925] = 1'b0;  addr_rom[18925]='h00000000;  wr_data_rom[18925]='h00000000;
    rd_cycle[18926] = 1'b0;  wr_cycle[18926] = 1'b0;  addr_rom[18926]='h00000000;  wr_data_rom[18926]='h00000000;
    rd_cycle[18927] = 1'b0;  wr_cycle[18927] = 1'b0;  addr_rom[18927]='h00000000;  wr_data_rom[18927]='h00000000;
    rd_cycle[18928] = 1'b0;  wr_cycle[18928] = 1'b0;  addr_rom[18928]='h00000000;  wr_data_rom[18928]='h00000000;
    rd_cycle[18929] = 1'b0;  wr_cycle[18929] = 1'b0;  addr_rom[18929]='h00000000;  wr_data_rom[18929]='h00000000;
    rd_cycle[18930] = 1'b0;  wr_cycle[18930] = 1'b0;  addr_rom[18930]='h00000000;  wr_data_rom[18930]='h00000000;
    rd_cycle[18931] = 1'b0;  wr_cycle[18931] = 1'b0;  addr_rom[18931]='h00000000;  wr_data_rom[18931]='h00000000;
    rd_cycle[18932] = 1'b0;  wr_cycle[18932] = 1'b0;  addr_rom[18932]='h00000000;  wr_data_rom[18932]='h00000000;
    rd_cycle[18933] = 1'b0;  wr_cycle[18933] = 1'b0;  addr_rom[18933]='h00000000;  wr_data_rom[18933]='h00000000;
    rd_cycle[18934] = 1'b0;  wr_cycle[18934] = 1'b0;  addr_rom[18934]='h00000000;  wr_data_rom[18934]='h00000000;
    rd_cycle[18935] = 1'b0;  wr_cycle[18935] = 1'b0;  addr_rom[18935]='h00000000;  wr_data_rom[18935]='h00000000;
    rd_cycle[18936] = 1'b0;  wr_cycle[18936] = 1'b0;  addr_rom[18936]='h00000000;  wr_data_rom[18936]='h00000000;
    rd_cycle[18937] = 1'b0;  wr_cycle[18937] = 1'b0;  addr_rom[18937]='h00000000;  wr_data_rom[18937]='h00000000;
    rd_cycle[18938] = 1'b0;  wr_cycle[18938] = 1'b0;  addr_rom[18938]='h00000000;  wr_data_rom[18938]='h00000000;
    rd_cycle[18939] = 1'b0;  wr_cycle[18939] = 1'b0;  addr_rom[18939]='h00000000;  wr_data_rom[18939]='h00000000;
    rd_cycle[18940] = 1'b0;  wr_cycle[18940] = 1'b0;  addr_rom[18940]='h00000000;  wr_data_rom[18940]='h00000000;
    rd_cycle[18941] = 1'b0;  wr_cycle[18941] = 1'b0;  addr_rom[18941]='h00000000;  wr_data_rom[18941]='h00000000;
    rd_cycle[18942] = 1'b0;  wr_cycle[18942] = 1'b0;  addr_rom[18942]='h00000000;  wr_data_rom[18942]='h00000000;
    rd_cycle[18943] = 1'b0;  wr_cycle[18943] = 1'b0;  addr_rom[18943]='h00000000;  wr_data_rom[18943]='h00000000;
    rd_cycle[18944] = 1'b0;  wr_cycle[18944] = 1'b0;  addr_rom[18944]='h00000000;  wr_data_rom[18944]='h00000000;
    rd_cycle[18945] = 1'b0;  wr_cycle[18945] = 1'b0;  addr_rom[18945]='h00000000;  wr_data_rom[18945]='h00000000;
    rd_cycle[18946] = 1'b0;  wr_cycle[18946] = 1'b0;  addr_rom[18946]='h00000000;  wr_data_rom[18946]='h00000000;
    rd_cycle[18947] = 1'b0;  wr_cycle[18947] = 1'b0;  addr_rom[18947]='h00000000;  wr_data_rom[18947]='h00000000;
    rd_cycle[18948] = 1'b0;  wr_cycle[18948] = 1'b0;  addr_rom[18948]='h00000000;  wr_data_rom[18948]='h00000000;
    rd_cycle[18949] = 1'b0;  wr_cycle[18949] = 1'b0;  addr_rom[18949]='h00000000;  wr_data_rom[18949]='h00000000;
    rd_cycle[18950] = 1'b0;  wr_cycle[18950] = 1'b0;  addr_rom[18950]='h00000000;  wr_data_rom[18950]='h00000000;
    rd_cycle[18951] = 1'b0;  wr_cycle[18951] = 1'b0;  addr_rom[18951]='h00000000;  wr_data_rom[18951]='h00000000;
    rd_cycle[18952] = 1'b0;  wr_cycle[18952] = 1'b0;  addr_rom[18952]='h00000000;  wr_data_rom[18952]='h00000000;
    rd_cycle[18953] = 1'b0;  wr_cycle[18953] = 1'b0;  addr_rom[18953]='h00000000;  wr_data_rom[18953]='h00000000;
    rd_cycle[18954] = 1'b0;  wr_cycle[18954] = 1'b0;  addr_rom[18954]='h00000000;  wr_data_rom[18954]='h00000000;
    rd_cycle[18955] = 1'b0;  wr_cycle[18955] = 1'b0;  addr_rom[18955]='h00000000;  wr_data_rom[18955]='h00000000;
    rd_cycle[18956] = 1'b0;  wr_cycle[18956] = 1'b0;  addr_rom[18956]='h00000000;  wr_data_rom[18956]='h00000000;
    rd_cycle[18957] = 1'b0;  wr_cycle[18957] = 1'b0;  addr_rom[18957]='h00000000;  wr_data_rom[18957]='h00000000;
    rd_cycle[18958] = 1'b0;  wr_cycle[18958] = 1'b0;  addr_rom[18958]='h00000000;  wr_data_rom[18958]='h00000000;
    rd_cycle[18959] = 1'b0;  wr_cycle[18959] = 1'b0;  addr_rom[18959]='h00000000;  wr_data_rom[18959]='h00000000;
    rd_cycle[18960] = 1'b0;  wr_cycle[18960] = 1'b0;  addr_rom[18960]='h00000000;  wr_data_rom[18960]='h00000000;
    rd_cycle[18961] = 1'b0;  wr_cycle[18961] = 1'b0;  addr_rom[18961]='h00000000;  wr_data_rom[18961]='h00000000;
    rd_cycle[18962] = 1'b0;  wr_cycle[18962] = 1'b0;  addr_rom[18962]='h00000000;  wr_data_rom[18962]='h00000000;
    rd_cycle[18963] = 1'b0;  wr_cycle[18963] = 1'b0;  addr_rom[18963]='h00000000;  wr_data_rom[18963]='h00000000;
    rd_cycle[18964] = 1'b0;  wr_cycle[18964] = 1'b0;  addr_rom[18964]='h00000000;  wr_data_rom[18964]='h00000000;
    rd_cycle[18965] = 1'b0;  wr_cycle[18965] = 1'b0;  addr_rom[18965]='h00000000;  wr_data_rom[18965]='h00000000;
    rd_cycle[18966] = 1'b0;  wr_cycle[18966] = 1'b0;  addr_rom[18966]='h00000000;  wr_data_rom[18966]='h00000000;
    rd_cycle[18967] = 1'b0;  wr_cycle[18967] = 1'b0;  addr_rom[18967]='h00000000;  wr_data_rom[18967]='h00000000;
    rd_cycle[18968] = 1'b0;  wr_cycle[18968] = 1'b0;  addr_rom[18968]='h00000000;  wr_data_rom[18968]='h00000000;
    rd_cycle[18969] = 1'b0;  wr_cycle[18969] = 1'b0;  addr_rom[18969]='h00000000;  wr_data_rom[18969]='h00000000;
    rd_cycle[18970] = 1'b0;  wr_cycle[18970] = 1'b0;  addr_rom[18970]='h00000000;  wr_data_rom[18970]='h00000000;
    rd_cycle[18971] = 1'b0;  wr_cycle[18971] = 1'b0;  addr_rom[18971]='h00000000;  wr_data_rom[18971]='h00000000;
    rd_cycle[18972] = 1'b0;  wr_cycle[18972] = 1'b0;  addr_rom[18972]='h00000000;  wr_data_rom[18972]='h00000000;
    rd_cycle[18973] = 1'b0;  wr_cycle[18973] = 1'b0;  addr_rom[18973]='h00000000;  wr_data_rom[18973]='h00000000;
    rd_cycle[18974] = 1'b0;  wr_cycle[18974] = 1'b0;  addr_rom[18974]='h00000000;  wr_data_rom[18974]='h00000000;
    rd_cycle[18975] = 1'b0;  wr_cycle[18975] = 1'b0;  addr_rom[18975]='h00000000;  wr_data_rom[18975]='h00000000;
    rd_cycle[18976] = 1'b0;  wr_cycle[18976] = 1'b0;  addr_rom[18976]='h00000000;  wr_data_rom[18976]='h00000000;
    rd_cycle[18977] = 1'b0;  wr_cycle[18977] = 1'b0;  addr_rom[18977]='h00000000;  wr_data_rom[18977]='h00000000;
    rd_cycle[18978] = 1'b0;  wr_cycle[18978] = 1'b0;  addr_rom[18978]='h00000000;  wr_data_rom[18978]='h00000000;
    rd_cycle[18979] = 1'b0;  wr_cycle[18979] = 1'b0;  addr_rom[18979]='h00000000;  wr_data_rom[18979]='h00000000;
    rd_cycle[18980] = 1'b0;  wr_cycle[18980] = 1'b0;  addr_rom[18980]='h00000000;  wr_data_rom[18980]='h00000000;
    rd_cycle[18981] = 1'b0;  wr_cycle[18981] = 1'b0;  addr_rom[18981]='h00000000;  wr_data_rom[18981]='h00000000;
    rd_cycle[18982] = 1'b0;  wr_cycle[18982] = 1'b0;  addr_rom[18982]='h00000000;  wr_data_rom[18982]='h00000000;
    rd_cycle[18983] = 1'b0;  wr_cycle[18983] = 1'b0;  addr_rom[18983]='h00000000;  wr_data_rom[18983]='h00000000;
    rd_cycle[18984] = 1'b0;  wr_cycle[18984] = 1'b0;  addr_rom[18984]='h00000000;  wr_data_rom[18984]='h00000000;
    rd_cycle[18985] = 1'b0;  wr_cycle[18985] = 1'b0;  addr_rom[18985]='h00000000;  wr_data_rom[18985]='h00000000;
    rd_cycle[18986] = 1'b0;  wr_cycle[18986] = 1'b0;  addr_rom[18986]='h00000000;  wr_data_rom[18986]='h00000000;
    rd_cycle[18987] = 1'b0;  wr_cycle[18987] = 1'b0;  addr_rom[18987]='h00000000;  wr_data_rom[18987]='h00000000;
    rd_cycle[18988] = 1'b0;  wr_cycle[18988] = 1'b0;  addr_rom[18988]='h00000000;  wr_data_rom[18988]='h00000000;
    rd_cycle[18989] = 1'b0;  wr_cycle[18989] = 1'b0;  addr_rom[18989]='h00000000;  wr_data_rom[18989]='h00000000;
    rd_cycle[18990] = 1'b0;  wr_cycle[18990] = 1'b0;  addr_rom[18990]='h00000000;  wr_data_rom[18990]='h00000000;
    rd_cycle[18991] = 1'b0;  wr_cycle[18991] = 1'b0;  addr_rom[18991]='h00000000;  wr_data_rom[18991]='h00000000;
    rd_cycle[18992] = 1'b0;  wr_cycle[18992] = 1'b0;  addr_rom[18992]='h00000000;  wr_data_rom[18992]='h00000000;
    rd_cycle[18993] = 1'b0;  wr_cycle[18993] = 1'b0;  addr_rom[18993]='h00000000;  wr_data_rom[18993]='h00000000;
    rd_cycle[18994] = 1'b0;  wr_cycle[18994] = 1'b0;  addr_rom[18994]='h00000000;  wr_data_rom[18994]='h00000000;
    rd_cycle[18995] = 1'b0;  wr_cycle[18995] = 1'b0;  addr_rom[18995]='h00000000;  wr_data_rom[18995]='h00000000;
    rd_cycle[18996] = 1'b0;  wr_cycle[18996] = 1'b0;  addr_rom[18996]='h00000000;  wr_data_rom[18996]='h00000000;
    rd_cycle[18997] = 1'b0;  wr_cycle[18997] = 1'b0;  addr_rom[18997]='h00000000;  wr_data_rom[18997]='h00000000;
    rd_cycle[18998] = 1'b0;  wr_cycle[18998] = 1'b0;  addr_rom[18998]='h00000000;  wr_data_rom[18998]='h00000000;
    rd_cycle[18999] = 1'b0;  wr_cycle[18999] = 1'b0;  addr_rom[18999]='h00000000;  wr_data_rom[18999]='h00000000;
    rd_cycle[19000] = 1'b0;  wr_cycle[19000] = 1'b0;  addr_rom[19000]='h00000000;  wr_data_rom[19000]='h00000000;
    rd_cycle[19001] = 1'b0;  wr_cycle[19001] = 1'b0;  addr_rom[19001]='h00000000;  wr_data_rom[19001]='h00000000;
    rd_cycle[19002] = 1'b0;  wr_cycle[19002] = 1'b0;  addr_rom[19002]='h00000000;  wr_data_rom[19002]='h00000000;
    rd_cycle[19003] = 1'b0;  wr_cycle[19003] = 1'b0;  addr_rom[19003]='h00000000;  wr_data_rom[19003]='h00000000;
    rd_cycle[19004] = 1'b0;  wr_cycle[19004] = 1'b0;  addr_rom[19004]='h00000000;  wr_data_rom[19004]='h00000000;
    rd_cycle[19005] = 1'b0;  wr_cycle[19005] = 1'b0;  addr_rom[19005]='h00000000;  wr_data_rom[19005]='h00000000;
    rd_cycle[19006] = 1'b0;  wr_cycle[19006] = 1'b0;  addr_rom[19006]='h00000000;  wr_data_rom[19006]='h00000000;
    rd_cycle[19007] = 1'b0;  wr_cycle[19007] = 1'b0;  addr_rom[19007]='h00000000;  wr_data_rom[19007]='h00000000;
    rd_cycle[19008] = 1'b0;  wr_cycle[19008] = 1'b0;  addr_rom[19008]='h00000000;  wr_data_rom[19008]='h00000000;
    rd_cycle[19009] = 1'b0;  wr_cycle[19009] = 1'b0;  addr_rom[19009]='h00000000;  wr_data_rom[19009]='h00000000;
    rd_cycle[19010] = 1'b0;  wr_cycle[19010] = 1'b0;  addr_rom[19010]='h00000000;  wr_data_rom[19010]='h00000000;
    rd_cycle[19011] = 1'b0;  wr_cycle[19011] = 1'b0;  addr_rom[19011]='h00000000;  wr_data_rom[19011]='h00000000;
    rd_cycle[19012] = 1'b0;  wr_cycle[19012] = 1'b0;  addr_rom[19012]='h00000000;  wr_data_rom[19012]='h00000000;
    rd_cycle[19013] = 1'b0;  wr_cycle[19013] = 1'b0;  addr_rom[19013]='h00000000;  wr_data_rom[19013]='h00000000;
    rd_cycle[19014] = 1'b0;  wr_cycle[19014] = 1'b0;  addr_rom[19014]='h00000000;  wr_data_rom[19014]='h00000000;
    rd_cycle[19015] = 1'b0;  wr_cycle[19015] = 1'b0;  addr_rom[19015]='h00000000;  wr_data_rom[19015]='h00000000;
    rd_cycle[19016] = 1'b0;  wr_cycle[19016] = 1'b0;  addr_rom[19016]='h00000000;  wr_data_rom[19016]='h00000000;
    rd_cycle[19017] = 1'b0;  wr_cycle[19017] = 1'b0;  addr_rom[19017]='h00000000;  wr_data_rom[19017]='h00000000;
    rd_cycle[19018] = 1'b0;  wr_cycle[19018] = 1'b0;  addr_rom[19018]='h00000000;  wr_data_rom[19018]='h00000000;
    rd_cycle[19019] = 1'b0;  wr_cycle[19019] = 1'b0;  addr_rom[19019]='h00000000;  wr_data_rom[19019]='h00000000;
    rd_cycle[19020] = 1'b0;  wr_cycle[19020] = 1'b0;  addr_rom[19020]='h00000000;  wr_data_rom[19020]='h00000000;
    rd_cycle[19021] = 1'b0;  wr_cycle[19021] = 1'b0;  addr_rom[19021]='h00000000;  wr_data_rom[19021]='h00000000;
    rd_cycle[19022] = 1'b0;  wr_cycle[19022] = 1'b0;  addr_rom[19022]='h00000000;  wr_data_rom[19022]='h00000000;
    rd_cycle[19023] = 1'b0;  wr_cycle[19023] = 1'b0;  addr_rom[19023]='h00000000;  wr_data_rom[19023]='h00000000;
    rd_cycle[19024] = 1'b0;  wr_cycle[19024] = 1'b0;  addr_rom[19024]='h00000000;  wr_data_rom[19024]='h00000000;
    rd_cycle[19025] = 1'b0;  wr_cycle[19025] = 1'b0;  addr_rom[19025]='h00000000;  wr_data_rom[19025]='h00000000;
    rd_cycle[19026] = 1'b0;  wr_cycle[19026] = 1'b0;  addr_rom[19026]='h00000000;  wr_data_rom[19026]='h00000000;
    rd_cycle[19027] = 1'b0;  wr_cycle[19027] = 1'b0;  addr_rom[19027]='h00000000;  wr_data_rom[19027]='h00000000;
    rd_cycle[19028] = 1'b0;  wr_cycle[19028] = 1'b0;  addr_rom[19028]='h00000000;  wr_data_rom[19028]='h00000000;
    rd_cycle[19029] = 1'b0;  wr_cycle[19029] = 1'b0;  addr_rom[19029]='h00000000;  wr_data_rom[19029]='h00000000;
    rd_cycle[19030] = 1'b0;  wr_cycle[19030] = 1'b0;  addr_rom[19030]='h00000000;  wr_data_rom[19030]='h00000000;
    rd_cycle[19031] = 1'b0;  wr_cycle[19031] = 1'b0;  addr_rom[19031]='h00000000;  wr_data_rom[19031]='h00000000;
    rd_cycle[19032] = 1'b0;  wr_cycle[19032] = 1'b0;  addr_rom[19032]='h00000000;  wr_data_rom[19032]='h00000000;
    rd_cycle[19033] = 1'b0;  wr_cycle[19033] = 1'b0;  addr_rom[19033]='h00000000;  wr_data_rom[19033]='h00000000;
    rd_cycle[19034] = 1'b0;  wr_cycle[19034] = 1'b0;  addr_rom[19034]='h00000000;  wr_data_rom[19034]='h00000000;
    rd_cycle[19035] = 1'b0;  wr_cycle[19035] = 1'b0;  addr_rom[19035]='h00000000;  wr_data_rom[19035]='h00000000;
    rd_cycle[19036] = 1'b0;  wr_cycle[19036] = 1'b0;  addr_rom[19036]='h00000000;  wr_data_rom[19036]='h00000000;
    rd_cycle[19037] = 1'b0;  wr_cycle[19037] = 1'b0;  addr_rom[19037]='h00000000;  wr_data_rom[19037]='h00000000;
    rd_cycle[19038] = 1'b0;  wr_cycle[19038] = 1'b0;  addr_rom[19038]='h00000000;  wr_data_rom[19038]='h00000000;
    rd_cycle[19039] = 1'b0;  wr_cycle[19039] = 1'b0;  addr_rom[19039]='h00000000;  wr_data_rom[19039]='h00000000;
    rd_cycle[19040] = 1'b0;  wr_cycle[19040] = 1'b0;  addr_rom[19040]='h00000000;  wr_data_rom[19040]='h00000000;
    rd_cycle[19041] = 1'b0;  wr_cycle[19041] = 1'b0;  addr_rom[19041]='h00000000;  wr_data_rom[19041]='h00000000;
    rd_cycle[19042] = 1'b0;  wr_cycle[19042] = 1'b0;  addr_rom[19042]='h00000000;  wr_data_rom[19042]='h00000000;
    rd_cycle[19043] = 1'b0;  wr_cycle[19043] = 1'b0;  addr_rom[19043]='h00000000;  wr_data_rom[19043]='h00000000;
    rd_cycle[19044] = 1'b0;  wr_cycle[19044] = 1'b0;  addr_rom[19044]='h00000000;  wr_data_rom[19044]='h00000000;
    rd_cycle[19045] = 1'b0;  wr_cycle[19045] = 1'b0;  addr_rom[19045]='h00000000;  wr_data_rom[19045]='h00000000;
    rd_cycle[19046] = 1'b0;  wr_cycle[19046] = 1'b0;  addr_rom[19046]='h00000000;  wr_data_rom[19046]='h00000000;
    rd_cycle[19047] = 1'b0;  wr_cycle[19047] = 1'b0;  addr_rom[19047]='h00000000;  wr_data_rom[19047]='h00000000;
    rd_cycle[19048] = 1'b0;  wr_cycle[19048] = 1'b0;  addr_rom[19048]='h00000000;  wr_data_rom[19048]='h00000000;
    rd_cycle[19049] = 1'b0;  wr_cycle[19049] = 1'b0;  addr_rom[19049]='h00000000;  wr_data_rom[19049]='h00000000;
    rd_cycle[19050] = 1'b0;  wr_cycle[19050] = 1'b0;  addr_rom[19050]='h00000000;  wr_data_rom[19050]='h00000000;
    rd_cycle[19051] = 1'b0;  wr_cycle[19051] = 1'b0;  addr_rom[19051]='h00000000;  wr_data_rom[19051]='h00000000;
    rd_cycle[19052] = 1'b0;  wr_cycle[19052] = 1'b0;  addr_rom[19052]='h00000000;  wr_data_rom[19052]='h00000000;
    rd_cycle[19053] = 1'b0;  wr_cycle[19053] = 1'b0;  addr_rom[19053]='h00000000;  wr_data_rom[19053]='h00000000;
    rd_cycle[19054] = 1'b0;  wr_cycle[19054] = 1'b0;  addr_rom[19054]='h00000000;  wr_data_rom[19054]='h00000000;
    rd_cycle[19055] = 1'b0;  wr_cycle[19055] = 1'b0;  addr_rom[19055]='h00000000;  wr_data_rom[19055]='h00000000;
    rd_cycle[19056] = 1'b0;  wr_cycle[19056] = 1'b0;  addr_rom[19056]='h00000000;  wr_data_rom[19056]='h00000000;
    rd_cycle[19057] = 1'b0;  wr_cycle[19057] = 1'b0;  addr_rom[19057]='h00000000;  wr_data_rom[19057]='h00000000;
    rd_cycle[19058] = 1'b0;  wr_cycle[19058] = 1'b0;  addr_rom[19058]='h00000000;  wr_data_rom[19058]='h00000000;
    rd_cycle[19059] = 1'b0;  wr_cycle[19059] = 1'b0;  addr_rom[19059]='h00000000;  wr_data_rom[19059]='h00000000;
    rd_cycle[19060] = 1'b0;  wr_cycle[19060] = 1'b0;  addr_rom[19060]='h00000000;  wr_data_rom[19060]='h00000000;
    rd_cycle[19061] = 1'b0;  wr_cycle[19061] = 1'b0;  addr_rom[19061]='h00000000;  wr_data_rom[19061]='h00000000;
    rd_cycle[19062] = 1'b0;  wr_cycle[19062] = 1'b0;  addr_rom[19062]='h00000000;  wr_data_rom[19062]='h00000000;
    rd_cycle[19063] = 1'b0;  wr_cycle[19063] = 1'b0;  addr_rom[19063]='h00000000;  wr_data_rom[19063]='h00000000;
    rd_cycle[19064] = 1'b0;  wr_cycle[19064] = 1'b0;  addr_rom[19064]='h00000000;  wr_data_rom[19064]='h00000000;
    rd_cycle[19065] = 1'b0;  wr_cycle[19065] = 1'b0;  addr_rom[19065]='h00000000;  wr_data_rom[19065]='h00000000;
    rd_cycle[19066] = 1'b0;  wr_cycle[19066] = 1'b0;  addr_rom[19066]='h00000000;  wr_data_rom[19066]='h00000000;
    rd_cycle[19067] = 1'b0;  wr_cycle[19067] = 1'b0;  addr_rom[19067]='h00000000;  wr_data_rom[19067]='h00000000;
    rd_cycle[19068] = 1'b0;  wr_cycle[19068] = 1'b0;  addr_rom[19068]='h00000000;  wr_data_rom[19068]='h00000000;
    rd_cycle[19069] = 1'b0;  wr_cycle[19069] = 1'b0;  addr_rom[19069]='h00000000;  wr_data_rom[19069]='h00000000;
    rd_cycle[19070] = 1'b0;  wr_cycle[19070] = 1'b0;  addr_rom[19070]='h00000000;  wr_data_rom[19070]='h00000000;
    rd_cycle[19071] = 1'b0;  wr_cycle[19071] = 1'b0;  addr_rom[19071]='h00000000;  wr_data_rom[19071]='h00000000;
    rd_cycle[19072] = 1'b0;  wr_cycle[19072] = 1'b0;  addr_rom[19072]='h00000000;  wr_data_rom[19072]='h00000000;
    rd_cycle[19073] = 1'b0;  wr_cycle[19073] = 1'b0;  addr_rom[19073]='h00000000;  wr_data_rom[19073]='h00000000;
    rd_cycle[19074] = 1'b0;  wr_cycle[19074] = 1'b0;  addr_rom[19074]='h00000000;  wr_data_rom[19074]='h00000000;
    rd_cycle[19075] = 1'b0;  wr_cycle[19075] = 1'b0;  addr_rom[19075]='h00000000;  wr_data_rom[19075]='h00000000;
    rd_cycle[19076] = 1'b0;  wr_cycle[19076] = 1'b0;  addr_rom[19076]='h00000000;  wr_data_rom[19076]='h00000000;
    rd_cycle[19077] = 1'b0;  wr_cycle[19077] = 1'b0;  addr_rom[19077]='h00000000;  wr_data_rom[19077]='h00000000;
    rd_cycle[19078] = 1'b0;  wr_cycle[19078] = 1'b0;  addr_rom[19078]='h00000000;  wr_data_rom[19078]='h00000000;
    rd_cycle[19079] = 1'b0;  wr_cycle[19079] = 1'b0;  addr_rom[19079]='h00000000;  wr_data_rom[19079]='h00000000;
    rd_cycle[19080] = 1'b0;  wr_cycle[19080] = 1'b0;  addr_rom[19080]='h00000000;  wr_data_rom[19080]='h00000000;
    rd_cycle[19081] = 1'b0;  wr_cycle[19081] = 1'b0;  addr_rom[19081]='h00000000;  wr_data_rom[19081]='h00000000;
    rd_cycle[19082] = 1'b0;  wr_cycle[19082] = 1'b0;  addr_rom[19082]='h00000000;  wr_data_rom[19082]='h00000000;
    rd_cycle[19083] = 1'b0;  wr_cycle[19083] = 1'b0;  addr_rom[19083]='h00000000;  wr_data_rom[19083]='h00000000;
    rd_cycle[19084] = 1'b0;  wr_cycle[19084] = 1'b0;  addr_rom[19084]='h00000000;  wr_data_rom[19084]='h00000000;
    rd_cycle[19085] = 1'b0;  wr_cycle[19085] = 1'b0;  addr_rom[19085]='h00000000;  wr_data_rom[19085]='h00000000;
    rd_cycle[19086] = 1'b0;  wr_cycle[19086] = 1'b0;  addr_rom[19086]='h00000000;  wr_data_rom[19086]='h00000000;
    rd_cycle[19087] = 1'b0;  wr_cycle[19087] = 1'b0;  addr_rom[19087]='h00000000;  wr_data_rom[19087]='h00000000;
    rd_cycle[19088] = 1'b0;  wr_cycle[19088] = 1'b0;  addr_rom[19088]='h00000000;  wr_data_rom[19088]='h00000000;
    rd_cycle[19089] = 1'b0;  wr_cycle[19089] = 1'b0;  addr_rom[19089]='h00000000;  wr_data_rom[19089]='h00000000;
    rd_cycle[19090] = 1'b0;  wr_cycle[19090] = 1'b0;  addr_rom[19090]='h00000000;  wr_data_rom[19090]='h00000000;
    rd_cycle[19091] = 1'b0;  wr_cycle[19091] = 1'b0;  addr_rom[19091]='h00000000;  wr_data_rom[19091]='h00000000;
    rd_cycle[19092] = 1'b0;  wr_cycle[19092] = 1'b0;  addr_rom[19092]='h00000000;  wr_data_rom[19092]='h00000000;
    rd_cycle[19093] = 1'b0;  wr_cycle[19093] = 1'b0;  addr_rom[19093]='h00000000;  wr_data_rom[19093]='h00000000;
    rd_cycle[19094] = 1'b0;  wr_cycle[19094] = 1'b0;  addr_rom[19094]='h00000000;  wr_data_rom[19094]='h00000000;
    rd_cycle[19095] = 1'b0;  wr_cycle[19095] = 1'b0;  addr_rom[19095]='h00000000;  wr_data_rom[19095]='h00000000;
    rd_cycle[19096] = 1'b0;  wr_cycle[19096] = 1'b0;  addr_rom[19096]='h00000000;  wr_data_rom[19096]='h00000000;
    rd_cycle[19097] = 1'b0;  wr_cycle[19097] = 1'b0;  addr_rom[19097]='h00000000;  wr_data_rom[19097]='h00000000;
    rd_cycle[19098] = 1'b0;  wr_cycle[19098] = 1'b0;  addr_rom[19098]='h00000000;  wr_data_rom[19098]='h00000000;
    rd_cycle[19099] = 1'b0;  wr_cycle[19099] = 1'b0;  addr_rom[19099]='h00000000;  wr_data_rom[19099]='h00000000;
    rd_cycle[19100] = 1'b0;  wr_cycle[19100] = 1'b0;  addr_rom[19100]='h00000000;  wr_data_rom[19100]='h00000000;
    rd_cycle[19101] = 1'b0;  wr_cycle[19101] = 1'b0;  addr_rom[19101]='h00000000;  wr_data_rom[19101]='h00000000;
    rd_cycle[19102] = 1'b0;  wr_cycle[19102] = 1'b0;  addr_rom[19102]='h00000000;  wr_data_rom[19102]='h00000000;
    rd_cycle[19103] = 1'b0;  wr_cycle[19103] = 1'b0;  addr_rom[19103]='h00000000;  wr_data_rom[19103]='h00000000;
    rd_cycle[19104] = 1'b0;  wr_cycle[19104] = 1'b0;  addr_rom[19104]='h00000000;  wr_data_rom[19104]='h00000000;
    rd_cycle[19105] = 1'b0;  wr_cycle[19105] = 1'b0;  addr_rom[19105]='h00000000;  wr_data_rom[19105]='h00000000;
    rd_cycle[19106] = 1'b0;  wr_cycle[19106] = 1'b0;  addr_rom[19106]='h00000000;  wr_data_rom[19106]='h00000000;
    rd_cycle[19107] = 1'b0;  wr_cycle[19107] = 1'b0;  addr_rom[19107]='h00000000;  wr_data_rom[19107]='h00000000;
    rd_cycle[19108] = 1'b0;  wr_cycle[19108] = 1'b0;  addr_rom[19108]='h00000000;  wr_data_rom[19108]='h00000000;
    rd_cycle[19109] = 1'b0;  wr_cycle[19109] = 1'b0;  addr_rom[19109]='h00000000;  wr_data_rom[19109]='h00000000;
    rd_cycle[19110] = 1'b0;  wr_cycle[19110] = 1'b0;  addr_rom[19110]='h00000000;  wr_data_rom[19110]='h00000000;
    rd_cycle[19111] = 1'b0;  wr_cycle[19111] = 1'b0;  addr_rom[19111]='h00000000;  wr_data_rom[19111]='h00000000;
    rd_cycle[19112] = 1'b0;  wr_cycle[19112] = 1'b0;  addr_rom[19112]='h00000000;  wr_data_rom[19112]='h00000000;
    rd_cycle[19113] = 1'b0;  wr_cycle[19113] = 1'b0;  addr_rom[19113]='h00000000;  wr_data_rom[19113]='h00000000;
    rd_cycle[19114] = 1'b0;  wr_cycle[19114] = 1'b0;  addr_rom[19114]='h00000000;  wr_data_rom[19114]='h00000000;
    rd_cycle[19115] = 1'b0;  wr_cycle[19115] = 1'b0;  addr_rom[19115]='h00000000;  wr_data_rom[19115]='h00000000;
    rd_cycle[19116] = 1'b0;  wr_cycle[19116] = 1'b0;  addr_rom[19116]='h00000000;  wr_data_rom[19116]='h00000000;
    rd_cycle[19117] = 1'b0;  wr_cycle[19117] = 1'b0;  addr_rom[19117]='h00000000;  wr_data_rom[19117]='h00000000;
    rd_cycle[19118] = 1'b0;  wr_cycle[19118] = 1'b0;  addr_rom[19118]='h00000000;  wr_data_rom[19118]='h00000000;
    rd_cycle[19119] = 1'b0;  wr_cycle[19119] = 1'b0;  addr_rom[19119]='h00000000;  wr_data_rom[19119]='h00000000;
    rd_cycle[19120] = 1'b0;  wr_cycle[19120] = 1'b0;  addr_rom[19120]='h00000000;  wr_data_rom[19120]='h00000000;
    rd_cycle[19121] = 1'b0;  wr_cycle[19121] = 1'b0;  addr_rom[19121]='h00000000;  wr_data_rom[19121]='h00000000;
    rd_cycle[19122] = 1'b0;  wr_cycle[19122] = 1'b0;  addr_rom[19122]='h00000000;  wr_data_rom[19122]='h00000000;
    rd_cycle[19123] = 1'b0;  wr_cycle[19123] = 1'b0;  addr_rom[19123]='h00000000;  wr_data_rom[19123]='h00000000;
    rd_cycle[19124] = 1'b0;  wr_cycle[19124] = 1'b0;  addr_rom[19124]='h00000000;  wr_data_rom[19124]='h00000000;
    rd_cycle[19125] = 1'b0;  wr_cycle[19125] = 1'b0;  addr_rom[19125]='h00000000;  wr_data_rom[19125]='h00000000;
    rd_cycle[19126] = 1'b0;  wr_cycle[19126] = 1'b0;  addr_rom[19126]='h00000000;  wr_data_rom[19126]='h00000000;
    rd_cycle[19127] = 1'b0;  wr_cycle[19127] = 1'b0;  addr_rom[19127]='h00000000;  wr_data_rom[19127]='h00000000;
    rd_cycle[19128] = 1'b0;  wr_cycle[19128] = 1'b0;  addr_rom[19128]='h00000000;  wr_data_rom[19128]='h00000000;
    rd_cycle[19129] = 1'b0;  wr_cycle[19129] = 1'b0;  addr_rom[19129]='h00000000;  wr_data_rom[19129]='h00000000;
    rd_cycle[19130] = 1'b0;  wr_cycle[19130] = 1'b0;  addr_rom[19130]='h00000000;  wr_data_rom[19130]='h00000000;
    rd_cycle[19131] = 1'b0;  wr_cycle[19131] = 1'b0;  addr_rom[19131]='h00000000;  wr_data_rom[19131]='h00000000;
    rd_cycle[19132] = 1'b0;  wr_cycle[19132] = 1'b0;  addr_rom[19132]='h00000000;  wr_data_rom[19132]='h00000000;
    rd_cycle[19133] = 1'b0;  wr_cycle[19133] = 1'b0;  addr_rom[19133]='h00000000;  wr_data_rom[19133]='h00000000;
    rd_cycle[19134] = 1'b0;  wr_cycle[19134] = 1'b0;  addr_rom[19134]='h00000000;  wr_data_rom[19134]='h00000000;
    rd_cycle[19135] = 1'b0;  wr_cycle[19135] = 1'b0;  addr_rom[19135]='h00000000;  wr_data_rom[19135]='h00000000;
    rd_cycle[19136] = 1'b0;  wr_cycle[19136] = 1'b0;  addr_rom[19136]='h00000000;  wr_data_rom[19136]='h00000000;
    rd_cycle[19137] = 1'b0;  wr_cycle[19137] = 1'b0;  addr_rom[19137]='h00000000;  wr_data_rom[19137]='h00000000;
    rd_cycle[19138] = 1'b0;  wr_cycle[19138] = 1'b0;  addr_rom[19138]='h00000000;  wr_data_rom[19138]='h00000000;
    rd_cycle[19139] = 1'b0;  wr_cycle[19139] = 1'b0;  addr_rom[19139]='h00000000;  wr_data_rom[19139]='h00000000;
    rd_cycle[19140] = 1'b0;  wr_cycle[19140] = 1'b0;  addr_rom[19140]='h00000000;  wr_data_rom[19140]='h00000000;
    rd_cycle[19141] = 1'b0;  wr_cycle[19141] = 1'b0;  addr_rom[19141]='h00000000;  wr_data_rom[19141]='h00000000;
    rd_cycle[19142] = 1'b0;  wr_cycle[19142] = 1'b0;  addr_rom[19142]='h00000000;  wr_data_rom[19142]='h00000000;
    rd_cycle[19143] = 1'b0;  wr_cycle[19143] = 1'b0;  addr_rom[19143]='h00000000;  wr_data_rom[19143]='h00000000;
    rd_cycle[19144] = 1'b0;  wr_cycle[19144] = 1'b0;  addr_rom[19144]='h00000000;  wr_data_rom[19144]='h00000000;
    rd_cycle[19145] = 1'b0;  wr_cycle[19145] = 1'b0;  addr_rom[19145]='h00000000;  wr_data_rom[19145]='h00000000;
    rd_cycle[19146] = 1'b0;  wr_cycle[19146] = 1'b0;  addr_rom[19146]='h00000000;  wr_data_rom[19146]='h00000000;
    rd_cycle[19147] = 1'b0;  wr_cycle[19147] = 1'b0;  addr_rom[19147]='h00000000;  wr_data_rom[19147]='h00000000;
    rd_cycle[19148] = 1'b0;  wr_cycle[19148] = 1'b0;  addr_rom[19148]='h00000000;  wr_data_rom[19148]='h00000000;
    rd_cycle[19149] = 1'b0;  wr_cycle[19149] = 1'b0;  addr_rom[19149]='h00000000;  wr_data_rom[19149]='h00000000;
    rd_cycle[19150] = 1'b0;  wr_cycle[19150] = 1'b0;  addr_rom[19150]='h00000000;  wr_data_rom[19150]='h00000000;
    rd_cycle[19151] = 1'b0;  wr_cycle[19151] = 1'b0;  addr_rom[19151]='h00000000;  wr_data_rom[19151]='h00000000;
    rd_cycle[19152] = 1'b0;  wr_cycle[19152] = 1'b0;  addr_rom[19152]='h00000000;  wr_data_rom[19152]='h00000000;
    rd_cycle[19153] = 1'b0;  wr_cycle[19153] = 1'b0;  addr_rom[19153]='h00000000;  wr_data_rom[19153]='h00000000;
    rd_cycle[19154] = 1'b0;  wr_cycle[19154] = 1'b0;  addr_rom[19154]='h00000000;  wr_data_rom[19154]='h00000000;
    rd_cycle[19155] = 1'b0;  wr_cycle[19155] = 1'b0;  addr_rom[19155]='h00000000;  wr_data_rom[19155]='h00000000;
    rd_cycle[19156] = 1'b0;  wr_cycle[19156] = 1'b0;  addr_rom[19156]='h00000000;  wr_data_rom[19156]='h00000000;
    rd_cycle[19157] = 1'b0;  wr_cycle[19157] = 1'b0;  addr_rom[19157]='h00000000;  wr_data_rom[19157]='h00000000;
    rd_cycle[19158] = 1'b0;  wr_cycle[19158] = 1'b0;  addr_rom[19158]='h00000000;  wr_data_rom[19158]='h00000000;
    rd_cycle[19159] = 1'b0;  wr_cycle[19159] = 1'b0;  addr_rom[19159]='h00000000;  wr_data_rom[19159]='h00000000;
    rd_cycle[19160] = 1'b0;  wr_cycle[19160] = 1'b0;  addr_rom[19160]='h00000000;  wr_data_rom[19160]='h00000000;
    rd_cycle[19161] = 1'b0;  wr_cycle[19161] = 1'b0;  addr_rom[19161]='h00000000;  wr_data_rom[19161]='h00000000;
    rd_cycle[19162] = 1'b0;  wr_cycle[19162] = 1'b0;  addr_rom[19162]='h00000000;  wr_data_rom[19162]='h00000000;
    rd_cycle[19163] = 1'b0;  wr_cycle[19163] = 1'b0;  addr_rom[19163]='h00000000;  wr_data_rom[19163]='h00000000;
    rd_cycle[19164] = 1'b0;  wr_cycle[19164] = 1'b0;  addr_rom[19164]='h00000000;  wr_data_rom[19164]='h00000000;
    rd_cycle[19165] = 1'b0;  wr_cycle[19165] = 1'b0;  addr_rom[19165]='h00000000;  wr_data_rom[19165]='h00000000;
    rd_cycle[19166] = 1'b0;  wr_cycle[19166] = 1'b0;  addr_rom[19166]='h00000000;  wr_data_rom[19166]='h00000000;
    rd_cycle[19167] = 1'b0;  wr_cycle[19167] = 1'b0;  addr_rom[19167]='h00000000;  wr_data_rom[19167]='h00000000;
    rd_cycle[19168] = 1'b0;  wr_cycle[19168] = 1'b0;  addr_rom[19168]='h00000000;  wr_data_rom[19168]='h00000000;
    rd_cycle[19169] = 1'b0;  wr_cycle[19169] = 1'b0;  addr_rom[19169]='h00000000;  wr_data_rom[19169]='h00000000;
    rd_cycle[19170] = 1'b0;  wr_cycle[19170] = 1'b0;  addr_rom[19170]='h00000000;  wr_data_rom[19170]='h00000000;
    rd_cycle[19171] = 1'b0;  wr_cycle[19171] = 1'b0;  addr_rom[19171]='h00000000;  wr_data_rom[19171]='h00000000;
    rd_cycle[19172] = 1'b0;  wr_cycle[19172] = 1'b0;  addr_rom[19172]='h00000000;  wr_data_rom[19172]='h00000000;
    rd_cycle[19173] = 1'b0;  wr_cycle[19173] = 1'b0;  addr_rom[19173]='h00000000;  wr_data_rom[19173]='h00000000;
    rd_cycle[19174] = 1'b0;  wr_cycle[19174] = 1'b0;  addr_rom[19174]='h00000000;  wr_data_rom[19174]='h00000000;
    rd_cycle[19175] = 1'b0;  wr_cycle[19175] = 1'b0;  addr_rom[19175]='h00000000;  wr_data_rom[19175]='h00000000;
    rd_cycle[19176] = 1'b0;  wr_cycle[19176] = 1'b0;  addr_rom[19176]='h00000000;  wr_data_rom[19176]='h00000000;
    rd_cycle[19177] = 1'b0;  wr_cycle[19177] = 1'b0;  addr_rom[19177]='h00000000;  wr_data_rom[19177]='h00000000;
    rd_cycle[19178] = 1'b0;  wr_cycle[19178] = 1'b0;  addr_rom[19178]='h00000000;  wr_data_rom[19178]='h00000000;
    rd_cycle[19179] = 1'b0;  wr_cycle[19179] = 1'b0;  addr_rom[19179]='h00000000;  wr_data_rom[19179]='h00000000;
    rd_cycle[19180] = 1'b0;  wr_cycle[19180] = 1'b0;  addr_rom[19180]='h00000000;  wr_data_rom[19180]='h00000000;
    rd_cycle[19181] = 1'b0;  wr_cycle[19181] = 1'b0;  addr_rom[19181]='h00000000;  wr_data_rom[19181]='h00000000;
    rd_cycle[19182] = 1'b0;  wr_cycle[19182] = 1'b0;  addr_rom[19182]='h00000000;  wr_data_rom[19182]='h00000000;
    rd_cycle[19183] = 1'b0;  wr_cycle[19183] = 1'b0;  addr_rom[19183]='h00000000;  wr_data_rom[19183]='h00000000;
    rd_cycle[19184] = 1'b0;  wr_cycle[19184] = 1'b0;  addr_rom[19184]='h00000000;  wr_data_rom[19184]='h00000000;
    rd_cycle[19185] = 1'b0;  wr_cycle[19185] = 1'b0;  addr_rom[19185]='h00000000;  wr_data_rom[19185]='h00000000;
    rd_cycle[19186] = 1'b0;  wr_cycle[19186] = 1'b0;  addr_rom[19186]='h00000000;  wr_data_rom[19186]='h00000000;
    rd_cycle[19187] = 1'b0;  wr_cycle[19187] = 1'b0;  addr_rom[19187]='h00000000;  wr_data_rom[19187]='h00000000;
    rd_cycle[19188] = 1'b0;  wr_cycle[19188] = 1'b0;  addr_rom[19188]='h00000000;  wr_data_rom[19188]='h00000000;
    rd_cycle[19189] = 1'b0;  wr_cycle[19189] = 1'b0;  addr_rom[19189]='h00000000;  wr_data_rom[19189]='h00000000;
    rd_cycle[19190] = 1'b0;  wr_cycle[19190] = 1'b0;  addr_rom[19190]='h00000000;  wr_data_rom[19190]='h00000000;
    rd_cycle[19191] = 1'b0;  wr_cycle[19191] = 1'b0;  addr_rom[19191]='h00000000;  wr_data_rom[19191]='h00000000;
    rd_cycle[19192] = 1'b0;  wr_cycle[19192] = 1'b0;  addr_rom[19192]='h00000000;  wr_data_rom[19192]='h00000000;
    rd_cycle[19193] = 1'b0;  wr_cycle[19193] = 1'b0;  addr_rom[19193]='h00000000;  wr_data_rom[19193]='h00000000;
    rd_cycle[19194] = 1'b0;  wr_cycle[19194] = 1'b0;  addr_rom[19194]='h00000000;  wr_data_rom[19194]='h00000000;
    rd_cycle[19195] = 1'b0;  wr_cycle[19195] = 1'b0;  addr_rom[19195]='h00000000;  wr_data_rom[19195]='h00000000;
    rd_cycle[19196] = 1'b0;  wr_cycle[19196] = 1'b0;  addr_rom[19196]='h00000000;  wr_data_rom[19196]='h00000000;
    rd_cycle[19197] = 1'b0;  wr_cycle[19197] = 1'b0;  addr_rom[19197]='h00000000;  wr_data_rom[19197]='h00000000;
    rd_cycle[19198] = 1'b0;  wr_cycle[19198] = 1'b0;  addr_rom[19198]='h00000000;  wr_data_rom[19198]='h00000000;
    rd_cycle[19199] = 1'b0;  wr_cycle[19199] = 1'b0;  addr_rom[19199]='h00000000;  wr_data_rom[19199]='h00000000;
    rd_cycle[19200] = 1'b0;  wr_cycle[19200] = 1'b0;  addr_rom[19200]='h00000000;  wr_data_rom[19200]='h00000000;
    rd_cycle[19201] = 1'b0;  wr_cycle[19201] = 1'b0;  addr_rom[19201]='h00000000;  wr_data_rom[19201]='h00000000;
    rd_cycle[19202] = 1'b0;  wr_cycle[19202] = 1'b0;  addr_rom[19202]='h00000000;  wr_data_rom[19202]='h00000000;
    rd_cycle[19203] = 1'b0;  wr_cycle[19203] = 1'b0;  addr_rom[19203]='h00000000;  wr_data_rom[19203]='h00000000;
    rd_cycle[19204] = 1'b0;  wr_cycle[19204] = 1'b0;  addr_rom[19204]='h00000000;  wr_data_rom[19204]='h00000000;
    rd_cycle[19205] = 1'b0;  wr_cycle[19205] = 1'b0;  addr_rom[19205]='h00000000;  wr_data_rom[19205]='h00000000;
    rd_cycle[19206] = 1'b0;  wr_cycle[19206] = 1'b0;  addr_rom[19206]='h00000000;  wr_data_rom[19206]='h00000000;
    rd_cycle[19207] = 1'b0;  wr_cycle[19207] = 1'b0;  addr_rom[19207]='h00000000;  wr_data_rom[19207]='h00000000;
    rd_cycle[19208] = 1'b0;  wr_cycle[19208] = 1'b0;  addr_rom[19208]='h00000000;  wr_data_rom[19208]='h00000000;
    rd_cycle[19209] = 1'b0;  wr_cycle[19209] = 1'b0;  addr_rom[19209]='h00000000;  wr_data_rom[19209]='h00000000;
    rd_cycle[19210] = 1'b0;  wr_cycle[19210] = 1'b0;  addr_rom[19210]='h00000000;  wr_data_rom[19210]='h00000000;
    rd_cycle[19211] = 1'b0;  wr_cycle[19211] = 1'b0;  addr_rom[19211]='h00000000;  wr_data_rom[19211]='h00000000;
    rd_cycle[19212] = 1'b0;  wr_cycle[19212] = 1'b0;  addr_rom[19212]='h00000000;  wr_data_rom[19212]='h00000000;
    rd_cycle[19213] = 1'b0;  wr_cycle[19213] = 1'b0;  addr_rom[19213]='h00000000;  wr_data_rom[19213]='h00000000;
    rd_cycle[19214] = 1'b0;  wr_cycle[19214] = 1'b0;  addr_rom[19214]='h00000000;  wr_data_rom[19214]='h00000000;
    rd_cycle[19215] = 1'b0;  wr_cycle[19215] = 1'b0;  addr_rom[19215]='h00000000;  wr_data_rom[19215]='h00000000;
    rd_cycle[19216] = 1'b0;  wr_cycle[19216] = 1'b0;  addr_rom[19216]='h00000000;  wr_data_rom[19216]='h00000000;
    rd_cycle[19217] = 1'b0;  wr_cycle[19217] = 1'b0;  addr_rom[19217]='h00000000;  wr_data_rom[19217]='h00000000;
    rd_cycle[19218] = 1'b0;  wr_cycle[19218] = 1'b0;  addr_rom[19218]='h00000000;  wr_data_rom[19218]='h00000000;
    rd_cycle[19219] = 1'b0;  wr_cycle[19219] = 1'b0;  addr_rom[19219]='h00000000;  wr_data_rom[19219]='h00000000;
    rd_cycle[19220] = 1'b0;  wr_cycle[19220] = 1'b0;  addr_rom[19220]='h00000000;  wr_data_rom[19220]='h00000000;
    rd_cycle[19221] = 1'b0;  wr_cycle[19221] = 1'b0;  addr_rom[19221]='h00000000;  wr_data_rom[19221]='h00000000;
    rd_cycle[19222] = 1'b0;  wr_cycle[19222] = 1'b0;  addr_rom[19222]='h00000000;  wr_data_rom[19222]='h00000000;
    rd_cycle[19223] = 1'b0;  wr_cycle[19223] = 1'b0;  addr_rom[19223]='h00000000;  wr_data_rom[19223]='h00000000;
    rd_cycle[19224] = 1'b0;  wr_cycle[19224] = 1'b0;  addr_rom[19224]='h00000000;  wr_data_rom[19224]='h00000000;
    rd_cycle[19225] = 1'b0;  wr_cycle[19225] = 1'b0;  addr_rom[19225]='h00000000;  wr_data_rom[19225]='h00000000;
    rd_cycle[19226] = 1'b0;  wr_cycle[19226] = 1'b0;  addr_rom[19226]='h00000000;  wr_data_rom[19226]='h00000000;
    rd_cycle[19227] = 1'b0;  wr_cycle[19227] = 1'b0;  addr_rom[19227]='h00000000;  wr_data_rom[19227]='h00000000;
    rd_cycle[19228] = 1'b0;  wr_cycle[19228] = 1'b0;  addr_rom[19228]='h00000000;  wr_data_rom[19228]='h00000000;
    rd_cycle[19229] = 1'b0;  wr_cycle[19229] = 1'b0;  addr_rom[19229]='h00000000;  wr_data_rom[19229]='h00000000;
    rd_cycle[19230] = 1'b0;  wr_cycle[19230] = 1'b0;  addr_rom[19230]='h00000000;  wr_data_rom[19230]='h00000000;
    rd_cycle[19231] = 1'b0;  wr_cycle[19231] = 1'b0;  addr_rom[19231]='h00000000;  wr_data_rom[19231]='h00000000;
    rd_cycle[19232] = 1'b0;  wr_cycle[19232] = 1'b0;  addr_rom[19232]='h00000000;  wr_data_rom[19232]='h00000000;
    rd_cycle[19233] = 1'b0;  wr_cycle[19233] = 1'b0;  addr_rom[19233]='h00000000;  wr_data_rom[19233]='h00000000;
    rd_cycle[19234] = 1'b0;  wr_cycle[19234] = 1'b0;  addr_rom[19234]='h00000000;  wr_data_rom[19234]='h00000000;
    rd_cycle[19235] = 1'b0;  wr_cycle[19235] = 1'b0;  addr_rom[19235]='h00000000;  wr_data_rom[19235]='h00000000;
    rd_cycle[19236] = 1'b0;  wr_cycle[19236] = 1'b0;  addr_rom[19236]='h00000000;  wr_data_rom[19236]='h00000000;
    rd_cycle[19237] = 1'b0;  wr_cycle[19237] = 1'b0;  addr_rom[19237]='h00000000;  wr_data_rom[19237]='h00000000;
    rd_cycle[19238] = 1'b0;  wr_cycle[19238] = 1'b0;  addr_rom[19238]='h00000000;  wr_data_rom[19238]='h00000000;
    rd_cycle[19239] = 1'b0;  wr_cycle[19239] = 1'b0;  addr_rom[19239]='h00000000;  wr_data_rom[19239]='h00000000;
    rd_cycle[19240] = 1'b0;  wr_cycle[19240] = 1'b0;  addr_rom[19240]='h00000000;  wr_data_rom[19240]='h00000000;
    rd_cycle[19241] = 1'b0;  wr_cycle[19241] = 1'b0;  addr_rom[19241]='h00000000;  wr_data_rom[19241]='h00000000;
    rd_cycle[19242] = 1'b0;  wr_cycle[19242] = 1'b0;  addr_rom[19242]='h00000000;  wr_data_rom[19242]='h00000000;
    rd_cycle[19243] = 1'b0;  wr_cycle[19243] = 1'b0;  addr_rom[19243]='h00000000;  wr_data_rom[19243]='h00000000;
    rd_cycle[19244] = 1'b0;  wr_cycle[19244] = 1'b0;  addr_rom[19244]='h00000000;  wr_data_rom[19244]='h00000000;
    rd_cycle[19245] = 1'b0;  wr_cycle[19245] = 1'b0;  addr_rom[19245]='h00000000;  wr_data_rom[19245]='h00000000;
    rd_cycle[19246] = 1'b0;  wr_cycle[19246] = 1'b0;  addr_rom[19246]='h00000000;  wr_data_rom[19246]='h00000000;
    rd_cycle[19247] = 1'b0;  wr_cycle[19247] = 1'b0;  addr_rom[19247]='h00000000;  wr_data_rom[19247]='h00000000;
    rd_cycle[19248] = 1'b0;  wr_cycle[19248] = 1'b0;  addr_rom[19248]='h00000000;  wr_data_rom[19248]='h00000000;
    rd_cycle[19249] = 1'b0;  wr_cycle[19249] = 1'b0;  addr_rom[19249]='h00000000;  wr_data_rom[19249]='h00000000;
    rd_cycle[19250] = 1'b0;  wr_cycle[19250] = 1'b0;  addr_rom[19250]='h00000000;  wr_data_rom[19250]='h00000000;
    rd_cycle[19251] = 1'b0;  wr_cycle[19251] = 1'b0;  addr_rom[19251]='h00000000;  wr_data_rom[19251]='h00000000;
    rd_cycle[19252] = 1'b0;  wr_cycle[19252] = 1'b0;  addr_rom[19252]='h00000000;  wr_data_rom[19252]='h00000000;
    rd_cycle[19253] = 1'b0;  wr_cycle[19253] = 1'b0;  addr_rom[19253]='h00000000;  wr_data_rom[19253]='h00000000;
    rd_cycle[19254] = 1'b0;  wr_cycle[19254] = 1'b0;  addr_rom[19254]='h00000000;  wr_data_rom[19254]='h00000000;
    rd_cycle[19255] = 1'b0;  wr_cycle[19255] = 1'b0;  addr_rom[19255]='h00000000;  wr_data_rom[19255]='h00000000;
    rd_cycle[19256] = 1'b0;  wr_cycle[19256] = 1'b0;  addr_rom[19256]='h00000000;  wr_data_rom[19256]='h00000000;
    rd_cycle[19257] = 1'b0;  wr_cycle[19257] = 1'b0;  addr_rom[19257]='h00000000;  wr_data_rom[19257]='h00000000;
    rd_cycle[19258] = 1'b0;  wr_cycle[19258] = 1'b0;  addr_rom[19258]='h00000000;  wr_data_rom[19258]='h00000000;
    rd_cycle[19259] = 1'b0;  wr_cycle[19259] = 1'b0;  addr_rom[19259]='h00000000;  wr_data_rom[19259]='h00000000;
    rd_cycle[19260] = 1'b0;  wr_cycle[19260] = 1'b0;  addr_rom[19260]='h00000000;  wr_data_rom[19260]='h00000000;
    rd_cycle[19261] = 1'b0;  wr_cycle[19261] = 1'b0;  addr_rom[19261]='h00000000;  wr_data_rom[19261]='h00000000;
    rd_cycle[19262] = 1'b0;  wr_cycle[19262] = 1'b0;  addr_rom[19262]='h00000000;  wr_data_rom[19262]='h00000000;
    rd_cycle[19263] = 1'b0;  wr_cycle[19263] = 1'b0;  addr_rom[19263]='h00000000;  wr_data_rom[19263]='h00000000;
    rd_cycle[19264] = 1'b0;  wr_cycle[19264] = 1'b0;  addr_rom[19264]='h00000000;  wr_data_rom[19264]='h00000000;
    rd_cycle[19265] = 1'b0;  wr_cycle[19265] = 1'b0;  addr_rom[19265]='h00000000;  wr_data_rom[19265]='h00000000;
    rd_cycle[19266] = 1'b0;  wr_cycle[19266] = 1'b0;  addr_rom[19266]='h00000000;  wr_data_rom[19266]='h00000000;
    rd_cycle[19267] = 1'b0;  wr_cycle[19267] = 1'b0;  addr_rom[19267]='h00000000;  wr_data_rom[19267]='h00000000;
    rd_cycle[19268] = 1'b0;  wr_cycle[19268] = 1'b0;  addr_rom[19268]='h00000000;  wr_data_rom[19268]='h00000000;
    rd_cycle[19269] = 1'b0;  wr_cycle[19269] = 1'b0;  addr_rom[19269]='h00000000;  wr_data_rom[19269]='h00000000;
    rd_cycle[19270] = 1'b0;  wr_cycle[19270] = 1'b0;  addr_rom[19270]='h00000000;  wr_data_rom[19270]='h00000000;
    rd_cycle[19271] = 1'b0;  wr_cycle[19271] = 1'b0;  addr_rom[19271]='h00000000;  wr_data_rom[19271]='h00000000;
    rd_cycle[19272] = 1'b0;  wr_cycle[19272] = 1'b0;  addr_rom[19272]='h00000000;  wr_data_rom[19272]='h00000000;
    rd_cycle[19273] = 1'b0;  wr_cycle[19273] = 1'b0;  addr_rom[19273]='h00000000;  wr_data_rom[19273]='h00000000;
    rd_cycle[19274] = 1'b0;  wr_cycle[19274] = 1'b0;  addr_rom[19274]='h00000000;  wr_data_rom[19274]='h00000000;
    rd_cycle[19275] = 1'b0;  wr_cycle[19275] = 1'b0;  addr_rom[19275]='h00000000;  wr_data_rom[19275]='h00000000;
    rd_cycle[19276] = 1'b0;  wr_cycle[19276] = 1'b0;  addr_rom[19276]='h00000000;  wr_data_rom[19276]='h00000000;
    rd_cycle[19277] = 1'b0;  wr_cycle[19277] = 1'b0;  addr_rom[19277]='h00000000;  wr_data_rom[19277]='h00000000;
    rd_cycle[19278] = 1'b0;  wr_cycle[19278] = 1'b0;  addr_rom[19278]='h00000000;  wr_data_rom[19278]='h00000000;
    rd_cycle[19279] = 1'b0;  wr_cycle[19279] = 1'b0;  addr_rom[19279]='h00000000;  wr_data_rom[19279]='h00000000;
    rd_cycle[19280] = 1'b0;  wr_cycle[19280] = 1'b0;  addr_rom[19280]='h00000000;  wr_data_rom[19280]='h00000000;
    rd_cycle[19281] = 1'b0;  wr_cycle[19281] = 1'b0;  addr_rom[19281]='h00000000;  wr_data_rom[19281]='h00000000;
    rd_cycle[19282] = 1'b0;  wr_cycle[19282] = 1'b0;  addr_rom[19282]='h00000000;  wr_data_rom[19282]='h00000000;
    rd_cycle[19283] = 1'b0;  wr_cycle[19283] = 1'b0;  addr_rom[19283]='h00000000;  wr_data_rom[19283]='h00000000;
    rd_cycle[19284] = 1'b0;  wr_cycle[19284] = 1'b0;  addr_rom[19284]='h00000000;  wr_data_rom[19284]='h00000000;
    rd_cycle[19285] = 1'b0;  wr_cycle[19285] = 1'b0;  addr_rom[19285]='h00000000;  wr_data_rom[19285]='h00000000;
    rd_cycle[19286] = 1'b0;  wr_cycle[19286] = 1'b0;  addr_rom[19286]='h00000000;  wr_data_rom[19286]='h00000000;
    rd_cycle[19287] = 1'b0;  wr_cycle[19287] = 1'b0;  addr_rom[19287]='h00000000;  wr_data_rom[19287]='h00000000;
    rd_cycle[19288] = 1'b0;  wr_cycle[19288] = 1'b0;  addr_rom[19288]='h00000000;  wr_data_rom[19288]='h00000000;
    rd_cycle[19289] = 1'b0;  wr_cycle[19289] = 1'b0;  addr_rom[19289]='h00000000;  wr_data_rom[19289]='h00000000;
    rd_cycle[19290] = 1'b0;  wr_cycle[19290] = 1'b0;  addr_rom[19290]='h00000000;  wr_data_rom[19290]='h00000000;
    rd_cycle[19291] = 1'b0;  wr_cycle[19291] = 1'b0;  addr_rom[19291]='h00000000;  wr_data_rom[19291]='h00000000;
    rd_cycle[19292] = 1'b0;  wr_cycle[19292] = 1'b0;  addr_rom[19292]='h00000000;  wr_data_rom[19292]='h00000000;
    rd_cycle[19293] = 1'b0;  wr_cycle[19293] = 1'b0;  addr_rom[19293]='h00000000;  wr_data_rom[19293]='h00000000;
    rd_cycle[19294] = 1'b0;  wr_cycle[19294] = 1'b0;  addr_rom[19294]='h00000000;  wr_data_rom[19294]='h00000000;
    rd_cycle[19295] = 1'b0;  wr_cycle[19295] = 1'b0;  addr_rom[19295]='h00000000;  wr_data_rom[19295]='h00000000;
    rd_cycle[19296] = 1'b0;  wr_cycle[19296] = 1'b0;  addr_rom[19296]='h00000000;  wr_data_rom[19296]='h00000000;
    rd_cycle[19297] = 1'b0;  wr_cycle[19297] = 1'b0;  addr_rom[19297]='h00000000;  wr_data_rom[19297]='h00000000;
    rd_cycle[19298] = 1'b0;  wr_cycle[19298] = 1'b0;  addr_rom[19298]='h00000000;  wr_data_rom[19298]='h00000000;
    rd_cycle[19299] = 1'b0;  wr_cycle[19299] = 1'b0;  addr_rom[19299]='h00000000;  wr_data_rom[19299]='h00000000;
    rd_cycle[19300] = 1'b0;  wr_cycle[19300] = 1'b0;  addr_rom[19300]='h00000000;  wr_data_rom[19300]='h00000000;
    rd_cycle[19301] = 1'b0;  wr_cycle[19301] = 1'b0;  addr_rom[19301]='h00000000;  wr_data_rom[19301]='h00000000;
    rd_cycle[19302] = 1'b0;  wr_cycle[19302] = 1'b0;  addr_rom[19302]='h00000000;  wr_data_rom[19302]='h00000000;
    rd_cycle[19303] = 1'b0;  wr_cycle[19303] = 1'b0;  addr_rom[19303]='h00000000;  wr_data_rom[19303]='h00000000;
    rd_cycle[19304] = 1'b0;  wr_cycle[19304] = 1'b0;  addr_rom[19304]='h00000000;  wr_data_rom[19304]='h00000000;
    rd_cycle[19305] = 1'b0;  wr_cycle[19305] = 1'b0;  addr_rom[19305]='h00000000;  wr_data_rom[19305]='h00000000;
    rd_cycle[19306] = 1'b0;  wr_cycle[19306] = 1'b0;  addr_rom[19306]='h00000000;  wr_data_rom[19306]='h00000000;
    rd_cycle[19307] = 1'b0;  wr_cycle[19307] = 1'b0;  addr_rom[19307]='h00000000;  wr_data_rom[19307]='h00000000;
    rd_cycle[19308] = 1'b0;  wr_cycle[19308] = 1'b0;  addr_rom[19308]='h00000000;  wr_data_rom[19308]='h00000000;
    rd_cycle[19309] = 1'b0;  wr_cycle[19309] = 1'b0;  addr_rom[19309]='h00000000;  wr_data_rom[19309]='h00000000;
    rd_cycle[19310] = 1'b0;  wr_cycle[19310] = 1'b0;  addr_rom[19310]='h00000000;  wr_data_rom[19310]='h00000000;
    rd_cycle[19311] = 1'b0;  wr_cycle[19311] = 1'b0;  addr_rom[19311]='h00000000;  wr_data_rom[19311]='h00000000;
    rd_cycle[19312] = 1'b0;  wr_cycle[19312] = 1'b0;  addr_rom[19312]='h00000000;  wr_data_rom[19312]='h00000000;
    rd_cycle[19313] = 1'b0;  wr_cycle[19313] = 1'b0;  addr_rom[19313]='h00000000;  wr_data_rom[19313]='h00000000;
    rd_cycle[19314] = 1'b0;  wr_cycle[19314] = 1'b0;  addr_rom[19314]='h00000000;  wr_data_rom[19314]='h00000000;
    rd_cycle[19315] = 1'b0;  wr_cycle[19315] = 1'b0;  addr_rom[19315]='h00000000;  wr_data_rom[19315]='h00000000;
    rd_cycle[19316] = 1'b0;  wr_cycle[19316] = 1'b0;  addr_rom[19316]='h00000000;  wr_data_rom[19316]='h00000000;
    rd_cycle[19317] = 1'b0;  wr_cycle[19317] = 1'b0;  addr_rom[19317]='h00000000;  wr_data_rom[19317]='h00000000;
    rd_cycle[19318] = 1'b0;  wr_cycle[19318] = 1'b0;  addr_rom[19318]='h00000000;  wr_data_rom[19318]='h00000000;
    rd_cycle[19319] = 1'b0;  wr_cycle[19319] = 1'b0;  addr_rom[19319]='h00000000;  wr_data_rom[19319]='h00000000;
    rd_cycle[19320] = 1'b0;  wr_cycle[19320] = 1'b0;  addr_rom[19320]='h00000000;  wr_data_rom[19320]='h00000000;
    rd_cycle[19321] = 1'b0;  wr_cycle[19321] = 1'b0;  addr_rom[19321]='h00000000;  wr_data_rom[19321]='h00000000;
    rd_cycle[19322] = 1'b0;  wr_cycle[19322] = 1'b0;  addr_rom[19322]='h00000000;  wr_data_rom[19322]='h00000000;
    rd_cycle[19323] = 1'b0;  wr_cycle[19323] = 1'b0;  addr_rom[19323]='h00000000;  wr_data_rom[19323]='h00000000;
    rd_cycle[19324] = 1'b0;  wr_cycle[19324] = 1'b0;  addr_rom[19324]='h00000000;  wr_data_rom[19324]='h00000000;
    rd_cycle[19325] = 1'b0;  wr_cycle[19325] = 1'b0;  addr_rom[19325]='h00000000;  wr_data_rom[19325]='h00000000;
    rd_cycle[19326] = 1'b0;  wr_cycle[19326] = 1'b0;  addr_rom[19326]='h00000000;  wr_data_rom[19326]='h00000000;
    rd_cycle[19327] = 1'b0;  wr_cycle[19327] = 1'b0;  addr_rom[19327]='h00000000;  wr_data_rom[19327]='h00000000;
    rd_cycle[19328] = 1'b0;  wr_cycle[19328] = 1'b0;  addr_rom[19328]='h00000000;  wr_data_rom[19328]='h00000000;
    rd_cycle[19329] = 1'b0;  wr_cycle[19329] = 1'b0;  addr_rom[19329]='h00000000;  wr_data_rom[19329]='h00000000;
    rd_cycle[19330] = 1'b0;  wr_cycle[19330] = 1'b0;  addr_rom[19330]='h00000000;  wr_data_rom[19330]='h00000000;
    rd_cycle[19331] = 1'b0;  wr_cycle[19331] = 1'b0;  addr_rom[19331]='h00000000;  wr_data_rom[19331]='h00000000;
    rd_cycle[19332] = 1'b0;  wr_cycle[19332] = 1'b0;  addr_rom[19332]='h00000000;  wr_data_rom[19332]='h00000000;
    rd_cycle[19333] = 1'b0;  wr_cycle[19333] = 1'b0;  addr_rom[19333]='h00000000;  wr_data_rom[19333]='h00000000;
    rd_cycle[19334] = 1'b0;  wr_cycle[19334] = 1'b0;  addr_rom[19334]='h00000000;  wr_data_rom[19334]='h00000000;
    rd_cycle[19335] = 1'b0;  wr_cycle[19335] = 1'b0;  addr_rom[19335]='h00000000;  wr_data_rom[19335]='h00000000;
    rd_cycle[19336] = 1'b0;  wr_cycle[19336] = 1'b0;  addr_rom[19336]='h00000000;  wr_data_rom[19336]='h00000000;
    rd_cycle[19337] = 1'b0;  wr_cycle[19337] = 1'b0;  addr_rom[19337]='h00000000;  wr_data_rom[19337]='h00000000;
    rd_cycle[19338] = 1'b0;  wr_cycle[19338] = 1'b0;  addr_rom[19338]='h00000000;  wr_data_rom[19338]='h00000000;
    rd_cycle[19339] = 1'b0;  wr_cycle[19339] = 1'b0;  addr_rom[19339]='h00000000;  wr_data_rom[19339]='h00000000;
    rd_cycle[19340] = 1'b0;  wr_cycle[19340] = 1'b0;  addr_rom[19340]='h00000000;  wr_data_rom[19340]='h00000000;
    rd_cycle[19341] = 1'b0;  wr_cycle[19341] = 1'b0;  addr_rom[19341]='h00000000;  wr_data_rom[19341]='h00000000;
    rd_cycle[19342] = 1'b0;  wr_cycle[19342] = 1'b0;  addr_rom[19342]='h00000000;  wr_data_rom[19342]='h00000000;
    rd_cycle[19343] = 1'b0;  wr_cycle[19343] = 1'b0;  addr_rom[19343]='h00000000;  wr_data_rom[19343]='h00000000;
    rd_cycle[19344] = 1'b0;  wr_cycle[19344] = 1'b0;  addr_rom[19344]='h00000000;  wr_data_rom[19344]='h00000000;
    rd_cycle[19345] = 1'b0;  wr_cycle[19345] = 1'b0;  addr_rom[19345]='h00000000;  wr_data_rom[19345]='h00000000;
    rd_cycle[19346] = 1'b0;  wr_cycle[19346] = 1'b0;  addr_rom[19346]='h00000000;  wr_data_rom[19346]='h00000000;
    rd_cycle[19347] = 1'b0;  wr_cycle[19347] = 1'b0;  addr_rom[19347]='h00000000;  wr_data_rom[19347]='h00000000;
    rd_cycle[19348] = 1'b0;  wr_cycle[19348] = 1'b0;  addr_rom[19348]='h00000000;  wr_data_rom[19348]='h00000000;
    rd_cycle[19349] = 1'b0;  wr_cycle[19349] = 1'b0;  addr_rom[19349]='h00000000;  wr_data_rom[19349]='h00000000;
    rd_cycle[19350] = 1'b0;  wr_cycle[19350] = 1'b0;  addr_rom[19350]='h00000000;  wr_data_rom[19350]='h00000000;
    rd_cycle[19351] = 1'b0;  wr_cycle[19351] = 1'b0;  addr_rom[19351]='h00000000;  wr_data_rom[19351]='h00000000;
    rd_cycle[19352] = 1'b0;  wr_cycle[19352] = 1'b0;  addr_rom[19352]='h00000000;  wr_data_rom[19352]='h00000000;
    rd_cycle[19353] = 1'b0;  wr_cycle[19353] = 1'b0;  addr_rom[19353]='h00000000;  wr_data_rom[19353]='h00000000;
    rd_cycle[19354] = 1'b0;  wr_cycle[19354] = 1'b0;  addr_rom[19354]='h00000000;  wr_data_rom[19354]='h00000000;
    rd_cycle[19355] = 1'b0;  wr_cycle[19355] = 1'b0;  addr_rom[19355]='h00000000;  wr_data_rom[19355]='h00000000;
    rd_cycle[19356] = 1'b0;  wr_cycle[19356] = 1'b0;  addr_rom[19356]='h00000000;  wr_data_rom[19356]='h00000000;
    rd_cycle[19357] = 1'b0;  wr_cycle[19357] = 1'b0;  addr_rom[19357]='h00000000;  wr_data_rom[19357]='h00000000;
    rd_cycle[19358] = 1'b0;  wr_cycle[19358] = 1'b0;  addr_rom[19358]='h00000000;  wr_data_rom[19358]='h00000000;
    rd_cycle[19359] = 1'b0;  wr_cycle[19359] = 1'b0;  addr_rom[19359]='h00000000;  wr_data_rom[19359]='h00000000;
    rd_cycle[19360] = 1'b0;  wr_cycle[19360] = 1'b0;  addr_rom[19360]='h00000000;  wr_data_rom[19360]='h00000000;
    rd_cycle[19361] = 1'b0;  wr_cycle[19361] = 1'b0;  addr_rom[19361]='h00000000;  wr_data_rom[19361]='h00000000;
    rd_cycle[19362] = 1'b0;  wr_cycle[19362] = 1'b0;  addr_rom[19362]='h00000000;  wr_data_rom[19362]='h00000000;
    rd_cycle[19363] = 1'b0;  wr_cycle[19363] = 1'b0;  addr_rom[19363]='h00000000;  wr_data_rom[19363]='h00000000;
    rd_cycle[19364] = 1'b0;  wr_cycle[19364] = 1'b0;  addr_rom[19364]='h00000000;  wr_data_rom[19364]='h00000000;
    rd_cycle[19365] = 1'b0;  wr_cycle[19365] = 1'b0;  addr_rom[19365]='h00000000;  wr_data_rom[19365]='h00000000;
    rd_cycle[19366] = 1'b0;  wr_cycle[19366] = 1'b0;  addr_rom[19366]='h00000000;  wr_data_rom[19366]='h00000000;
    rd_cycle[19367] = 1'b0;  wr_cycle[19367] = 1'b0;  addr_rom[19367]='h00000000;  wr_data_rom[19367]='h00000000;
    rd_cycle[19368] = 1'b0;  wr_cycle[19368] = 1'b0;  addr_rom[19368]='h00000000;  wr_data_rom[19368]='h00000000;
    rd_cycle[19369] = 1'b0;  wr_cycle[19369] = 1'b0;  addr_rom[19369]='h00000000;  wr_data_rom[19369]='h00000000;
    rd_cycle[19370] = 1'b0;  wr_cycle[19370] = 1'b0;  addr_rom[19370]='h00000000;  wr_data_rom[19370]='h00000000;
    rd_cycle[19371] = 1'b0;  wr_cycle[19371] = 1'b0;  addr_rom[19371]='h00000000;  wr_data_rom[19371]='h00000000;
    rd_cycle[19372] = 1'b0;  wr_cycle[19372] = 1'b0;  addr_rom[19372]='h00000000;  wr_data_rom[19372]='h00000000;
    rd_cycle[19373] = 1'b0;  wr_cycle[19373] = 1'b0;  addr_rom[19373]='h00000000;  wr_data_rom[19373]='h00000000;
    rd_cycle[19374] = 1'b0;  wr_cycle[19374] = 1'b0;  addr_rom[19374]='h00000000;  wr_data_rom[19374]='h00000000;
    rd_cycle[19375] = 1'b0;  wr_cycle[19375] = 1'b0;  addr_rom[19375]='h00000000;  wr_data_rom[19375]='h00000000;
    rd_cycle[19376] = 1'b0;  wr_cycle[19376] = 1'b0;  addr_rom[19376]='h00000000;  wr_data_rom[19376]='h00000000;
    rd_cycle[19377] = 1'b0;  wr_cycle[19377] = 1'b0;  addr_rom[19377]='h00000000;  wr_data_rom[19377]='h00000000;
    rd_cycle[19378] = 1'b0;  wr_cycle[19378] = 1'b0;  addr_rom[19378]='h00000000;  wr_data_rom[19378]='h00000000;
    rd_cycle[19379] = 1'b0;  wr_cycle[19379] = 1'b0;  addr_rom[19379]='h00000000;  wr_data_rom[19379]='h00000000;
    rd_cycle[19380] = 1'b0;  wr_cycle[19380] = 1'b0;  addr_rom[19380]='h00000000;  wr_data_rom[19380]='h00000000;
    rd_cycle[19381] = 1'b0;  wr_cycle[19381] = 1'b0;  addr_rom[19381]='h00000000;  wr_data_rom[19381]='h00000000;
    rd_cycle[19382] = 1'b0;  wr_cycle[19382] = 1'b0;  addr_rom[19382]='h00000000;  wr_data_rom[19382]='h00000000;
    rd_cycle[19383] = 1'b0;  wr_cycle[19383] = 1'b0;  addr_rom[19383]='h00000000;  wr_data_rom[19383]='h00000000;
    rd_cycle[19384] = 1'b0;  wr_cycle[19384] = 1'b0;  addr_rom[19384]='h00000000;  wr_data_rom[19384]='h00000000;
    rd_cycle[19385] = 1'b0;  wr_cycle[19385] = 1'b0;  addr_rom[19385]='h00000000;  wr_data_rom[19385]='h00000000;
    rd_cycle[19386] = 1'b0;  wr_cycle[19386] = 1'b0;  addr_rom[19386]='h00000000;  wr_data_rom[19386]='h00000000;
    rd_cycle[19387] = 1'b0;  wr_cycle[19387] = 1'b0;  addr_rom[19387]='h00000000;  wr_data_rom[19387]='h00000000;
    rd_cycle[19388] = 1'b0;  wr_cycle[19388] = 1'b0;  addr_rom[19388]='h00000000;  wr_data_rom[19388]='h00000000;
    rd_cycle[19389] = 1'b0;  wr_cycle[19389] = 1'b0;  addr_rom[19389]='h00000000;  wr_data_rom[19389]='h00000000;
    rd_cycle[19390] = 1'b0;  wr_cycle[19390] = 1'b0;  addr_rom[19390]='h00000000;  wr_data_rom[19390]='h00000000;
    rd_cycle[19391] = 1'b0;  wr_cycle[19391] = 1'b0;  addr_rom[19391]='h00000000;  wr_data_rom[19391]='h00000000;
    rd_cycle[19392] = 1'b0;  wr_cycle[19392] = 1'b0;  addr_rom[19392]='h00000000;  wr_data_rom[19392]='h00000000;
    rd_cycle[19393] = 1'b0;  wr_cycle[19393] = 1'b0;  addr_rom[19393]='h00000000;  wr_data_rom[19393]='h00000000;
    rd_cycle[19394] = 1'b0;  wr_cycle[19394] = 1'b0;  addr_rom[19394]='h00000000;  wr_data_rom[19394]='h00000000;
    rd_cycle[19395] = 1'b0;  wr_cycle[19395] = 1'b0;  addr_rom[19395]='h00000000;  wr_data_rom[19395]='h00000000;
    rd_cycle[19396] = 1'b0;  wr_cycle[19396] = 1'b0;  addr_rom[19396]='h00000000;  wr_data_rom[19396]='h00000000;
    rd_cycle[19397] = 1'b0;  wr_cycle[19397] = 1'b0;  addr_rom[19397]='h00000000;  wr_data_rom[19397]='h00000000;
    rd_cycle[19398] = 1'b0;  wr_cycle[19398] = 1'b0;  addr_rom[19398]='h00000000;  wr_data_rom[19398]='h00000000;
    rd_cycle[19399] = 1'b0;  wr_cycle[19399] = 1'b0;  addr_rom[19399]='h00000000;  wr_data_rom[19399]='h00000000;
    rd_cycle[19400] = 1'b0;  wr_cycle[19400] = 1'b0;  addr_rom[19400]='h00000000;  wr_data_rom[19400]='h00000000;
    rd_cycle[19401] = 1'b0;  wr_cycle[19401] = 1'b0;  addr_rom[19401]='h00000000;  wr_data_rom[19401]='h00000000;
    rd_cycle[19402] = 1'b0;  wr_cycle[19402] = 1'b0;  addr_rom[19402]='h00000000;  wr_data_rom[19402]='h00000000;
    rd_cycle[19403] = 1'b0;  wr_cycle[19403] = 1'b0;  addr_rom[19403]='h00000000;  wr_data_rom[19403]='h00000000;
    rd_cycle[19404] = 1'b0;  wr_cycle[19404] = 1'b0;  addr_rom[19404]='h00000000;  wr_data_rom[19404]='h00000000;
    rd_cycle[19405] = 1'b0;  wr_cycle[19405] = 1'b0;  addr_rom[19405]='h00000000;  wr_data_rom[19405]='h00000000;
    rd_cycle[19406] = 1'b0;  wr_cycle[19406] = 1'b0;  addr_rom[19406]='h00000000;  wr_data_rom[19406]='h00000000;
    rd_cycle[19407] = 1'b0;  wr_cycle[19407] = 1'b0;  addr_rom[19407]='h00000000;  wr_data_rom[19407]='h00000000;
    rd_cycle[19408] = 1'b0;  wr_cycle[19408] = 1'b0;  addr_rom[19408]='h00000000;  wr_data_rom[19408]='h00000000;
    rd_cycle[19409] = 1'b0;  wr_cycle[19409] = 1'b0;  addr_rom[19409]='h00000000;  wr_data_rom[19409]='h00000000;
    rd_cycle[19410] = 1'b0;  wr_cycle[19410] = 1'b0;  addr_rom[19410]='h00000000;  wr_data_rom[19410]='h00000000;
    rd_cycle[19411] = 1'b0;  wr_cycle[19411] = 1'b0;  addr_rom[19411]='h00000000;  wr_data_rom[19411]='h00000000;
    rd_cycle[19412] = 1'b0;  wr_cycle[19412] = 1'b0;  addr_rom[19412]='h00000000;  wr_data_rom[19412]='h00000000;
    rd_cycle[19413] = 1'b0;  wr_cycle[19413] = 1'b0;  addr_rom[19413]='h00000000;  wr_data_rom[19413]='h00000000;
    rd_cycle[19414] = 1'b0;  wr_cycle[19414] = 1'b0;  addr_rom[19414]='h00000000;  wr_data_rom[19414]='h00000000;
    rd_cycle[19415] = 1'b0;  wr_cycle[19415] = 1'b0;  addr_rom[19415]='h00000000;  wr_data_rom[19415]='h00000000;
    rd_cycle[19416] = 1'b0;  wr_cycle[19416] = 1'b0;  addr_rom[19416]='h00000000;  wr_data_rom[19416]='h00000000;
    rd_cycle[19417] = 1'b0;  wr_cycle[19417] = 1'b0;  addr_rom[19417]='h00000000;  wr_data_rom[19417]='h00000000;
    rd_cycle[19418] = 1'b0;  wr_cycle[19418] = 1'b0;  addr_rom[19418]='h00000000;  wr_data_rom[19418]='h00000000;
    rd_cycle[19419] = 1'b0;  wr_cycle[19419] = 1'b0;  addr_rom[19419]='h00000000;  wr_data_rom[19419]='h00000000;
    rd_cycle[19420] = 1'b0;  wr_cycle[19420] = 1'b0;  addr_rom[19420]='h00000000;  wr_data_rom[19420]='h00000000;
    rd_cycle[19421] = 1'b0;  wr_cycle[19421] = 1'b0;  addr_rom[19421]='h00000000;  wr_data_rom[19421]='h00000000;
    rd_cycle[19422] = 1'b0;  wr_cycle[19422] = 1'b0;  addr_rom[19422]='h00000000;  wr_data_rom[19422]='h00000000;
    rd_cycle[19423] = 1'b0;  wr_cycle[19423] = 1'b0;  addr_rom[19423]='h00000000;  wr_data_rom[19423]='h00000000;
    rd_cycle[19424] = 1'b0;  wr_cycle[19424] = 1'b0;  addr_rom[19424]='h00000000;  wr_data_rom[19424]='h00000000;
    rd_cycle[19425] = 1'b0;  wr_cycle[19425] = 1'b0;  addr_rom[19425]='h00000000;  wr_data_rom[19425]='h00000000;
    rd_cycle[19426] = 1'b0;  wr_cycle[19426] = 1'b0;  addr_rom[19426]='h00000000;  wr_data_rom[19426]='h00000000;
    rd_cycle[19427] = 1'b0;  wr_cycle[19427] = 1'b0;  addr_rom[19427]='h00000000;  wr_data_rom[19427]='h00000000;
    rd_cycle[19428] = 1'b0;  wr_cycle[19428] = 1'b0;  addr_rom[19428]='h00000000;  wr_data_rom[19428]='h00000000;
    rd_cycle[19429] = 1'b0;  wr_cycle[19429] = 1'b0;  addr_rom[19429]='h00000000;  wr_data_rom[19429]='h00000000;
    rd_cycle[19430] = 1'b0;  wr_cycle[19430] = 1'b0;  addr_rom[19430]='h00000000;  wr_data_rom[19430]='h00000000;
    rd_cycle[19431] = 1'b0;  wr_cycle[19431] = 1'b0;  addr_rom[19431]='h00000000;  wr_data_rom[19431]='h00000000;
    rd_cycle[19432] = 1'b0;  wr_cycle[19432] = 1'b0;  addr_rom[19432]='h00000000;  wr_data_rom[19432]='h00000000;
    rd_cycle[19433] = 1'b0;  wr_cycle[19433] = 1'b0;  addr_rom[19433]='h00000000;  wr_data_rom[19433]='h00000000;
    rd_cycle[19434] = 1'b0;  wr_cycle[19434] = 1'b0;  addr_rom[19434]='h00000000;  wr_data_rom[19434]='h00000000;
    rd_cycle[19435] = 1'b0;  wr_cycle[19435] = 1'b0;  addr_rom[19435]='h00000000;  wr_data_rom[19435]='h00000000;
    rd_cycle[19436] = 1'b0;  wr_cycle[19436] = 1'b0;  addr_rom[19436]='h00000000;  wr_data_rom[19436]='h00000000;
    rd_cycle[19437] = 1'b0;  wr_cycle[19437] = 1'b0;  addr_rom[19437]='h00000000;  wr_data_rom[19437]='h00000000;
    rd_cycle[19438] = 1'b0;  wr_cycle[19438] = 1'b0;  addr_rom[19438]='h00000000;  wr_data_rom[19438]='h00000000;
    rd_cycle[19439] = 1'b0;  wr_cycle[19439] = 1'b0;  addr_rom[19439]='h00000000;  wr_data_rom[19439]='h00000000;
    rd_cycle[19440] = 1'b0;  wr_cycle[19440] = 1'b0;  addr_rom[19440]='h00000000;  wr_data_rom[19440]='h00000000;
    rd_cycle[19441] = 1'b0;  wr_cycle[19441] = 1'b0;  addr_rom[19441]='h00000000;  wr_data_rom[19441]='h00000000;
    rd_cycle[19442] = 1'b0;  wr_cycle[19442] = 1'b0;  addr_rom[19442]='h00000000;  wr_data_rom[19442]='h00000000;
    rd_cycle[19443] = 1'b0;  wr_cycle[19443] = 1'b0;  addr_rom[19443]='h00000000;  wr_data_rom[19443]='h00000000;
    rd_cycle[19444] = 1'b0;  wr_cycle[19444] = 1'b0;  addr_rom[19444]='h00000000;  wr_data_rom[19444]='h00000000;
    rd_cycle[19445] = 1'b0;  wr_cycle[19445] = 1'b0;  addr_rom[19445]='h00000000;  wr_data_rom[19445]='h00000000;
    rd_cycle[19446] = 1'b0;  wr_cycle[19446] = 1'b0;  addr_rom[19446]='h00000000;  wr_data_rom[19446]='h00000000;
    rd_cycle[19447] = 1'b0;  wr_cycle[19447] = 1'b0;  addr_rom[19447]='h00000000;  wr_data_rom[19447]='h00000000;
    rd_cycle[19448] = 1'b0;  wr_cycle[19448] = 1'b0;  addr_rom[19448]='h00000000;  wr_data_rom[19448]='h00000000;
    rd_cycle[19449] = 1'b0;  wr_cycle[19449] = 1'b0;  addr_rom[19449]='h00000000;  wr_data_rom[19449]='h00000000;
    rd_cycle[19450] = 1'b0;  wr_cycle[19450] = 1'b0;  addr_rom[19450]='h00000000;  wr_data_rom[19450]='h00000000;
    rd_cycle[19451] = 1'b0;  wr_cycle[19451] = 1'b0;  addr_rom[19451]='h00000000;  wr_data_rom[19451]='h00000000;
    rd_cycle[19452] = 1'b0;  wr_cycle[19452] = 1'b0;  addr_rom[19452]='h00000000;  wr_data_rom[19452]='h00000000;
    rd_cycle[19453] = 1'b0;  wr_cycle[19453] = 1'b0;  addr_rom[19453]='h00000000;  wr_data_rom[19453]='h00000000;
    rd_cycle[19454] = 1'b0;  wr_cycle[19454] = 1'b0;  addr_rom[19454]='h00000000;  wr_data_rom[19454]='h00000000;
    rd_cycle[19455] = 1'b0;  wr_cycle[19455] = 1'b0;  addr_rom[19455]='h00000000;  wr_data_rom[19455]='h00000000;
    rd_cycle[19456] = 1'b0;  wr_cycle[19456] = 1'b0;  addr_rom[19456]='h00000000;  wr_data_rom[19456]='h00000000;
    rd_cycle[19457] = 1'b0;  wr_cycle[19457] = 1'b0;  addr_rom[19457]='h00000000;  wr_data_rom[19457]='h00000000;
    rd_cycle[19458] = 1'b0;  wr_cycle[19458] = 1'b0;  addr_rom[19458]='h00000000;  wr_data_rom[19458]='h00000000;
    rd_cycle[19459] = 1'b0;  wr_cycle[19459] = 1'b0;  addr_rom[19459]='h00000000;  wr_data_rom[19459]='h00000000;
    rd_cycle[19460] = 1'b0;  wr_cycle[19460] = 1'b0;  addr_rom[19460]='h00000000;  wr_data_rom[19460]='h00000000;
    rd_cycle[19461] = 1'b0;  wr_cycle[19461] = 1'b0;  addr_rom[19461]='h00000000;  wr_data_rom[19461]='h00000000;
    rd_cycle[19462] = 1'b0;  wr_cycle[19462] = 1'b0;  addr_rom[19462]='h00000000;  wr_data_rom[19462]='h00000000;
    rd_cycle[19463] = 1'b0;  wr_cycle[19463] = 1'b0;  addr_rom[19463]='h00000000;  wr_data_rom[19463]='h00000000;
    rd_cycle[19464] = 1'b0;  wr_cycle[19464] = 1'b0;  addr_rom[19464]='h00000000;  wr_data_rom[19464]='h00000000;
    rd_cycle[19465] = 1'b0;  wr_cycle[19465] = 1'b0;  addr_rom[19465]='h00000000;  wr_data_rom[19465]='h00000000;
    rd_cycle[19466] = 1'b0;  wr_cycle[19466] = 1'b0;  addr_rom[19466]='h00000000;  wr_data_rom[19466]='h00000000;
    rd_cycle[19467] = 1'b0;  wr_cycle[19467] = 1'b0;  addr_rom[19467]='h00000000;  wr_data_rom[19467]='h00000000;
    rd_cycle[19468] = 1'b0;  wr_cycle[19468] = 1'b0;  addr_rom[19468]='h00000000;  wr_data_rom[19468]='h00000000;
    rd_cycle[19469] = 1'b0;  wr_cycle[19469] = 1'b0;  addr_rom[19469]='h00000000;  wr_data_rom[19469]='h00000000;
    rd_cycle[19470] = 1'b0;  wr_cycle[19470] = 1'b0;  addr_rom[19470]='h00000000;  wr_data_rom[19470]='h00000000;
    rd_cycle[19471] = 1'b0;  wr_cycle[19471] = 1'b0;  addr_rom[19471]='h00000000;  wr_data_rom[19471]='h00000000;
    rd_cycle[19472] = 1'b0;  wr_cycle[19472] = 1'b0;  addr_rom[19472]='h00000000;  wr_data_rom[19472]='h00000000;
    rd_cycle[19473] = 1'b0;  wr_cycle[19473] = 1'b0;  addr_rom[19473]='h00000000;  wr_data_rom[19473]='h00000000;
    rd_cycle[19474] = 1'b0;  wr_cycle[19474] = 1'b0;  addr_rom[19474]='h00000000;  wr_data_rom[19474]='h00000000;
    rd_cycle[19475] = 1'b0;  wr_cycle[19475] = 1'b0;  addr_rom[19475]='h00000000;  wr_data_rom[19475]='h00000000;
    rd_cycle[19476] = 1'b0;  wr_cycle[19476] = 1'b0;  addr_rom[19476]='h00000000;  wr_data_rom[19476]='h00000000;
    rd_cycle[19477] = 1'b0;  wr_cycle[19477] = 1'b0;  addr_rom[19477]='h00000000;  wr_data_rom[19477]='h00000000;
    rd_cycle[19478] = 1'b0;  wr_cycle[19478] = 1'b0;  addr_rom[19478]='h00000000;  wr_data_rom[19478]='h00000000;
    rd_cycle[19479] = 1'b0;  wr_cycle[19479] = 1'b0;  addr_rom[19479]='h00000000;  wr_data_rom[19479]='h00000000;
    rd_cycle[19480] = 1'b0;  wr_cycle[19480] = 1'b0;  addr_rom[19480]='h00000000;  wr_data_rom[19480]='h00000000;
    rd_cycle[19481] = 1'b0;  wr_cycle[19481] = 1'b0;  addr_rom[19481]='h00000000;  wr_data_rom[19481]='h00000000;
    rd_cycle[19482] = 1'b0;  wr_cycle[19482] = 1'b0;  addr_rom[19482]='h00000000;  wr_data_rom[19482]='h00000000;
    rd_cycle[19483] = 1'b0;  wr_cycle[19483] = 1'b0;  addr_rom[19483]='h00000000;  wr_data_rom[19483]='h00000000;
    rd_cycle[19484] = 1'b0;  wr_cycle[19484] = 1'b0;  addr_rom[19484]='h00000000;  wr_data_rom[19484]='h00000000;
    rd_cycle[19485] = 1'b0;  wr_cycle[19485] = 1'b0;  addr_rom[19485]='h00000000;  wr_data_rom[19485]='h00000000;
    rd_cycle[19486] = 1'b0;  wr_cycle[19486] = 1'b0;  addr_rom[19486]='h00000000;  wr_data_rom[19486]='h00000000;
    rd_cycle[19487] = 1'b0;  wr_cycle[19487] = 1'b0;  addr_rom[19487]='h00000000;  wr_data_rom[19487]='h00000000;
    rd_cycle[19488] = 1'b0;  wr_cycle[19488] = 1'b0;  addr_rom[19488]='h00000000;  wr_data_rom[19488]='h00000000;
    rd_cycle[19489] = 1'b0;  wr_cycle[19489] = 1'b0;  addr_rom[19489]='h00000000;  wr_data_rom[19489]='h00000000;
    rd_cycle[19490] = 1'b0;  wr_cycle[19490] = 1'b0;  addr_rom[19490]='h00000000;  wr_data_rom[19490]='h00000000;
    rd_cycle[19491] = 1'b0;  wr_cycle[19491] = 1'b0;  addr_rom[19491]='h00000000;  wr_data_rom[19491]='h00000000;
    rd_cycle[19492] = 1'b0;  wr_cycle[19492] = 1'b0;  addr_rom[19492]='h00000000;  wr_data_rom[19492]='h00000000;
    rd_cycle[19493] = 1'b0;  wr_cycle[19493] = 1'b0;  addr_rom[19493]='h00000000;  wr_data_rom[19493]='h00000000;
    rd_cycle[19494] = 1'b0;  wr_cycle[19494] = 1'b0;  addr_rom[19494]='h00000000;  wr_data_rom[19494]='h00000000;
    rd_cycle[19495] = 1'b0;  wr_cycle[19495] = 1'b0;  addr_rom[19495]='h00000000;  wr_data_rom[19495]='h00000000;
    rd_cycle[19496] = 1'b0;  wr_cycle[19496] = 1'b0;  addr_rom[19496]='h00000000;  wr_data_rom[19496]='h00000000;
    rd_cycle[19497] = 1'b0;  wr_cycle[19497] = 1'b0;  addr_rom[19497]='h00000000;  wr_data_rom[19497]='h00000000;
    rd_cycle[19498] = 1'b0;  wr_cycle[19498] = 1'b0;  addr_rom[19498]='h00000000;  wr_data_rom[19498]='h00000000;
    rd_cycle[19499] = 1'b0;  wr_cycle[19499] = 1'b0;  addr_rom[19499]='h00000000;  wr_data_rom[19499]='h00000000;
    rd_cycle[19500] = 1'b0;  wr_cycle[19500] = 1'b0;  addr_rom[19500]='h00000000;  wr_data_rom[19500]='h00000000;
    rd_cycle[19501] = 1'b0;  wr_cycle[19501] = 1'b0;  addr_rom[19501]='h00000000;  wr_data_rom[19501]='h00000000;
    rd_cycle[19502] = 1'b0;  wr_cycle[19502] = 1'b0;  addr_rom[19502]='h00000000;  wr_data_rom[19502]='h00000000;
    rd_cycle[19503] = 1'b0;  wr_cycle[19503] = 1'b0;  addr_rom[19503]='h00000000;  wr_data_rom[19503]='h00000000;
    rd_cycle[19504] = 1'b0;  wr_cycle[19504] = 1'b0;  addr_rom[19504]='h00000000;  wr_data_rom[19504]='h00000000;
    rd_cycle[19505] = 1'b0;  wr_cycle[19505] = 1'b0;  addr_rom[19505]='h00000000;  wr_data_rom[19505]='h00000000;
    rd_cycle[19506] = 1'b0;  wr_cycle[19506] = 1'b0;  addr_rom[19506]='h00000000;  wr_data_rom[19506]='h00000000;
    rd_cycle[19507] = 1'b0;  wr_cycle[19507] = 1'b0;  addr_rom[19507]='h00000000;  wr_data_rom[19507]='h00000000;
    rd_cycle[19508] = 1'b0;  wr_cycle[19508] = 1'b0;  addr_rom[19508]='h00000000;  wr_data_rom[19508]='h00000000;
    rd_cycle[19509] = 1'b0;  wr_cycle[19509] = 1'b0;  addr_rom[19509]='h00000000;  wr_data_rom[19509]='h00000000;
    rd_cycle[19510] = 1'b0;  wr_cycle[19510] = 1'b0;  addr_rom[19510]='h00000000;  wr_data_rom[19510]='h00000000;
    rd_cycle[19511] = 1'b0;  wr_cycle[19511] = 1'b0;  addr_rom[19511]='h00000000;  wr_data_rom[19511]='h00000000;
    rd_cycle[19512] = 1'b0;  wr_cycle[19512] = 1'b0;  addr_rom[19512]='h00000000;  wr_data_rom[19512]='h00000000;
    rd_cycle[19513] = 1'b0;  wr_cycle[19513] = 1'b0;  addr_rom[19513]='h00000000;  wr_data_rom[19513]='h00000000;
    rd_cycle[19514] = 1'b0;  wr_cycle[19514] = 1'b0;  addr_rom[19514]='h00000000;  wr_data_rom[19514]='h00000000;
    rd_cycle[19515] = 1'b0;  wr_cycle[19515] = 1'b0;  addr_rom[19515]='h00000000;  wr_data_rom[19515]='h00000000;
    rd_cycle[19516] = 1'b0;  wr_cycle[19516] = 1'b0;  addr_rom[19516]='h00000000;  wr_data_rom[19516]='h00000000;
    rd_cycle[19517] = 1'b0;  wr_cycle[19517] = 1'b0;  addr_rom[19517]='h00000000;  wr_data_rom[19517]='h00000000;
    rd_cycle[19518] = 1'b0;  wr_cycle[19518] = 1'b0;  addr_rom[19518]='h00000000;  wr_data_rom[19518]='h00000000;
    rd_cycle[19519] = 1'b0;  wr_cycle[19519] = 1'b0;  addr_rom[19519]='h00000000;  wr_data_rom[19519]='h00000000;
    rd_cycle[19520] = 1'b0;  wr_cycle[19520] = 1'b0;  addr_rom[19520]='h00000000;  wr_data_rom[19520]='h00000000;
    rd_cycle[19521] = 1'b0;  wr_cycle[19521] = 1'b0;  addr_rom[19521]='h00000000;  wr_data_rom[19521]='h00000000;
    rd_cycle[19522] = 1'b0;  wr_cycle[19522] = 1'b0;  addr_rom[19522]='h00000000;  wr_data_rom[19522]='h00000000;
    rd_cycle[19523] = 1'b0;  wr_cycle[19523] = 1'b0;  addr_rom[19523]='h00000000;  wr_data_rom[19523]='h00000000;
    rd_cycle[19524] = 1'b0;  wr_cycle[19524] = 1'b0;  addr_rom[19524]='h00000000;  wr_data_rom[19524]='h00000000;
    rd_cycle[19525] = 1'b0;  wr_cycle[19525] = 1'b0;  addr_rom[19525]='h00000000;  wr_data_rom[19525]='h00000000;
    rd_cycle[19526] = 1'b0;  wr_cycle[19526] = 1'b0;  addr_rom[19526]='h00000000;  wr_data_rom[19526]='h00000000;
    rd_cycle[19527] = 1'b0;  wr_cycle[19527] = 1'b0;  addr_rom[19527]='h00000000;  wr_data_rom[19527]='h00000000;
    rd_cycle[19528] = 1'b0;  wr_cycle[19528] = 1'b0;  addr_rom[19528]='h00000000;  wr_data_rom[19528]='h00000000;
    rd_cycle[19529] = 1'b0;  wr_cycle[19529] = 1'b0;  addr_rom[19529]='h00000000;  wr_data_rom[19529]='h00000000;
    rd_cycle[19530] = 1'b0;  wr_cycle[19530] = 1'b0;  addr_rom[19530]='h00000000;  wr_data_rom[19530]='h00000000;
    rd_cycle[19531] = 1'b0;  wr_cycle[19531] = 1'b0;  addr_rom[19531]='h00000000;  wr_data_rom[19531]='h00000000;
    rd_cycle[19532] = 1'b0;  wr_cycle[19532] = 1'b0;  addr_rom[19532]='h00000000;  wr_data_rom[19532]='h00000000;
    rd_cycle[19533] = 1'b0;  wr_cycle[19533] = 1'b0;  addr_rom[19533]='h00000000;  wr_data_rom[19533]='h00000000;
    rd_cycle[19534] = 1'b0;  wr_cycle[19534] = 1'b0;  addr_rom[19534]='h00000000;  wr_data_rom[19534]='h00000000;
    rd_cycle[19535] = 1'b0;  wr_cycle[19535] = 1'b0;  addr_rom[19535]='h00000000;  wr_data_rom[19535]='h00000000;
    rd_cycle[19536] = 1'b0;  wr_cycle[19536] = 1'b0;  addr_rom[19536]='h00000000;  wr_data_rom[19536]='h00000000;
    rd_cycle[19537] = 1'b0;  wr_cycle[19537] = 1'b0;  addr_rom[19537]='h00000000;  wr_data_rom[19537]='h00000000;
    rd_cycle[19538] = 1'b0;  wr_cycle[19538] = 1'b0;  addr_rom[19538]='h00000000;  wr_data_rom[19538]='h00000000;
    rd_cycle[19539] = 1'b0;  wr_cycle[19539] = 1'b0;  addr_rom[19539]='h00000000;  wr_data_rom[19539]='h00000000;
    rd_cycle[19540] = 1'b0;  wr_cycle[19540] = 1'b0;  addr_rom[19540]='h00000000;  wr_data_rom[19540]='h00000000;
    rd_cycle[19541] = 1'b0;  wr_cycle[19541] = 1'b0;  addr_rom[19541]='h00000000;  wr_data_rom[19541]='h00000000;
    rd_cycle[19542] = 1'b0;  wr_cycle[19542] = 1'b0;  addr_rom[19542]='h00000000;  wr_data_rom[19542]='h00000000;
    rd_cycle[19543] = 1'b0;  wr_cycle[19543] = 1'b0;  addr_rom[19543]='h00000000;  wr_data_rom[19543]='h00000000;
    rd_cycle[19544] = 1'b0;  wr_cycle[19544] = 1'b0;  addr_rom[19544]='h00000000;  wr_data_rom[19544]='h00000000;
    rd_cycle[19545] = 1'b0;  wr_cycle[19545] = 1'b0;  addr_rom[19545]='h00000000;  wr_data_rom[19545]='h00000000;
    rd_cycle[19546] = 1'b0;  wr_cycle[19546] = 1'b0;  addr_rom[19546]='h00000000;  wr_data_rom[19546]='h00000000;
    rd_cycle[19547] = 1'b0;  wr_cycle[19547] = 1'b0;  addr_rom[19547]='h00000000;  wr_data_rom[19547]='h00000000;
    rd_cycle[19548] = 1'b0;  wr_cycle[19548] = 1'b0;  addr_rom[19548]='h00000000;  wr_data_rom[19548]='h00000000;
    rd_cycle[19549] = 1'b0;  wr_cycle[19549] = 1'b0;  addr_rom[19549]='h00000000;  wr_data_rom[19549]='h00000000;
    rd_cycle[19550] = 1'b0;  wr_cycle[19550] = 1'b0;  addr_rom[19550]='h00000000;  wr_data_rom[19550]='h00000000;
    rd_cycle[19551] = 1'b0;  wr_cycle[19551] = 1'b0;  addr_rom[19551]='h00000000;  wr_data_rom[19551]='h00000000;
    rd_cycle[19552] = 1'b0;  wr_cycle[19552] = 1'b0;  addr_rom[19552]='h00000000;  wr_data_rom[19552]='h00000000;
    rd_cycle[19553] = 1'b0;  wr_cycle[19553] = 1'b0;  addr_rom[19553]='h00000000;  wr_data_rom[19553]='h00000000;
    rd_cycle[19554] = 1'b0;  wr_cycle[19554] = 1'b0;  addr_rom[19554]='h00000000;  wr_data_rom[19554]='h00000000;
    rd_cycle[19555] = 1'b0;  wr_cycle[19555] = 1'b0;  addr_rom[19555]='h00000000;  wr_data_rom[19555]='h00000000;
    rd_cycle[19556] = 1'b0;  wr_cycle[19556] = 1'b0;  addr_rom[19556]='h00000000;  wr_data_rom[19556]='h00000000;
    rd_cycle[19557] = 1'b0;  wr_cycle[19557] = 1'b0;  addr_rom[19557]='h00000000;  wr_data_rom[19557]='h00000000;
    rd_cycle[19558] = 1'b0;  wr_cycle[19558] = 1'b0;  addr_rom[19558]='h00000000;  wr_data_rom[19558]='h00000000;
    rd_cycle[19559] = 1'b0;  wr_cycle[19559] = 1'b0;  addr_rom[19559]='h00000000;  wr_data_rom[19559]='h00000000;
    rd_cycle[19560] = 1'b0;  wr_cycle[19560] = 1'b0;  addr_rom[19560]='h00000000;  wr_data_rom[19560]='h00000000;
    rd_cycle[19561] = 1'b0;  wr_cycle[19561] = 1'b0;  addr_rom[19561]='h00000000;  wr_data_rom[19561]='h00000000;
    rd_cycle[19562] = 1'b0;  wr_cycle[19562] = 1'b0;  addr_rom[19562]='h00000000;  wr_data_rom[19562]='h00000000;
    rd_cycle[19563] = 1'b0;  wr_cycle[19563] = 1'b0;  addr_rom[19563]='h00000000;  wr_data_rom[19563]='h00000000;
    rd_cycle[19564] = 1'b0;  wr_cycle[19564] = 1'b0;  addr_rom[19564]='h00000000;  wr_data_rom[19564]='h00000000;
    rd_cycle[19565] = 1'b0;  wr_cycle[19565] = 1'b0;  addr_rom[19565]='h00000000;  wr_data_rom[19565]='h00000000;
    rd_cycle[19566] = 1'b0;  wr_cycle[19566] = 1'b0;  addr_rom[19566]='h00000000;  wr_data_rom[19566]='h00000000;
    rd_cycle[19567] = 1'b0;  wr_cycle[19567] = 1'b0;  addr_rom[19567]='h00000000;  wr_data_rom[19567]='h00000000;
    rd_cycle[19568] = 1'b0;  wr_cycle[19568] = 1'b0;  addr_rom[19568]='h00000000;  wr_data_rom[19568]='h00000000;
    rd_cycle[19569] = 1'b0;  wr_cycle[19569] = 1'b0;  addr_rom[19569]='h00000000;  wr_data_rom[19569]='h00000000;
    rd_cycle[19570] = 1'b0;  wr_cycle[19570] = 1'b0;  addr_rom[19570]='h00000000;  wr_data_rom[19570]='h00000000;
    rd_cycle[19571] = 1'b0;  wr_cycle[19571] = 1'b0;  addr_rom[19571]='h00000000;  wr_data_rom[19571]='h00000000;
    rd_cycle[19572] = 1'b0;  wr_cycle[19572] = 1'b0;  addr_rom[19572]='h00000000;  wr_data_rom[19572]='h00000000;
    rd_cycle[19573] = 1'b0;  wr_cycle[19573] = 1'b0;  addr_rom[19573]='h00000000;  wr_data_rom[19573]='h00000000;
    rd_cycle[19574] = 1'b0;  wr_cycle[19574] = 1'b0;  addr_rom[19574]='h00000000;  wr_data_rom[19574]='h00000000;
    rd_cycle[19575] = 1'b0;  wr_cycle[19575] = 1'b0;  addr_rom[19575]='h00000000;  wr_data_rom[19575]='h00000000;
    rd_cycle[19576] = 1'b0;  wr_cycle[19576] = 1'b0;  addr_rom[19576]='h00000000;  wr_data_rom[19576]='h00000000;
    rd_cycle[19577] = 1'b0;  wr_cycle[19577] = 1'b0;  addr_rom[19577]='h00000000;  wr_data_rom[19577]='h00000000;
    rd_cycle[19578] = 1'b0;  wr_cycle[19578] = 1'b0;  addr_rom[19578]='h00000000;  wr_data_rom[19578]='h00000000;
    rd_cycle[19579] = 1'b0;  wr_cycle[19579] = 1'b0;  addr_rom[19579]='h00000000;  wr_data_rom[19579]='h00000000;
    rd_cycle[19580] = 1'b0;  wr_cycle[19580] = 1'b0;  addr_rom[19580]='h00000000;  wr_data_rom[19580]='h00000000;
    rd_cycle[19581] = 1'b0;  wr_cycle[19581] = 1'b0;  addr_rom[19581]='h00000000;  wr_data_rom[19581]='h00000000;
    rd_cycle[19582] = 1'b0;  wr_cycle[19582] = 1'b0;  addr_rom[19582]='h00000000;  wr_data_rom[19582]='h00000000;
    rd_cycle[19583] = 1'b0;  wr_cycle[19583] = 1'b0;  addr_rom[19583]='h00000000;  wr_data_rom[19583]='h00000000;
    rd_cycle[19584] = 1'b0;  wr_cycle[19584] = 1'b0;  addr_rom[19584]='h00000000;  wr_data_rom[19584]='h00000000;
    rd_cycle[19585] = 1'b0;  wr_cycle[19585] = 1'b0;  addr_rom[19585]='h00000000;  wr_data_rom[19585]='h00000000;
    rd_cycle[19586] = 1'b0;  wr_cycle[19586] = 1'b0;  addr_rom[19586]='h00000000;  wr_data_rom[19586]='h00000000;
    rd_cycle[19587] = 1'b0;  wr_cycle[19587] = 1'b0;  addr_rom[19587]='h00000000;  wr_data_rom[19587]='h00000000;
    rd_cycle[19588] = 1'b0;  wr_cycle[19588] = 1'b0;  addr_rom[19588]='h00000000;  wr_data_rom[19588]='h00000000;
    rd_cycle[19589] = 1'b0;  wr_cycle[19589] = 1'b0;  addr_rom[19589]='h00000000;  wr_data_rom[19589]='h00000000;
    rd_cycle[19590] = 1'b0;  wr_cycle[19590] = 1'b0;  addr_rom[19590]='h00000000;  wr_data_rom[19590]='h00000000;
    rd_cycle[19591] = 1'b0;  wr_cycle[19591] = 1'b0;  addr_rom[19591]='h00000000;  wr_data_rom[19591]='h00000000;
    rd_cycle[19592] = 1'b0;  wr_cycle[19592] = 1'b0;  addr_rom[19592]='h00000000;  wr_data_rom[19592]='h00000000;
    rd_cycle[19593] = 1'b0;  wr_cycle[19593] = 1'b0;  addr_rom[19593]='h00000000;  wr_data_rom[19593]='h00000000;
    rd_cycle[19594] = 1'b0;  wr_cycle[19594] = 1'b0;  addr_rom[19594]='h00000000;  wr_data_rom[19594]='h00000000;
    rd_cycle[19595] = 1'b0;  wr_cycle[19595] = 1'b0;  addr_rom[19595]='h00000000;  wr_data_rom[19595]='h00000000;
    rd_cycle[19596] = 1'b0;  wr_cycle[19596] = 1'b0;  addr_rom[19596]='h00000000;  wr_data_rom[19596]='h00000000;
    rd_cycle[19597] = 1'b0;  wr_cycle[19597] = 1'b0;  addr_rom[19597]='h00000000;  wr_data_rom[19597]='h00000000;
    rd_cycle[19598] = 1'b0;  wr_cycle[19598] = 1'b0;  addr_rom[19598]='h00000000;  wr_data_rom[19598]='h00000000;
    rd_cycle[19599] = 1'b0;  wr_cycle[19599] = 1'b0;  addr_rom[19599]='h00000000;  wr_data_rom[19599]='h00000000;
    rd_cycle[19600] = 1'b0;  wr_cycle[19600] = 1'b0;  addr_rom[19600]='h00000000;  wr_data_rom[19600]='h00000000;
    rd_cycle[19601] = 1'b0;  wr_cycle[19601] = 1'b0;  addr_rom[19601]='h00000000;  wr_data_rom[19601]='h00000000;
    rd_cycle[19602] = 1'b0;  wr_cycle[19602] = 1'b0;  addr_rom[19602]='h00000000;  wr_data_rom[19602]='h00000000;
    rd_cycle[19603] = 1'b0;  wr_cycle[19603] = 1'b0;  addr_rom[19603]='h00000000;  wr_data_rom[19603]='h00000000;
    rd_cycle[19604] = 1'b0;  wr_cycle[19604] = 1'b0;  addr_rom[19604]='h00000000;  wr_data_rom[19604]='h00000000;
    rd_cycle[19605] = 1'b0;  wr_cycle[19605] = 1'b0;  addr_rom[19605]='h00000000;  wr_data_rom[19605]='h00000000;
    rd_cycle[19606] = 1'b0;  wr_cycle[19606] = 1'b0;  addr_rom[19606]='h00000000;  wr_data_rom[19606]='h00000000;
    rd_cycle[19607] = 1'b0;  wr_cycle[19607] = 1'b0;  addr_rom[19607]='h00000000;  wr_data_rom[19607]='h00000000;
    rd_cycle[19608] = 1'b0;  wr_cycle[19608] = 1'b0;  addr_rom[19608]='h00000000;  wr_data_rom[19608]='h00000000;
    rd_cycle[19609] = 1'b0;  wr_cycle[19609] = 1'b0;  addr_rom[19609]='h00000000;  wr_data_rom[19609]='h00000000;
    rd_cycle[19610] = 1'b0;  wr_cycle[19610] = 1'b0;  addr_rom[19610]='h00000000;  wr_data_rom[19610]='h00000000;
    rd_cycle[19611] = 1'b0;  wr_cycle[19611] = 1'b0;  addr_rom[19611]='h00000000;  wr_data_rom[19611]='h00000000;
    rd_cycle[19612] = 1'b0;  wr_cycle[19612] = 1'b0;  addr_rom[19612]='h00000000;  wr_data_rom[19612]='h00000000;
    rd_cycle[19613] = 1'b0;  wr_cycle[19613] = 1'b0;  addr_rom[19613]='h00000000;  wr_data_rom[19613]='h00000000;
    rd_cycle[19614] = 1'b0;  wr_cycle[19614] = 1'b0;  addr_rom[19614]='h00000000;  wr_data_rom[19614]='h00000000;
    rd_cycle[19615] = 1'b0;  wr_cycle[19615] = 1'b0;  addr_rom[19615]='h00000000;  wr_data_rom[19615]='h00000000;
    rd_cycle[19616] = 1'b0;  wr_cycle[19616] = 1'b0;  addr_rom[19616]='h00000000;  wr_data_rom[19616]='h00000000;
    rd_cycle[19617] = 1'b0;  wr_cycle[19617] = 1'b0;  addr_rom[19617]='h00000000;  wr_data_rom[19617]='h00000000;
    rd_cycle[19618] = 1'b0;  wr_cycle[19618] = 1'b0;  addr_rom[19618]='h00000000;  wr_data_rom[19618]='h00000000;
    rd_cycle[19619] = 1'b0;  wr_cycle[19619] = 1'b0;  addr_rom[19619]='h00000000;  wr_data_rom[19619]='h00000000;
    rd_cycle[19620] = 1'b0;  wr_cycle[19620] = 1'b0;  addr_rom[19620]='h00000000;  wr_data_rom[19620]='h00000000;
    rd_cycle[19621] = 1'b0;  wr_cycle[19621] = 1'b0;  addr_rom[19621]='h00000000;  wr_data_rom[19621]='h00000000;
    rd_cycle[19622] = 1'b0;  wr_cycle[19622] = 1'b0;  addr_rom[19622]='h00000000;  wr_data_rom[19622]='h00000000;
    rd_cycle[19623] = 1'b0;  wr_cycle[19623] = 1'b0;  addr_rom[19623]='h00000000;  wr_data_rom[19623]='h00000000;
    rd_cycle[19624] = 1'b0;  wr_cycle[19624] = 1'b0;  addr_rom[19624]='h00000000;  wr_data_rom[19624]='h00000000;
    rd_cycle[19625] = 1'b0;  wr_cycle[19625] = 1'b0;  addr_rom[19625]='h00000000;  wr_data_rom[19625]='h00000000;
    rd_cycle[19626] = 1'b0;  wr_cycle[19626] = 1'b0;  addr_rom[19626]='h00000000;  wr_data_rom[19626]='h00000000;
    rd_cycle[19627] = 1'b0;  wr_cycle[19627] = 1'b0;  addr_rom[19627]='h00000000;  wr_data_rom[19627]='h00000000;
    rd_cycle[19628] = 1'b0;  wr_cycle[19628] = 1'b0;  addr_rom[19628]='h00000000;  wr_data_rom[19628]='h00000000;
    rd_cycle[19629] = 1'b0;  wr_cycle[19629] = 1'b0;  addr_rom[19629]='h00000000;  wr_data_rom[19629]='h00000000;
    rd_cycle[19630] = 1'b0;  wr_cycle[19630] = 1'b0;  addr_rom[19630]='h00000000;  wr_data_rom[19630]='h00000000;
    rd_cycle[19631] = 1'b0;  wr_cycle[19631] = 1'b0;  addr_rom[19631]='h00000000;  wr_data_rom[19631]='h00000000;
    rd_cycle[19632] = 1'b0;  wr_cycle[19632] = 1'b0;  addr_rom[19632]='h00000000;  wr_data_rom[19632]='h00000000;
    rd_cycle[19633] = 1'b0;  wr_cycle[19633] = 1'b0;  addr_rom[19633]='h00000000;  wr_data_rom[19633]='h00000000;
    rd_cycle[19634] = 1'b0;  wr_cycle[19634] = 1'b0;  addr_rom[19634]='h00000000;  wr_data_rom[19634]='h00000000;
    rd_cycle[19635] = 1'b0;  wr_cycle[19635] = 1'b0;  addr_rom[19635]='h00000000;  wr_data_rom[19635]='h00000000;
    rd_cycle[19636] = 1'b0;  wr_cycle[19636] = 1'b0;  addr_rom[19636]='h00000000;  wr_data_rom[19636]='h00000000;
    rd_cycle[19637] = 1'b0;  wr_cycle[19637] = 1'b0;  addr_rom[19637]='h00000000;  wr_data_rom[19637]='h00000000;
    rd_cycle[19638] = 1'b0;  wr_cycle[19638] = 1'b0;  addr_rom[19638]='h00000000;  wr_data_rom[19638]='h00000000;
    rd_cycle[19639] = 1'b0;  wr_cycle[19639] = 1'b0;  addr_rom[19639]='h00000000;  wr_data_rom[19639]='h00000000;
    rd_cycle[19640] = 1'b0;  wr_cycle[19640] = 1'b0;  addr_rom[19640]='h00000000;  wr_data_rom[19640]='h00000000;
    rd_cycle[19641] = 1'b0;  wr_cycle[19641] = 1'b0;  addr_rom[19641]='h00000000;  wr_data_rom[19641]='h00000000;
    rd_cycle[19642] = 1'b0;  wr_cycle[19642] = 1'b0;  addr_rom[19642]='h00000000;  wr_data_rom[19642]='h00000000;
    rd_cycle[19643] = 1'b0;  wr_cycle[19643] = 1'b0;  addr_rom[19643]='h00000000;  wr_data_rom[19643]='h00000000;
    rd_cycle[19644] = 1'b0;  wr_cycle[19644] = 1'b0;  addr_rom[19644]='h00000000;  wr_data_rom[19644]='h00000000;
    rd_cycle[19645] = 1'b0;  wr_cycle[19645] = 1'b0;  addr_rom[19645]='h00000000;  wr_data_rom[19645]='h00000000;
    rd_cycle[19646] = 1'b0;  wr_cycle[19646] = 1'b0;  addr_rom[19646]='h00000000;  wr_data_rom[19646]='h00000000;
    rd_cycle[19647] = 1'b0;  wr_cycle[19647] = 1'b0;  addr_rom[19647]='h00000000;  wr_data_rom[19647]='h00000000;
    rd_cycle[19648] = 1'b0;  wr_cycle[19648] = 1'b0;  addr_rom[19648]='h00000000;  wr_data_rom[19648]='h00000000;
    rd_cycle[19649] = 1'b0;  wr_cycle[19649] = 1'b0;  addr_rom[19649]='h00000000;  wr_data_rom[19649]='h00000000;
    rd_cycle[19650] = 1'b0;  wr_cycle[19650] = 1'b0;  addr_rom[19650]='h00000000;  wr_data_rom[19650]='h00000000;
    rd_cycle[19651] = 1'b0;  wr_cycle[19651] = 1'b0;  addr_rom[19651]='h00000000;  wr_data_rom[19651]='h00000000;
    rd_cycle[19652] = 1'b0;  wr_cycle[19652] = 1'b0;  addr_rom[19652]='h00000000;  wr_data_rom[19652]='h00000000;
    rd_cycle[19653] = 1'b0;  wr_cycle[19653] = 1'b0;  addr_rom[19653]='h00000000;  wr_data_rom[19653]='h00000000;
    rd_cycle[19654] = 1'b0;  wr_cycle[19654] = 1'b0;  addr_rom[19654]='h00000000;  wr_data_rom[19654]='h00000000;
    rd_cycle[19655] = 1'b0;  wr_cycle[19655] = 1'b0;  addr_rom[19655]='h00000000;  wr_data_rom[19655]='h00000000;
    rd_cycle[19656] = 1'b0;  wr_cycle[19656] = 1'b0;  addr_rom[19656]='h00000000;  wr_data_rom[19656]='h00000000;
    rd_cycle[19657] = 1'b0;  wr_cycle[19657] = 1'b0;  addr_rom[19657]='h00000000;  wr_data_rom[19657]='h00000000;
    rd_cycle[19658] = 1'b0;  wr_cycle[19658] = 1'b0;  addr_rom[19658]='h00000000;  wr_data_rom[19658]='h00000000;
    rd_cycle[19659] = 1'b0;  wr_cycle[19659] = 1'b0;  addr_rom[19659]='h00000000;  wr_data_rom[19659]='h00000000;
    rd_cycle[19660] = 1'b0;  wr_cycle[19660] = 1'b0;  addr_rom[19660]='h00000000;  wr_data_rom[19660]='h00000000;
    rd_cycle[19661] = 1'b0;  wr_cycle[19661] = 1'b0;  addr_rom[19661]='h00000000;  wr_data_rom[19661]='h00000000;
    rd_cycle[19662] = 1'b0;  wr_cycle[19662] = 1'b0;  addr_rom[19662]='h00000000;  wr_data_rom[19662]='h00000000;
    rd_cycle[19663] = 1'b0;  wr_cycle[19663] = 1'b0;  addr_rom[19663]='h00000000;  wr_data_rom[19663]='h00000000;
    rd_cycle[19664] = 1'b0;  wr_cycle[19664] = 1'b0;  addr_rom[19664]='h00000000;  wr_data_rom[19664]='h00000000;
    rd_cycle[19665] = 1'b0;  wr_cycle[19665] = 1'b0;  addr_rom[19665]='h00000000;  wr_data_rom[19665]='h00000000;
    rd_cycle[19666] = 1'b0;  wr_cycle[19666] = 1'b0;  addr_rom[19666]='h00000000;  wr_data_rom[19666]='h00000000;
    rd_cycle[19667] = 1'b0;  wr_cycle[19667] = 1'b0;  addr_rom[19667]='h00000000;  wr_data_rom[19667]='h00000000;
    rd_cycle[19668] = 1'b0;  wr_cycle[19668] = 1'b0;  addr_rom[19668]='h00000000;  wr_data_rom[19668]='h00000000;
    rd_cycle[19669] = 1'b0;  wr_cycle[19669] = 1'b0;  addr_rom[19669]='h00000000;  wr_data_rom[19669]='h00000000;
    rd_cycle[19670] = 1'b0;  wr_cycle[19670] = 1'b0;  addr_rom[19670]='h00000000;  wr_data_rom[19670]='h00000000;
    rd_cycle[19671] = 1'b0;  wr_cycle[19671] = 1'b0;  addr_rom[19671]='h00000000;  wr_data_rom[19671]='h00000000;
    rd_cycle[19672] = 1'b0;  wr_cycle[19672] = 1'b0;  addr_rom[19672]='h00000000;  wr_data_rom[19672]='h00000000;
    rd_cycle[19673] = 1'b0;  wr_cycle[19673] = 1'b0;  addr_rom[19673]='h00000000;  wr_data_rom[19673]='h00000000;
    rd_cycle[19674] = 1'b0;  wr_cycle[19674] = 1'b0;  addr_rom[19674]='h00000000;  wr_data_rom[19674]='h00000000;
    rd_cycle[19675] = 1'b0;  wr_cycle[19675] = 1'b0;  addr_rom[19675]='h00000000;  wr_data_rom[19675]='h00000000;
    rd_cycle[19676] = 1'b0;  wr_cycle[19676] = 1'b0;  addr_rom[19676]='h00000000;  wr_data_rom[19676]='h00000000;
    rd_cycle[19677] = 1'b0;  wr_cycle[19677] = 1'b0;  addr_rom[19677]='h00000000;  wr_data_rom[19677]='h00000000;
    rd_cycle[19678] = 1'b0;  wr_cycle[19678] = 1'b0;  addr_rom[19678]='h00000000;  wr_data_rom[19678]='h00000000;
    rd_cycle[19679] = 1'b0;  wr_cycle[19679] = 1'b0;  addr_rom[19679]='h00000000;  wr_data_rom[19679]='h00000000;
    rd_cycle[19680] = 1'b0;  wr_cycle[19680] = 1'b0;  addr_rom[19680]='h00000000;  wr_data_rom[19680]='h00000000;
    rd_cycle[19681] = 1'b0;  wr_cycle[19681] = 1'b0;  addr_rom[19681]='h00000000;  wr_data_rom[19681]='h00000000;
    rd_cycle[19682] = 1'b0;  wr_cycle[19682] = 1'b0;  addr_rom[19682]='h00000000;  wr_data_rom[19682]='h00000000;
    rd_cycle[19683] = 1'b0;  wr_cycle[19683] = 1'b0;  addr_rom[19683]='h00000000;  wr_data_rom[19683]='h00000000;
    rd_cycle[19684] = 1'b0;  wr_cycle[19684] = 1'b0;  addr_rom[19684]='h00000000;  wr_data_rom[19684]='h00000000;
    rd_cycle[19685] = 1'b0;  wr_cycle[19685] = 1'b0;  addr_rom[19685]='h00000000;  wr_data_rom[19685]='h00000000;
    rd_cycle[19686] = 1'b0;  wr_cycle[19686] = 1'b0;  addr_rom[19686]='h00000000;  wr_data_rom[19686]='h00000000;
    rd_cycle[19687] = 1'b0;  wr_cycle[19687] = 1'b0;  addr_rom[19687]='h00000000;  wr_data_rom[19687]='h00000000;
    rd_cycle[19688] = 1'b0;  wr_cycle[19688] = 1'b0;  addr_rom[19688]='h00000000;  wr_data_rom[19688]='h00000000;
    rd_cycle[19689] = 1'b0;  wr_cycle[19689] = 1'b0;  addr_rom[19689]='h00000000;  wr_data_rom[19689]='h00000000;
    rd_cycle[19690] = 1'b0;  wr_cycle[19690] = 1'b0;  addr_rom[19690]='h00000000;  wr_data_rom[19690]='h00000000;
    rd_cycle[19691] = 1'b0;  wr_cycle[19691] = 1'b0;  addr_rom[19691]='h00000000;  wr_data_rom[19691]='h00000000;
    rd_cycle[19692] = 1'b0;  wr_cycle[19692] = 1'b0;  addr_rom[19692]='h00000000;  wr_data_rom[19692]='h00000000;
    rd_cycle[19693] = 1'b0;  wr_cycle[19693] = 1'b0;  addr_rom[19693]='h00000000;  wr_data_rom[19693]='h00000000;
    rd_cycle[19694] = 1'b0;  wr_cycle[19694] = 1'b0;  addr_rom[19694]='h00000000;  wr_data_rom[19694]='h00000000;
    rd_cycle[19695] = 1'b0;  wr_cycle[19695] = 1'b0;  addr_rom[19695]='h00000000;  wr_data_rom[19695]='h00000000;
    rd_cycle[19696] = 1'b0;  wr_cycle[19696] = 1'b0;  addr_rom[19696]='h00000000;  wr_data_rom[19696]='h00000000;
    rd_cycle[19697] = 1'b0;  wr_cycle[19697] = 1'b0;  addr_rom[19697]='h00000000;  wr_data_rom[19697]='h00000000;
    rd_cycle[19698] = 1'b0;  wr_cycle[19698] = 1'b0;  addr_rom[19698]='h00000000;  wr_data_rom[19698]='h00000000;
    rd_cycle[19699] = 1'b0;  wr_cycle[19699] = 1'b0;  addr_rom[19699]='h00000000;  wr_data_rom[19699]='h00000000;
    rd_cycle[19700] = 1'b0;  wr_cycle[19700] = 1'b0;  addr_rom[19700]='h00000000;  wr_data_rom[19700]='h00000000;
    rd_cycle[19701] = 1'b0;  wr_cycle[19701] = 1'b0;  addr_rom[19701]='h00000000;  wr_data_rom[19701]='h00000000;
    rd_cycle[19702] = 1'b0;  wr_cycle[19702] = 1'b0;  addr_rom[19702]='h00000000;  wr_data_rom[19702]='h00000000;
    rd_cycle[19703] = 1'b0;  wr_cycle[19703] = 1'b0;  addr_rom[19703]='h00000000;  wr_data_rom[19703]='h00000000;
    rd_cycle[19704] = 1'b0;  wr_cycle[19704] = 1'b0;  addr_rom[19704]='h00000000;  wr_data_rom[19704]='h00000000;
    rd_cycle[19705] = 1'b0;  wr_cycle[19705] = 1'b0;  addr_rom[19705]='h00000000;  wr_data_rom[19705]='h00000000;
    rd_cycle[19706] = 1'b0;  wr_cycle[19706] = 1'b0;  addr_rom[19706]='h00000000;  wr_data_rom[19706]='h00000000;
    rd_cycle[19707] = 1'b0;  wr_cycle[19707] = 1'b0;  addr_rom[19707]='h00000000;  wr_data_rom[19707]='h00000000;
    rd_cycle[19708] = 1'b0;  wr_cycle[19708] = 1'b0;  addr_rom[19708]='h00000000;  wr_data_rom[19708]='h00000000;
    rd_cycle[19709] = 1'b0;  wr_cycle[19709] = 1'b0;  addr_rom[19709]='h00000000;  wr_data_rom[19709]='h00000000;
    rd_cycle[19710] = 1'b0;  wr_cycle[19710] = 1'b0;  addr_rom[19710]='h00000000;  wr_data_rom[19710]='h00000000;
    rd_cycle[19711] = 1'b0;  wr_cycle[19711] = 1'b0;  addr_rom[19711]='h00000000;  wr_data_rom[19711]='h00000000;
    rd_cycle[19712] = 1'b0;  wr_cycle[19712] = 1'b0;  addr_rom[19712]='h00000000;  wr_data_rom[19712]='h00000000;
    rd_cycle[19713] = 1'b0;  wr_cycle[19713] = 1'b0;  addr_rom[19713]='h00000000;  wr_data_rom[19713]='h00000000;
    rd_cycle[19714] = 1'b0;  wr_cycle[19714] = 1'b0;  addr_rom[19714]='h00000000;  wr_data_rom[19714]='h00000000;
    rd_cycle[19715] = 1'b0;  wr_cycle[19715] = 1'b0;  addr_rom[19715]='h00000000;  wr_data_rom[19715]='h00000000;
    rd_cycle[19716] = 1'b0;  wr_cycle[19716] = 1'b0;  addr_rom[19716]='h00000000;  wr_data_rom[19716]='h00000000;
    rd_cycle[19717] = 1'b0;  wr_cycle[19717] = 1'b0;  addr_rom[19717]='h00000000;  wr_data_rom[19717]='h00000000;
    rd_cycle[19718] = 1'b0;  wr_cycle[19718] = 1'b0;  addr_rom[19718]='h00000000;  wr_data_rom[19718]='h00000000;
    rd_cycle[19719] = 1'b0;  wr_cycle[19719] = 1'b0;  addr_rom[19719]='h00000000;  wr_data_rom[19719]='h00000000;
    rd_cycle[19720] = 1'b0;  wr_cycle[19720] = 1'b0;  addr_rom[19720]='h00000000;  wr_data_rom[19720]='h00000000;
    rd_cycle[19721] = 1'b0;  wr_cycle[19721] = 1'b0;  addr_rom[19721]='h00000000;  wr_data_rom[19721]='h00000000;
    rd_cycle[19722] = 1'b0;  wr_cycle[19722] = 1'b0;  addr_rom[19722]='h00000000;  wr_data_rom[19722]='h00000000;
    rd_cycle[19723] = 1'b0;  wr_cycle[19723] = 1'b0;  addr_rom[19723]='h00000000;  wr_data_rom[19723]='h00000000;
    rd_cycle[19724] = 1'b0;  wr_cycle[19724] = 1'b0;  addr_rom[19724]='h00000000;  wr_data_rom[19724]='h00000000;
    rd_cycle[19725] = 1'b0;  wr_cycle[19725] = 1'b0;  addr_rom[19725]='h00000000;  wr_data_rom[19725]='h00000000;
    rd_cycle[19726] = 1'b0;  wr_cycle[19726] = 1'b0;  addr_rom[19726]='h00000000;  wr_data_rom[19726]='h00000000;
    rd_cycle[19727] = 1'b0;  wr_cycle[19727] = 1'b0;  addr_rom[19727]='h00000000;  wr_data_rom[19727]='h00000000;
    rd_cycle[19728] = 1'b0;  wr_cycle[19728] = 1'b0;  addr_rom[19728]='h00000000;  wr_data_rom[19728]='h00000000;
    rd_cycle[19729] = 1'b0;  wr_cycle[19729] = 1'b0;  addr_rom[19729]='h00000000;  wr_data_rom[19729]='h00000000;
    rd_cycle[19730] = 1'b0;  wr_cycle[19730] = 1'b0;  addr_rom[19730]='h00000000;  wr_data_rom[19730]='h00000000;
    rd_cycle[19731] = 1'b0;  wr_cycle[19731] = 1'b0;  addr_rom[19731]='h00000000;  wr_data_rom[19731]='h00000000;
    rd_cycle[19732] = 1'b0;  wr_cycle[19732] = 1'b0;  addr_rom[19732]='h00000000;  wr_data_rom[19732]='h00000000;
    rd_cycle[19733] = 1'b0;  wr_cycle[19733] = 1'b0;  addr_rom[19733]='h00000000;  wr_data_rom[19733]='h00000000;
    rd_cycle[19734] = 1'b0;  wr_cycle[19734] = 1'b0;  addr_rom[19734]='h00000000;  wr_data_rom[19734]='h00000000;
    rd_cycle[19735] = 1'b0;  wr_cycle[19735] = 1'b0;  addr_rom[19735]='h00000000;  wr_data_rom[19735]='h00000000;
    rd_cycle[19736] = 1'b0;  wr_cycle[19736] = 1'b0;  addr_rom[19736]='h00000000;  wr_data_rom[19736]='h00000000;
    rd_cycle[19737] = 1'b0;  wr_cycle[19737] = 1'b0;  addr_rom[19737]='h00000000;  wr_data_rom[19737]='h00000000;
    rd_cycle[19738] = 1'b0;  wr_cycle[19738] = 1'b0;  addr_rom[19738]='h00000000;  wr_data_rom[19738]='h00000000;
    rd_cycle[19739] = 1'b0;  wr_cycle[19739] = 1'b0;  addr_rom[19739]='h00000000;  wr_data_rom[19739]='h00000000;
    rd_cycle[19740] = 1'b0;  wr_cycle[19740] = 1'b0;  addr_rom[19740]='h00000000;  wr_data_rom[19740]='h00000000;
    rd_cycle[19741] = 1'b0;  wr_cycle[19741] = 1'b0;  addr_rom[19741]='h00000000;  wr_data_rom[19741]='h00000000;
    rd_cycle[19742] = 1'b0;  wr_cycle[19742] = 1'b0;  addr_rom[19742]='h00000000;  wr_data_rom[19742]='h00000000;
    rd_cycle[19743] = 1'b0;  wr_cycle[19743] = 1'b0;  addr_rom[19743]='h00000000;  wr_data_rom[19743]='h00000000;
    rd_cycle[19744] = 1'b0;  wr_cycle[19744] = 1'b0;  addr_rom[19744]='h00000000;  wr_data_rom[19744]='h00000000;
    rd_cycle[19745] = 1'b0;  wr_cycle[19745] = 1'b0;  addr_rom[19745]='h00000000;  wr_data_rom[19745]='h00000000;
    rd_cycle[19746] = 1'b0;  wr_cycle[19746] = 1'b0;  addr_rom[19746]='h00000000;  wr_data_rom[19746]='h00000000;
    rd_cycle[19747] = 1'b0;  wr_cycle[19747] = 1'b0;  addr_rom[19747]='h00000000;  wr_data_rom[19747]='h00000000;
    rd_cycle[19748] = 1'b0;  wr_cycle[19748] = 1'b0;  addr_rom[19748]='h00000000;  wr_data_rom[19748]='h00000000;
    rd_cycle[19749] = 1'b0;  wr_cycle[19749] = 1'b0;  addr_rom[19749]='h00000000;  wr_data_rom[19749]='h00000000;
    rd_cycle[19750] = 1'b0;  wr_cycle[19750] = 1'b0;  addr_rom[19750]='h00000000;  wr_data_rom[19750]='h00000000;
    rd_cycle[19751] = 1'b0;  wr_cycle[19751] = 1'b0;  addr_rom[19751]='h00000000;  wr_data_rom[19751]='h00000000;
    rd_cycle[19752] = 1'b0;  wr_cycle[19752] = 1'b0;  addr_rom[19752]='h00000000;  wr_data_rom[19752]='h00000000;
    rd_cycle[19753] = 1'b0;  wr_cycle[19753] = 1'b0;  addr_rom[19753]='h00000000;  wr_data_rom[19753]='h00000000;
    rd_cycle[19754] = 1'b0;  wr_cycle[19754] = 1'b0;  addr_rom[19754]='h00000000;  wr_data_rom[19754]='h00000000;
    rd_cycle[19755] = 1'b0;  wr_cycle[19755] = 1'b0;  addr_rom[19755]='h00000000;  wr_data_rom[19755]='h00000000;
    rd_cycle[19756] = 1'b0;  wr_cycle[19756] = 1'b0;  addr_rom[19756]='h00000000;  wr_data_rom[19756]='h00000000;
    rd_cycle[19757] = 1'b0;  wr_cycle[19757] = 1'b0;  addr_rom[19757]='h00000000;  wr_data_rom[19757]='h00000000;
    rd_cycle[19758] = 1'b0;  wr_cycle[19758] = 1'b0;  addr_rom[19758]='h00000000;  wr_data_rom[19758]='h00000000;
    rd_cycle[19759] = 1'b0;  wr_cycle[19759] = 1'b0;  addr_rom[19759]='h00000000;  wr_data_rom[19759]='h00000000;
    rd_cycle[19760] = 1'b0;  wr_cycle[19760] = 1'b0;  addr_rom[19760]='h00000000;  wr_data_rom[19760]='h00000000;
    rd_cycle[19761] = 1'b0;  wr_cycle[19761] = 1'b0;  addr_rom[19761]='h00000000;  wr_data_rom[19761]='h00000000;
    rd_cycle[19762] = 1'b0;  wr_cycle[19762] = 1'b0;  addr_rom[19762]='h00000000;  wr_data_rom[19762]='h00000000;
    rd_cycle[19763] = 1'b0;  wr_cycle[19763] = 1'b0;  addr_rom[19763]='h00000000;  wr_data_rom[19763]='h00000000;
    rd_cycle[19764] = 1'b0;  wr_cycle[19764] = 1'b0;  addr_rom[19764]='h00000000;  wr_data_rom[19764]='h00000000;
    rd_cycle[19765] = 1'b0;  wr_cycle[19765] = 1'b0;  addr_rom[19765]='h00000000;  wr_data_rom[19765]='h00000000;
    rd_cycle[19766] = 1'b0;  wr_cycle[19766] = 1'b0;  addr_rom[19766]='h00000000;  wr_data_rom[19766]='h00000000;
    rd_cycle[19767] = 1'b0;  wr_cycle[19767] = 1'b0;  addr_rom[19767]='h00000000;  wr_data_rom[19767]='h00000000;
    rd_cycle[19768] = 1'b0;  wr_cycle[19768] = 1'b0;  addr_rom[19768]='h00000000;  wr_data_rom[19768]='h00000000;
    rd_cycle[19769] = 1'b0;  wr_cycle[19769] = 1'b0;  addr_rom[19769]='h00000000;  wr_data_rom[19769]='h00000000;
    rd_cycle[19770] = 1'b0;  wr_cycle[19770] = 1'b0;  addr_rom[19770]='h00000000;  wr_data_rom[19770]='h00000000;
    rd_cycle[19771] = 1'b0;  wr_cycle[19771] = 1'b0;  addr_rom[19771]='h00000000;  wr_data_rom[19771]='h00000000;
    rd_cycle[19772] = 1'b0;  wr_cycle[19772] = 1'b0;  addr_rom[19772]='h00000000;  wr_data_rom[19772]='h00000000;
    rd_cycle[19773] = 1'b0;  wr_cycle[19773] = 1'b0;  addr_rom[19773]='h00000000;  wr_data_rom[19773]='h00000000;
    rd_cycle[19774] = 1'b0;  wr_cycle[19774] = 1'b0;  addr_rom[19774]='h00000000;  wr_data_rom[19774]='h00000000;
    rd_cycle[19775] = 1'b0;  wr_cycle[19775] = 1'b0;  addr_rom[19775]='h00000000;  wr_data_rom[19775]='h00000000;
    rd_cycle[19776] = 1'b0;  wr_cycle[19776] = 1'b0;  addr_rom[19776]='h00000000;  wr_data_rom[19776]='h00000000;
    rd_cycle[19777] = 1'b0;  wr_cycle[19777] = 1'b0;  addr_rom[19777]='h00000000;  wr_data_rom[19777]='h00000000;
    rd_cycle[19778] = 1'b0;  wr_cycle[19778] = 1'b0;  addr_rom[19778]='h00000000;  wr_data_rom[19778]='h00000000;
    rd_cycle[19779] = 1'b0;  wr_cycle[19779] = 1'b0;  addr_rom[19779]='h00000000;  wr_data_rom[19779]='h00000000;
    rd_cycle[19780] = 1'b0;  wr_cycle[19780] = 1'b0;  addr_rom[19780]='h00000000;  wr_data_rom[19780]='h00000000;
    rd_cycle[19781] = 1'b0;  wr_cycle[19781] = 1'b0;  addr_rom[19781]='h00000000;  wr_data_rom[19781]='h00000000;
    rd_cycle[19782] = 1'b0;  wr_cycle[19782] = 1'b0;  addr_rom[19782]='h00000000;  wr_data_rom[19782]='h00000000;
    rd_cycle[19783] = 1'b0;  wr_cycle[19783] = 1'b0;  addr_rom[19783]='h00000000;  wr_data_rom[19783]='h00000000;
    rd_cycle[19784] = 1'b0;  wr_cycle[19784] = 1'b0;  addr_rom[19784]='h00000000;  wr_data_rom[19784]='h00000000;
    rd_cycle[19785] = 1'b0;  wr_cycle[19785] = 1'b0;  addr_rom[19785]='h00000000;  wr_data_rom[19785]='h00000000;
    rd_cycle[19786] = 1'b0;  wr_cycle[19786] = 1'b0;  addr_rom[19786]='h00000000;  wr_data_rom[19786]='h00000000;
    rd_cycle[19787] = 1'b0;  wr_cycle[19787] = 1'b0;  addr_rom[19787]='h00000000;  wr_data_rom[19787]='h00000000;
    rd_cycle[19788] = 1'b0;  wr_cycle[19788] = 1'b0;  addr_rom[19788]='h00000000;  wr_data_rom[19788]='h00000000;
    rd_cycle[19789] = 1'b0;  wr_cycle[19789] = 1'b0;  addr_rom[19789]='h00000000;  wr_data_rom[19789]='h00000000;
    rd_cycle[19790] = 1'b0;  wr_cycle[19790] = 1'b0;  addr_rom[19790]='h00000000;  wr_data_rom[19790]='h00000000;
    rd_cycle[19791] = 1'b0;  wr_cycle[19791] = 1'b0;  addr_rom[19791]='h00000000;  wr_data_rom[19791]='h00000000;
    rd_cycle[19792] = 1'b0;  wr_cycle[19792] = 1'b0;  addr_rom[19792]='h00000000;  wr_data_rom[19792]='h00000000;
    rd_cycle[19793] = 1'b0;  wr_cycle[19793] = 1'b0;  addr_rom[19793]='h00000000;  wr_data_rom[19793]='h00000000;
    rd_cycle[19794] = 1'b0;  wr_cycle[19794] = 1'b0;  addr_rom[19794]='h00000000;  wr_data_rom[19794]='h00000000;
    rd_cycle[19795] = 1'b0;  wr_cycle[19795] = 1'b0;  addr_rom[19795]='h00000000;  wr_data_rom[19795]='h00000000;
    rd_cycle[19796] = 1'b0;  wr_cycle[19796] = 1'b0;  addr_rom[19796]='h00000000;  wr_data_rom[19796]='h00000000;
    rd_cycle[19797] = 1'b0;  wr_cycle[19797] = 1'b0;  addr_rom[19797]='h00000000;  wr_data_rom[19797]='h00000000;
    rd_cycle[19798] = 1'b0;  wr_cycle[19798] = 1'b0;  addr_rom[19798]='h00000000;  wr_data_rom[19798]='h00000000;
    rd_cycle[19799] = 1'b0;  wr_cycle[19799] = 1'b0;  addr_rom[19799]='h00000000;  wr_data_rom[19799]='h00000000;
    rd_cycle[19800] = 1'b0;  wr_cycle[19800] = 1'b0;  addr_rom[19800]='h00000000;  wr_data_rom[19800]='h00000000;
    rd_cycle[19801] = 1'b0;  wr_cycle[19801] = 1'b0;  addr_rom[19801]='h00000000;  wr_data_rom[19801]='h00000000;
    rd_cycle[19802] = 1'b0;  wr_cycle[19802] = 1'b0;  addr_rom[19802]='h00000000;  wr_data_rom[19802]='h00000000;
    rd_cycle[19803] = 1'b0;  wr_cycle[19803] = 1'b0;  addr_rom[19803]='h00000000;  wr_data_rom[19803]='h00000000;
    rd_cycle[19804] = 1'b0;  wr_cycle[19804] = 1'b0;  addr_rom[19804]='h00000000;  wr_data_rom[19804]='h00000000;
    rd_cycle[19805] = 1'b0;  wr_cycle[19805] = 1'b0;  addr_rom[19805]='h00000000;  wr_data_rom[19805]='h00000000;
    rd_cycle[19806] = 1'b0;  wr_cycle[19806] = 1'b0;  addr_rom[19806]='h00000000;  wr_data_rom[19806]='h00000000;
    rd_cycle[19807] = 1'b0;  wr_cycle[19807] = 1'b0;  addr_rom[19807]='h00000000;  wr_data_rom[19807]='h00000000;
    rd_cycle[19808] = 1'b0;  wr_cycle[19808] = 1'b0;  addr_rom[19808]='h00000000;  wr_data_rom[19808]='h00000000;
    rd_cycle[19809] = 1'b0;  wr_cycle[19809] = 1'b0;  addr_rom[19809]='h00000000;  wr_data_rom[19809]='h00000000;
    rd_cycle[19810] = 1'b0;  wr_cycle[19810] = 1'b0;  addr_rom[19810]='h00000000;  wr_data_rom[19810]='h00000000;
    rd_cycle[19811] = 1'b0;  wr_cycle[19811] = 1'b0;  addr_rom[19811]='h00000000;  wr_data_rom[19811]='h00000000;
    rd_cycle[19812] = 1'b0;  wr_cycle[19812] = 1'b0;  addr_rom[19812]='h00000000;  wr_data_rom[19812]='h00000000;
    rd_cycle[19813] = 1'b0;  wr_cycle[19813] = 1'b0;  addr_rom[19813]='h00000000;  wr_data_rom[19813]='h00000000;
    rd_cycle[19814] = 1'b0;  wr_cycle[19814] = 1'b0;  addr_rom[19814]='h00000000;  wr_data_rom[19814]='h00000000;
    rd_cycle[19815] = 1'b0;  wr_cycle[19815] = 1'b0;  addr_rom[19815]='h00000000;  wr_data_rom[19815]='h00000000;
    rd_cycle[19816] = 1'b0;  wr_cycle[19816] = 1'b0;  addr_rom[19816]='h00000000;  wr_data_rom[19816]='h00000000;
    rd_cycle[19817] = 1'b0;  wr_cycle[19817] = 1'b0;  addr_rom[19817]='h00000000;  wr_data_rom[19817]='h00000000;
    rd_cycle[19818] = 1'b0;  wr_cycle[19818] = 1'b0;  addr_rom[19818]='h00000000;  wr_data_rom[19818]='h00000000;
    rd_cycle[19819] = 1'b0;  wr_cycle[19819] = 1'b0;  addr_rom[19819]='h00000000;  wr_data_rom[19819]='h00000000;
    rd_cycle[19820] = 1'b0;  wr_cycle[19820] = 1'b0;  addr_rom[19820]='h00000000;  wr_data_rom[19820]='h00000000;
    rd_cycle[19821] = 1'b0;  wr_cycle[19821] = 1'b0;  addr_rom[19821]='h00000000;  wr_data_rom[19821]='h00000000;
    rd_cycle[19822] = 1'b0;  wr_cycle[19822] = 1'b0;  addr_rom[19822]='h00000000;  wr_data_rom[19822]='h00000000;
    rd_cycle[19823] = 1'b0;  wr_cycle[19823] = 1'b0;  addr_rom[19823]='h00000000;  wr_data_rom[19823]='h00000000;
    rd_cycle[19824] = 1'b0;  wr_cycle[19824] = 1'b0;  addr_rom[19824]='h00000000;  wr_data_rom[19824]='h00000000;
    rd_cycle[19825] = 1'b0;  wr_cycle[19825] = 1'b0;  addr_rom[19825]='h00000000;  wr_data_rom[19825]='h00000000;
    rd_cycle[19826] = 1'b0;  wr_cycle[19826] = 1'b0;  addr_rom[19826]='h00000000;  wr_data_rom[19826]='h00000000;
    rd_cycle[19827] = 1'b0;  wr_cycle[19827] = 1'b0;  addr_rom[19827]='h00000000;  wr_data_rom[19827]='h00000000;
    rd_cycle[19828] = 1'b0;  wr_cycle[19828] = 1'b0;  addr_rom[19828]='h00000000;  wr_data_rom[19828]='h00000000;
    rd_cycle[19829] = 1'b0;  wr_cycle[19829] = 1'b0;  addr_rom[19829]='h00000000;  wr_data_rom[19829]='h00000000;
    rd_cycle[19830] = 1'b0;  wr_cycle[19830] = 1'b0;  addr_rom[19830]='h00000000;  wr_data_rom[19830]='h00000000;
    rd_cycle[19831] = 1'b0;  wr_cycle[19831] = 1'b0;  addr_rom[19831]='h00000000;  wr_data_rom[19831]='h00000000;
    rd_cycle[19832] = 1'b0;  wr_cycle[19832] = 1'b0;  addr_rom[19832]='h00000000;  wr_data_rom[19832]='h00000000;
    rd_cycle[19833] = 1'b0;  wr_cycle[19833] = 1'b0;  addr_rom[19833]='h00000000;  wr_data_rom[19833]='h00000000;
    rd_cycle[19834] = 1'b0;  wr_cycle[19834] = 1'b0;  addr_rom[19834]='h00000000;  wr_data_rom[19834]='h00000000;
    rd_cycle[19835] = 1'b0;  wr_cycle[19835] = 1'b0;  addr_rom[19835]='h00000000;  wr_data_rom[19835]='h00000000;
    rd_cycle[19836] = 1'b0;  wr_cycle[19836] = 1'b0;  addr_rom[19836]='h00000000;  wr_data_rom[19836]='h00000000;
    rd_cycle[19837] = 1'b0;  wr_cycle[19837] = 1'b0;  addr_rom[19837]='h00000000;  wr_data_rom[19837]='h00000000;
    rd_cycle[19838] = 1'b0;  wr_cycle[19838] = 1'b0;  addr_rom[19838]='h00000000;  wr_data_rom[19838]='h00000000;
    rd_cycle[19839] = 1'b0;  wr_cycle[19839] = 1'b0;  addr_rom[19839]='h00000000;  wr_data_rom[19839]='h00000000;
    rd_cycle[19840] = 1'b0;  wr_cycle[19840] = 1'b0;  addr_rom[19840]='h00000000;  wr_data_rom[19840]='h00000000;
    rd_cycle[19841] = 1'b0;  wr_cycle[19841] = 1'b0;  addr_rom[19841]='h00000000;  wr_data_rom[19841]='h00000000;
    rd_cycle[19842] = 1'b0;  wr_cycle[19842] = 1'b0;  addr_rom[19842]='h00000000;  wr_data_rom[19842]='h00000000;
    rd_cycle[19843] = 1'b0;  wr_cycle[19843] = 1'b0;  addr_rom[19843]='h00000000;  wr_data_rom[19843]='h00000000;
    rd_cycle[19844] = 1'b0;  wr_cycle[19844] = 1'b0;  addr_rom[19844]='h00000000;  wr_data_rom[19844]='h00000000;
    rd_cycle[19845] = 1'b0;  wr_cycle[19845] = 1'b0;  addr_rom[19845]='h00000000;  wr_data_rom[19845]='h00000000;
    rd_cycle[19846] = 1'b0;  wr_cycle[19846] = 1'b0;  addr_rom[19846]='h00000000;  wr_data_rom[19846]='h00000000;
    rd_cycle[19847] = 1'b0;  wr_cycle[19847] = 1'b0;  addr_rom[19847]='h00000000;  wr_data_rom[19847]='h00000000;
    rd_cycle[19848] = 1'b0;  wr_cycle[19848] = 1'b0;  addr_rom[19848]='h00000000;  wr_data_rom[19848]='h00000000;
    rd_cycle[19849] = 1'b0;  wr_cycle[19849] = 1'b0;  addr_rom[19849]='h00000000;  wr_data_rom[19849]='h00000000;
    rd_cycle[19850] = 1'b0;  wr_cycle[19850] = 1'b0;  addr_rom[19850]='h00000000;  wr_data_rom[19850]='h00000000;
    rd_cycle[19851] = 1'b0;  wr_cycle[19851] = 1'b0;  addr_rom[19851]='h00000000;  wr_data_rom[19851]='h00000000;
    rd_cycle[19852] = 1'b0;  wr_cycle[19852] = 1'b0;  addr_rom[19852]='h00000000;  wr_data_rom[19852]='h00000000;
    rd_cycle[19853] = 1'b0;  wr_cycle[19853] = 1'b0;  addr_rom[19853]='h00000000;  wr_data_rom[19853]='h00000000;
    rd_cycle[19854] = 1'b0;  wr_cycle[19854] = 1'b0;  addr_rom[19854]='h00000000;  wr_data_rom[19854]='h00000000;
    rd_cycle[19855] = 1'b0;  wr_cycle[19855] = 1'b0;  addr_rom[19855]='h00000000;  wr_data_rom[19855]='h00000000;
    rd_cycle[19856] = 1'b0;  wr_cycle[19856] = 1'b0;  addr_rom[19856]='h00000000;  wr_data_rom[19856]='h00000000;
    rd_cycle[19857] = 1'b0;  wr_cycle[19857] = 1'b0;  addr_rom[19857]='h00000000;  wr_data_rom[19857]='h00000000;
    rd_cycle[19858] = 1'b0;  wr_cycle[19858] = 1'b0;  addr_rom[19858]='h00000000;  wr_data_rom[19858]='h00000000;
    rd_cycle[19859] = 1'b0;  wr_cycle[19859] = 1'b0;  addr_rom[19859]='h00000000;  wr_data_rom[19859]='h00000000;
    rd_cycle[19860] = 1'b0;  wr_cycle[19860] = 1'b0;  addr_rom[19860]='h00000000;  wr_data_rom[19860]='h00000000;
    rd_cycle[19861] = 1'b0;  wr_cycle[19861] = 1'b0;  addr_rom[19861]='h00000000;  wr_data_rom[19861]='h00000000;
    rd_cycle[19862] = 1'b0;  wr_cycle[19862] = 1'b0;  addr_rom[19862]='h00000000;  wr_data_rom[19862]='h00000000;
    rd_cycle[19863] = 1'b0;  wr_cycle[19863] = 1'b0;  addr_rom[19863]='h00000000;  wr_data_rom[19863]='h00000000;
    rd_cycle[19864] = 1'b0;  wr_cycle[19864] = 1'b0;  addr_rom[19864]='h00000000;  wr_data_rom[19864]='h00000000;
    rd_cycle[19865] = 1'b0;  wr_cycle[19865] = 1'b0;  addr_rom[19865]='h00000000;  wr_data_rom[19865]='h00000000;
    rd_cycle[19866] = 1'b0;  wr_cycle[19866] = 1'b0;  addr_rom[19866]='h00000000;  wr_data_rom[19866]='h00000000;
    rd_cycle[19867] = 1'b0;  wr_cycle[19867] = 1'b0;  addr_rom[19867]='h00000000;  wr_data_rom[19867]='h00000000;
    rd_cycle[19868] = 1'b0;  wr_cycle[19868] = 1'b0;  addr_rom[19868]='h00000000;  wr_data_rom[19868]='h00000000;
    rd_cycle[19869] = 1'b0;  wr_cycle[19869] = 1'b0;  addr_rom[19869]='h00000000;  wr_data_rom[19869]='h00000000;
    rd_cycle[19870] = 1'b0;  wr_cycle[19870] = 1'b0;  addr_rom[19870]='h00000000;  wr_data_rom[19870]='h00000000;
    rd_cycle[19871] = 1'b0;  wr_cycle[19871] = 1'b0;  addr_rom[19871]='h00000000;  wr_data_rom[19871]='h00000000;
    rd_cycle[19872] = 1'b0;  wr_cycle[19872] = 1'b0;  addr_rom[19872]='h00000000;  wr_data_rom[19872]='h00000000;
    rd_cycle[19873] = 1'b0;  wr_cycle[19873] = 1'b0;  addr_rom[19873]='h00000000;  wr_data_rom[19873]='h00000000;
    rd_cycle[19874] = 1'b0;  wr_cycle[19874] = 1'b0;  addr_rom[19874]='h00000000;  wr_data_rom[19874]='h00000000;
    rd_cycle[19875] = 1'b0;  wr_cycle[19875] = 1'b0;  addr_rom[19875]='h00000000;  wr_data_rom[19875]='h00000000;
    rd_cycle[19876] = 1'b0;  wr_cycle[19876] = 1'b0;  addr_rom[19876]='h00000000;  wr_data_rom[19876]='h00000000;
    rd_cycle[19877] = 1'b0;  wr_cycle[19877] = 1'b0;  addr_rom[19877]='h00000000;  wr_data_rom[19877]='h00000000;
    rd_cycle[19878] = 1'b0;  wr_cycle[19878] = 1'b0;  addr_rom[19878]='h00000000;  wr_data_rom[19878]='h00000000;
    rd_cycle[19879] = 1'b0;  wr_cycle[19879] = 1'b0;  addr_rom[19879]='h00000000;  wr_data_rom[19879]='h00000000;
    rd_cycle[19880] = 1'b0;  wr_cycle[19880] = 1'b0;  addr_rom[19880]='h00000000;  wr_data_rom[19880]='h00000000;
    rd_cycle[19881] = 1'b0;  wr_cycle[19881] = 1'b0;  addr_rom[19881]='h00000000;  wr_data_rom[19881]='h00000000;
    rd_cycle[19882] = 1'b0;  wr_cycle[19882] = 1'b0;  addr_rom[19882]='h00000000;  wr_data_rom[19882]='h00000000;
    rd_cycle[19883] = 1'b0;  wr_cycle[19883] = 1'b0;  addr_rom[19883]='h00000000;  wr_data_rom[19883]='h00000000;
    rd_cycle[19884] = 1'b0;  wr_cycle[19884] = 1'b0;  addr_rom[19884]='h00000000;  wr_data_rom[19884]='h00000000;
    rd_cycle[19885] = 1'b0;  wr_cycle[19885] = 1'b0;  addr_rom[19885]='h00000000;  wr_data_rom[19885]='h00000000;
    rd_cycle[19886] = 1'b0;  wr_cycle[19886] = 1'b0;  addr_rom[19886]='h00000000;  wr_data_rom[19886]='h00000000;
    rd_cycle[19887] = 1'b0;  wr_cycle[19887] = 1'b0;  addr_rom[19887]='h00000000;  wr_data_rom[19887]='h00000000;
    rd_cycle[19888] = 1'b0;  wr_cycle[19888] = 1'b0;  addr_rom[19888]='h00000000;  wr_data_rom[19888]='h00000000;
    rd_cycle[19889] = 1'b0;  wr_cycle[19889] = 1'b0;  addr_rom[19889]='h00000000;  wr_data_rom[19889]='h00000000;
    rd_cycle[19890] = 1'b0;  wr_cycle[19890] = 1'b0;  addr_rom[19890]='h00000000;  wr_data_rom[19890]='h00000000;
    rd_cycle[19891] = 1'b0;  wr_cycle[19891] = 1'b0;  addr_rom[19891]='h00000000;  wr_data_rom[19891]='h00000000;
    rd_cycle[19892] = 1'b0;  wr_cycle[19892] = 1'b0;  addr_rom[19892]='h00000000;  wr_data_rom[19892]='h00000000;
    rd_cycle[19893] = 1'b0;  wr_cycle[19893] = 1'b0;  addr_rom[19893]='h00000000;  wr_data_rom[19893]='h00000000;
    rd_cycle[19894] = 1'b0;  wr_cycle[19894] = 1'b0;  addr_rom[19894]='h00000000;  wr_data_rom[19894]='h00000000;
    rd_cycle[19895] = 1'b0;  wr_cycle[19895] = 1'b0;  addr_rom[19895]='h00000000;  wr_data_rom[19895]='h00000000;
    rd_cycle[19896] = 1'b0;  wr_cycle[19896] = 1'b0;  addr_rom[19896]='h00000000;  wr_data_rom[19896]='h00000000;
    rd_cycle[19897] = 1'b0;  wr_cycle[19897] = 1'b0;  addr_rom[19897]='h00000000;  wr_data_rom[19897]='h00000000;
    rd_cycle[19898] = 1'b0;  wr_cycle[19898] = 1'b0;  addr_rom[19898]='h00000000;  wr_data_rom[19898]='h00000000;
    rd_cycle[19899] = 1'b0;  wr_cycle[19899] = 1'b0;  addr_rom[19899]='h00000000;  wr_data_rom[19899]='h00000000;
    rd_cycle[19900] = 1'b0;  wr_cycle[19900] = 1'b0;  addr_rom[19900]='h00000000;  wr_data_rom[19900]='h00000000;
    rd_cycle[19901] = 1'b0;  wr_cycle[19901] = 1'b0;  addr_rom[19901]='h00000000;  wr_data_rom[19901]='h00000000;
    rd_cycle[19902] = 1'b0;  wr_cycle[19902] = 1'b0;  addr_rom[19902]='h00000000;  wr_data_rom[19902]='h00000000;
    rd_cycle[19903] = 1'b0;  wr_cycle[19903] = 1'b0;  addr_rom[19903]='h00000000;  wr_data_rom[19903]='h00000000;
    rd_cycle[19904] = 1'b0;  wr_cycle[19904] = 1'b0;  addr_rom[19904]='h00000000;  wr_data_rom[19904]='h00000000;
    rd_cycle[19905] = 1'b0;  wr_cycle[19905] = 1'b0;  addr_rom[19905]='h00000000;  wr_data_rom[19905]='h00000000;
    rd_cycle[19906] = 1'b0;  wr_cycle[19906] = 1'b0;  addr_rom[19906]='h00000000;  wr_data_rom[19906]='h00000000;
    rd_cycle[19907] = 1'b0;  wr_cycle[19907] = 1'b0;  addr_rom[19907]='h00000000;  wr_data_rom[19907]='h00000000;
    rd_cycle[19908] = 1'b0;  wr_cycle[19908] = 1'b0;  addr_rom[19908]='h00000000;  wr_data_rom[19908]='h00000000;
    rd_cycle[19909] = 1'b0;  wr_cycle[19909] = 1'b0;  addr_rom[19909]='h00000000;  wr_data_rom[19909]='h00000000;
    rd_cycle[19910] = 1'b0;  wr_cycle[19910] = 1'b0;  addr_rom[19910]='h00000000;  wr_data_rom[19910]='h00000000;
    rd_cycle[19911] = 1'b0;  wr_cycle[19911] = 1'b0;  addr_rom[19911]='h00000000;  wr_data_rom[19911]='h00000000;
    rd_cycle[19912] = 1'b0;  wr_cycle[19912] = 1'b0;  addr_rom[19912]='h00000000;  wr_data_rom[19912]='h00000000;
    rd_cycle[19913] = 1'b0;  wr_cycle[19913] = 1'b0;  addr_rom[19913]='h00000000;  wr_data_rom[19913]='h00000000;
    rd_cycle[19914] = 1'b0;  wr_cycle[19914] = 1'b0;  addr_rom[19914]='h00000000;  wr_data_rom[19914]='h00000000;
    rd_cycle[19915] = 1'b0;  wr_cycle[19915] = 1'b0;  addr_rom[19915]='h00000000;  wr_data_rom[19915]='h00000000;
    rd_cycle[19916] = 1'b0;  wr_cycle[19916] = 1'b0;  addr_rom[19916]='h00000000;  wr_data_rom[19916]='h00000000;
    rd_cycle[19917] = 1'b0;  wr_cycle[19917] = 1'b0;  addr_rom[19917]='h00000000;  wr_data_rom[19917]='h00000000;
    rd_cycle[19918] = 1'b0;  wr_cycle[19918] = 1'b0;  addr_rom[19918]='h00000000;  wr_data_rom[19918]='h00000000;
    rd_cycle[19919] = 1'b0;  wr_cycle[19919] = 1'b0;  addr_rom[19919]='h00000000;  wr_data_rom[19919]='h00000000;
    rd_cycle[19920] = 1'b0;  wr_cycle[19920] = 1'b0;  addr_rom[19920]='h00000000;  wr_data_rom[19920]='h00000000;
    rd_cycle[19921] = 1'b0;  wr_cycle[19921] = 1'b0;  addr_rom[19921]='h00000000;  wr_data_rom[19921]='h00000000;
    rd_cycle[19922] = 1'b0;  wr_cycle[19922] = 1'b0;  addr_rom[19922]='h00000000;  wr_data_rom[19922]='h00000000;
    rd_cycle[19923] = 1'b0;  wr_cycle[19923] = 1'b0;  addr_rom[19923]='h00000000;  wr_data_rom[19923]='h00000000;
    rd_cycle[19924] = 1'b0;  wr_cycle[19924] = 1'b0;  addr_rom[19924]='h00000000;  wr_data_rom[19924]='h00000000;
    rd_cycle[19925] = 1'b0;  wr_cycle[19925] = 1'b0;  addr_rom[19925]='h00000000;  wr_data_rom[19925]='h00000000;
    rd_cycle[19926] = 1'b0;  wr_cycle[19926] = 1'b0;  addr_rom[19926]='h00000000;  wr_data_rom[19926]='h00000000;
    rd_cycle[19927] = 1'b0;  wr_cycle[19927] = 1'b0;  addr_rom[19927]='h00000000;  wr_data_rom[19927]='h00000000;
    rd_cycle[19928] = 1'b0;  wr_cycle[19928] = 1'b0;  addr_rom[19928]='h00000000;  wr_data_rom[19928]='h00000000;
    rd_cycle[19929] = 1'b0;  wr_cycle[19929] = 1'b0;  addr_rom[19929]='h00000000;  wr_data_rom[19929]='h00000000;
    rd_cycle[19930] = 1'b0;  wr_cycle[19930] = 1'b0;  addr_rom[19930]='h00000000;  wr_data_rom[19930]='h00000000;
    rd_cycle[19931] = 1'b0;  wr_cycle[19931] = 1'b0;  addr_rom[19931]='h00000000;  wr_data_rom[19931]='h00000000;
    rd_cycle[19932] = 1'b0;  wr_cycle[19932] = 1'b0;  addr_rom[19932]='h00000000;  wr_data_rom[19932]='h00000000;
    rd_cycle[19933] = 1'b0;  wr_cycle[19933] = 1'b0;  addr_rom[19933]='h00000000;  wr_data_rom[19933]='h00000000;
    rd_cycle[19934] = 1'b0;  wr_cycle[19934] = 1'b0;  addr_rom[19934]='h00000000;  wr_data_rom[19934]='h00000000;
    rd_cycle[19935] = 1'b0;  wr_cycle[19935] = 1'b0;  addr_rom[19935]='h00000000;  wr_data_rom[19935]='h00000000;
    rd_cycle[19936] = 1'b0;  wr_cycle[19936] = 1'b0;  addr_rom[19936]='h00000000;  wr_data_rom[19936]='h00000000;
    rd_cycle[19937] = 1'b0;  wr_cycle[19937] = 1'b0;  addr_rom[19937]='h00000000;  wr_data_rom[19937]='h00000000;
    rd_cycle[19938] = 1'b0;  wr_cycle[19938] = 1'b0;  addr_rom[19938]='h00000000;  wr_data_rom[19938]='h00000000;
    rd_cycle[19939] = 1'b0;  wr_cycle[19939] = 1'b0;  addr_rom[19939]='h00000000;  wr_data_rom[19939]='h00000000;
    rd_cycle[19940] = 1'b0;  wr_cycle[19940] = 1'b0;  addr_rom[19940]='h00000000;  wr_data_rom[19940]='h00000000;
    rd_cycle[19941] = 1'b0;  wr_cycle[19941] = 1'b0;  addr_rom[19941]='h00000000;  wr_data_rom[19941]='h00000000;
    rd_cycle[19942] = 1'b0;  wr_cycle[19942] = 1'b0;  addr_rom[19942]='h00000000;  wr_data_rom[19942]='h00000000;
    rd_cycle[19943] = 1'b0;  wr_cycle[19943] = 1'b0;  addr_rom[19943]='h00000000;  wr_data_rom[19943]='h00000000;
    rd_cycle[19944] = 1'b0;  wr_cycle[19944] = 1'b0;  addr_rom[19944]='h00000000;  wr_data_rom[19944]='h00000000;
    rd_cycle[19945] = 1'b0;  wr_cycle[19945] = 1'b0;  addr_rom[19945]='h00000000;  wr_data_rom[19945]='h00000000;
    rd_cycle[19946] = 1'b0;  wr_cycle[19946] = 1'b0;  addr_rom[19946]='h00000000;  wr_data_rom[19946]='h00000000;
    rd_cycle[19947] = 1'b0;  wr_cycle[19947] = 1'b0;  addr_rom[19947]='h00000000;  wr_data_rom[19947]='h00000000;
    rd_cycle[19948] = 1'b0;  wr_cycle[19948] = 1'b0;  addr_rom[19948]='h00000000;  wr_data_rom[19948]='h00000000;
    rd_cycle[19949] = 1'b0;  wr_cycle[19949] = 1'b0;  addr_rom[19949]='h00000000;  wr_data_rom[19949]='h00000000;
    rd_cycle[19950] = 1'b0;  wr_cycle[19950] = 1'b0;  addr_rom[19950]='h00000000;  wr_data_rom[19950]='h00000000;
    rd_cycle[19951] = 1'b0;  wr_cycle[19951] = 1'b0;  addr_rom[19951]='h00000000;  wr_data_rom[19951]='h00000000;
    rd_cycle[19952] = 1'b0;  wr_cycle[19952] = 1'b0;  addr_rom[19952]='h00000000;  wr_data_rom[19952]='h00000000;
    rd_cycle[19953] = 1'b0;  wr_cycle[19953] = 1'b0;  addr_rom[19953]='h00000000;  wr_data_rom[19953]='h00000000;
    rd_cycle[19954] = 1'b0;  wr_cycle[19954] = 1'b0;  addr_rom[19954]='h00000000;  wr_data_rom[19954]='h00000000;
    rd_cycle[19955] = 1'b0;  wr_cycle[19955] = 1'b0;  addr_rom[19955]='h00000000;  wr_data_rom[19955]='h00000000;
    rd_cycle[19956] = 1'b0;  wr_cycle[19956] = 1'b0;  addr_rom[19956]='h00000000;  wr_data_rom[19956]='h00000000;
    rd_cycle[19957] = 1'b0;  wr_cycle[19957] = 1'b0;  addr_rom[19957]='h00000000;  wr_data_rom[19957]='h00000000;
    rd_cycle[19958] = 1'b0;  wr_cycle[19958] = 1'b0;  addr_rom[19958]='h00000000;  wr_data_rom[19958]='h00000000;
    rd_cycle[19959] = 1'b0;  wr_cycle[19959] = 1'b0;  addr_rom[19959]='h00000000;  wr_data_rom[19959]='h00000000;
    rd_cycle[19960] = 1'b0;  wr_cycle[19960] = 1'b0;  addr_rom[19960]='h00000000;  wr_data_rom[19960]='h00000000;
    rd_cycle[19961] = 1'b0;  wr_cycle[19961] = 1'b0;  addr_rom[19961]='h00000000;  wr_data_rom[19961]='h00000000;
    rd_cycle[19962] = 1'b0;  wr_cycle[19962] = 1'b0;  addr_rom[19962]='h00000000;  wr_data_rom[19962]='h00000000;
    rd_cycle[19963] = 1'b0;  wr_cycle[19963] = 1'b0;  addr_rom[19963]='h00000000;  wr_data_rom[19963]='h00000000;
    rd_cycle[19964] = 1'b0;  wr_cycle[19964] = 1'b0;  addr_rom[19964]='h00000000;  wr_data_rom[19964]='h00000000;
    rd_cycle[19965] = 1'b0;  wr_cycle[19965] = 1'b0;  addr_rom[19965]='h00000000;  wr_data_rom[19965]='h00000000;
    rd_cycle[19966] = 1'b0;  wr_cycle[19966] = 1'b0;  addr_rom[19966]='h00000000;  wr_data_rom[19966]='h00000000;
    rd_cycle[19967] = 1'b0;  wr_cycle[19967] = 1'b0;  addr_rom[19967]='h00000000;  wr_data_rom[19967]='h00000000;
    rd_cycle[19968] = 1'b0;  wr_cycle[19968] = 1'b0;  addr_rom[19968]='h00000000;  wr_data_rom[19968]='h00000000;
    rd_cycle[19969] = 1'b0;  wr_cycle[19969] = 1'b0;  addr_rom[19969]='h00000000;  wr_data_rom[19969]='h00000000;
    rd_cycle[19970] = 1'b0;  wr_cycle[19970] = 1'b0;  addr_rom[19970]='h00000000;  wr_data_rom[19970]='h00000000;
    rd_cycle[19971] = 1'b0;  wr_cycle[19971] = 1'b0;  addr_rom[19971]='h00000000;  wr_data_rom[19971]='h00000000;
    rd_cycle[19972] = 1'b0;  wr_cycle[19972] = 1'b0;  addr_rom[19972]='h00000000;  wr_data_rom[19972]='h00000000;
    rd_cycle[19973] = 1'b0;  wr_cycle[19973] = 1'b0;  addr_rom[19973]='h00000000;  wr_data_rom[19973]='h00000000;
    rd_cycle[19974] = 1'b0;  wr_cycle[19974] = 1'b0;  addr_rom[19974]='h00000000;  wr_data_rom[19974]='h00000000;
    rd_cycle[19975] = 1'b0;  wr_cycle[19975] = 1'b0;  addr_rom[19975]='h00000000;  wr_data_rom[19975]='h00000000;
    rd_cycle[19976] = 1'b0;  wr_cycle[19976] = 1'b0;  addr_rom[19976]='h00000000;  wr_data_rom[19976]='h00000000;
    rd_cycle[19977] = 1'b0;  wr_cycle[19977] = 1'b0;  addr_rom[19977]='h00000000;  wr_data_rom[19977]='h00000000;
    rd_cycle[19978] = 1'b0;  wr_cycle[19978] = 1'b0;  addr_rom[19978]='h00000000;  wr_data_rom[19978]='h00000000;
    rd_cycle[19979] = 1'b0;  wr_cycle[19979] = 1'b0;  addr_rom[19979]='h00000000;  wr_data_rom[19979]='h00000000;
    rd_cycle[19980] = 1'b0;  wr_cycle[19980] = 1'b0;  addr_rom[19980]='h00000000;  wr_data_rom[19980]='h00000000;
    rd_cycle[19981] = 1'b0;  wr_cycle[19981] = 1'b0;  addr_rom[19981]='h00000000;  wr_data_rom[19981]='h00000000;
    rd_cycle[19982] = 1'b0;  wr_cycle[19982] = 1'b0;  addr_rom[19982]='h00000000;  wr_data_rom[19982]='h00000000;
    rd_cycle[19983] = 1'b0;  wr_cycle[19983] = 1'b0;  addr_rom[19983]='h00000000;  wr_data_rom[19983]='h00000000;
    rd_cycle[19984] = 1'b0;  wr_cycle[19984] = 1'b0;  addr_rom[19984]='h00000000;  wr_data_rom[19984]='h00000000;
    rd_cycle[19985] = 1'b0;  wr_cycle[19985] = 1'b0;  addr_rom[19985]='h00000000;  wr_data_rom[19985]='h00000000;
    rd_cycle[19986] = 1'b0;  wr_cycle[19986] = 1'b0;  addr_rom[19986]='h00000000;  wr_data_rom[19986]='h00000000;
    rd_cycle[19987] = 1'b0;  wr_cycle[19987] = 1'b0;  addr_rom[19987]='h00000000;  wr_data_rom[19987]='h00000000;
    rd_cycle[19988] = 1'b0;  wr_cycle[19988] = 1'b0;  addr_rom[19988]='h00000000;  wr_data_rom[19988]='h00000000;
    rd_cycle[19989] = 1'b0;  wr_cycle[19989] = 1'b0;  addr_rom[19989]='h00000000;  wr_data_rom[19989]='h00000000;
    rd_cycle[19990] = 1'b0;  wr_cycle[19990] = 1'b0;  addr_rom[19990]='h00000000;  wr_data_rom[19990]='h00000000;
    rd_cycle[19991] = 1'b0;  wr_cycle[19991] = 1'b0;  addr_rom[19991]='h00000000;  wr_data_rom[19991]='h00000000;
    rd_cycle[19992] = 1'b0;  wr_cycle[19992] = 1'b0;  addr_rom[19992]='h00000000;  wr_data_rom[19992]='h00000000;
    rd_cycle[19993] = 1'b0;  wr_cycle[19993] = 1'b0;  addr_rom[19993]='h00000000;  wr_data_rom[19993]='h00000000;
    rd_cycle[19994] = 1'b0;  wr_cycle[19994] = 1'b0;  addr_rom[19994]='h00000000;  wr_data_rom[19994]='h00000000;
    rd_cycle[19995] = 1'b0;  wr_cycle[19995] = 1'b0;  addr_rom[19995]='h00000000;  wr_data_rom[19995]='h00000000;
    rd_cycle[19996] = 1'b0;  wr_cycle[19996] = 1'b0;  addr_rom[19996]='h00000000;  wr_data_rom[19996]='h00000000;
    rd_cycle[19997] = 1'b0;  wr_cycle[19997] = 1'b0;  addr_rom[19997]='h00000000;  wr_data_rom[19997]='h00000000;
    rd_cycle[19998] = 1'b0;  wr_cycle[19998] = 1'b0;  addr_rom[19998]='h00000000;  wr_data_rom[19998]='h00000000;
    rd_cycle[19999] = 1'b0;  wr_cycle[19999] = 1'b0;  addr_rom[19999]='h00000000;  wr_data_rom[19999]='h00000000;
    rd_cycle[20000] = 1'b0;  wr_cycle[20000] = 1'b0;  addr_rom[20000]='h00000000;  wr_data_rom[20000]='h00000000;
    rd_cycle[20001] = 1'b0;  wr_cycle[20001] = 1'b0;  addr_rom[20001]='h00000000;  wr_data_rom[20001]='h00000000;
    rd_cycle[20002] = 1'b0;  wr_cycle[20002] = 1'b0;  addr_rom[20002]='h00000000;  wr_data_rom[20002]='h00000000;
    rd_cycle[20003] = 1'b0;  wr_cycle[20003] = 1'b0;  addr_rom[20003]='h00000000;  wr_data_rom[20003]='h00000000;
    rd_cycle[20004] = 1'b0;  wr_cycle[20004] = 1'b0;  addr_rom[20004]='h00000000;  wr_data_rom[20004]='h00000000;
    rd_cycle[20005] = 1'b0;  wr_cycle[20005] = 1'b0;  addr_rom[20005]='h00000000;  wr_data_rom[20005]='h00000000;
    rd_cycle[20006] = 1'b0;  wr_cycle[20006] = 1'b0;  addr_rom[20006]='h00000000;  wr_data_rom[20006]='h00000000;
    rd_cycle[20007] = 1'b0;  wr_cycle[20007] = 1'b0;  addr_rom[20007]='h00000000;  wr_data_rom[20007]='h00000000;
    rd_cycle[20008] = 1'b0;  wr_cycle[20008] = 1'b0;  addr_rom[20008]='h00000000;  wr_data_rom[20008]='h00000000;
    rd_cycle[20009] = 1'b0;  wr_cycle[20009] = 1'b0;  addr_rom[20009]='h00000000;  wr_data_rom[20009]='h00000000;
    rd_cycle[20010] = 1'b0;  wr_cycle[20010] = 1'b0;  addr_rom[20010]='h00000000;  wr_data_rom[20010]='h00000000;
    rd_cycle[20011] = 1'b0;  wr_cycle[20011] = 1'b0;  addr_rom[20011]='h00000000;  wr_data_rom[20011]='h00000000;
    rd_cycle[20012] = 1'b0;  wr_cycle[20012] = 1'b0;  addr_rom[20012]='h00000000;  wr_data_rom[20012]='h00000000;
    rd_cycle[20013] = 1'b0;  wr_cycle[20013] = 1'b0;  addr_rom[20013]='h00000000;  wr_data_rom[20013]='h00000000;
    rd_cycle[20014] = 1'b0;  wr_cycle[20014] = 1'b0;  addr_rom[20014]='h00000000;  wr_data_rom[20014]='h00000000;
    rd_cycle[20015] = 1'b0;  wr_cycle[20015] = 1'b0;  addr_rom[20015]='h00000000;  wr_data_rom[20015]='h00000000;
    rd_cycle[20016] = 1'b0;  wr_cycle[20016] = 1'b0;  addr_rom[20016]='h00000000;  wr_data_rom[20016]='h00000000;
    rd_cycle[20017] = 1'b0;  wr_cycle[20017] = 1'b0;  addr_rom[20017]='h00000000;  wr_data_rom[20017]='h00000000;
    rd_cycle[20018] = 1'b0;  wr_cycle[20018] = 1'b0;  addr_rom[20018]='h00000000;  wr_data_rom[20018]='h00000000;
    rd_cycle[20019] = 1'b0;  wr_cycle[20019] = 1'b0;  addr_rom[20019]='h00000000;  wr_data_rom[20019]='h00000000;
    rd_cycle[20020] = 1'b0;  wr_cycle[20020] = 1'b0;  addr_rom[20020]='h00000000;  wr_data_rom[20020]='h00000000;
    rd_cycle[20021] = 1'b0;  wr_cycle[20021] = 1'b0;  addr_rom[20021]='h00000000;  wr_data_rom[20021]='h00000000;
    rd_cycle[20022] = 1'b0;  wr_cycle[20022] = 1'b0;  addr_rom[20022]='h00000000;  wr_data_rom[20022]='h00000000;
    rd_cycle[20023] = 1'b0;  wr_cycle[20023] = 1'b0;  addr_rom[20023]='h00000000;  wr_data_rom[20023]='h00000000;
    rd_cycle[20024] = 1'b0;  wr_cycle[20024] = 1'b0;  addr_rom[20024]='h00000000;  wr_data_rom[20024]='h00000000;
    rd_cycle[20025] = 1'b0;  wr_cycle[20025] = 1'b0;  addr_rom[20025]='h00000000;  wr_data_rom[20025]='h00000000;
    rd_cycle[20026] = 1'b0;  wr_cycle[20026] = 1'b0;  addr_rom[20026]='h00000000;  wr_data_rom[20026]='h00000000;
    rd_cycle[20027] = 1'b0;  wr_cycle[20027] = 1'b0;  addr_rom[20027]='h00000000;  wr_data_rom[20027]='h00000000;
    rd_cycle[20028] = 1'b0;  wr_cycle[20028] = 1'b0;  addr_rom[20028]='h00000000;  wr_data_rom[20028]='h00000000;
    rd_cycle[20029] = 1'b0;  wr_cycle[20029] = 1'b0;  addr_rom[20029]='h00000000;  wr_data_rom[20029]='h00000000;
    rd_cycle[20030] = 1'b0;  wr_cycle[20030] = 1'b0;  addr_rom[20030]='h00000000;  wr_data_rom[20030]='h00000000;
    rd_cycle[20031] = 1'b0;  wr_cycle[20031] = 1'b0;  addr_rom[20031]='h00000000;  wr_data_rom[20031]='h00000000;
    rd_cycle[20032] = 1'b0;  wr_cycle[20032] = 1'b0;  addr_rom[20032]='h00000000;  wr_data_rom[20032]='h00000000;
    rd_cycle[20033] = 1'b0;  wr_cycle[20033] = 1'b0;  addr_rom[20033]='h00000000;  wr_data_rom[20033]='h00000000;
    rd_cycle[20034] = 1'b0;  wr_cycle[20034] = 1'b0;  addr_rom[20034]='h00000000;  wr_data_rom[20034]='h00000000;
    rd_cycle[20035] = 1'b0;  wr_cycle[20035] = 1'b0;  addr_rom[20035]='h00000000;  wr_data_rom[20035]='h00000000;
    rd_cycle[20036] = 1'b0;  wr_cycle[20036] = 1'b0;  addr_rom[20036]='h00000000;  wr_data_rom[20036]='h00000000;
    rd_cycle[20037] = 1'b0;  wr_cycle[20037] = 1'b0;  addr_rom[20037]='h00000000;  wr_data_rom[20037]='h00000000;
    rd_cycle[20038] = 1'b0;  wr_cycle[20038] = 1'b0;  addr_rom[20038]='h00000000;  wr_data_rom[20038]='h00000000;
    rd_cycle[20039] = 1'b0;  wr_cycle[20039] = 1'b0;  addr_rom[20039]='h00000000;  wr_data_rom[20039]='h00000000;
    rd_cycle[20040] = 1'b0;  wr_cycle[20040] = 1'b0;  addr_rom[20040]='h00000000;  wr_data_rom[20040]='h00000000;
    rd_cycle[20041] = 1'b0;  wr_cycle[20041] = 1'b0;  addr_rom[20041]='h00000000;  wr_data_rom[20041]='h00000000;
    rd_cycle[20042] = 1'b0;  wr_cycle[20042] = 1'b0;  addr_rom[20042]='h00000000;  wr_data_rom[20042]='h00000000;
    rd_cycle[20043] = 1'b0;  wr_cycle[20043] = 1'b0;  addr_rom[20043]='h00000000;  wr_data_rom[20043]='h00000000;
    rd_cycle[20044] = 1'b0;  wr_cycle[20044] = 1'b0;  addr_rom[20044]='h00000000;  wr_data_rom[20044]='h00000000;
    rd_cycle[20045] = 1'b0;  wr_cycle[20045] = 1'b0;  addr_rom[20045]='h00000000;  wr_data_rom[20045]='h00000000;
    rd_cycle[20046] = 1'b0;  wr_cycle[20046] = 1'b0;  addr_rom[20046]='h00000000;  wr_data_rom[20046]='h00000000;
    rd_cycle[20047] = 1'b0;  wr_cycle[20047] = 1'b0;  addr_rom[20047]='h00000000;  wr_data_rom[20047]='h00000000;
    rd_cycle[20048] = 1'b0;  wr_cycle[20048] = 1'b0;  addr_rom[20048]='h00000000;  wr_data_rom[20048]='h00000000;
    rd_cycle[20049] = 1'b0;  wr_cycle[20049] = 1'b0;  addr_rom[20049]='h00000000;  wr_data_rom[20049]='h00000000;
    rd_cycle[20050] = 1'b0;  wr_cycle[20050] = 1'b0;  addr_rom[20050]='h00000000;  wr_data_rom[20050]='h00000000;
    rd_cycle[20051] = 1'b0;  wr_cycle[20051] = 1'b0;  addr_rom[20051]='h00000000;  wr_data_rom[20051]='h00000000;
    rd_cycle[20052] = 1'b0;  wr_cycle[20052] = 1'b0;  addr_rom[20052]='h00000000;  wr_data_rom[20052]='h00000000;
    rd_cycle[20053] = 1'b0;  wr_cycle[20053] = 1'b0;  addr_rom[20053]='h00000000;  wr_data_rom[20053]='h00000000;
    rd_cycle[20054] = 1'b0;  wr_cycle[20054] = 1'b0;  addr_rom[20054]='h00000000;  wr_data_rom[20054]='h00000000;
    rd_cycle[20055] = 1'b0;  wr_cycle[20055] = 1'b0;  addr_rom[20055]='h00000000;  wr_data_rom[20055]='h00000000;
    rd_cycle[20056] = 1'b0;  wr_cycle[20056] = 1'b0;  addr_rom[20056]='h00000000;  wr_data_rom[20056]='h00000000;
    rd_cycle[20057] = 1'b0;  wr_cycle[20057] = 1'b0;  addr_rom[20057]='h00000000;  wr_data_rom[20057]='h00000000;
    rd_cycle[20058] = 1'b0;  wr_cycle[20058] = 1'b0;  addr_rom[20058]='h00000000;  wr_data_rom[20058]='h00000000;
    rd_cycle[20059] = 1'b0;  wr_cycle[20059] = 1'b0;  addr_rom[20059]='h00000000;  wr_data_rom[20059]='h00000000;
    rd_cycle[20060] = 1'b0;  wr_cycle[20060] = 1'b0;  addr_rom[20060]='h00000000;  wr_data_rom[20060]='h00000000;
    rd_cycle[20061] = 1'b0;  wr_cycle[20061] = 1'b0;  addr_rom[20061]='h00000000;  wr_data_rom[20061]='h00000000;
    rd_cycle[20062] = 1'b0;  wr_cycle[20062] = 1'b0;  addr_rom[20062]='h00000000;  wr_data_rom[20062]='h00000000;
    rd_cycle[20063] = 1'b0;  wr_cycle[20063] = 1'b0;  addr_rom[20063]='h00000000;  wr_data_rom[20063]='h00000000;
    rd_cycle[20064] = 1'b0;  wr_cycle[20064] = 1'b0;  addr_rom[20064]='h00000000;  wr_data_rom[20064]='h00000000;
    rd_cycle[20065] = 1'b0;  wr_cycle[20065] = 1'b0;  addr_rom[20065]='h00000000;  wr_data_rom[20065]='h00000000;
    rd_cycle[20066] = 1'b0;  wr_cycle[20066] = 1'b0;  addr_rom[20066]='h00000000;  wr_data_rom[20066]='h00000000;
    rd_cycle[20067] = 1'b0;  wr_cycle[20067] = 1'b0;  addr_rom[20067]='h00000000;  wr_data_rom[20067]='h00000000;
    rd_cycle[20068] = 1'b0;  wr_cycle[20068] = 1'b0;  addr_rom[20068]='h00000000;  wr_data_rom[20068]='h00000000;
    rd_cycle[20069] = 1'b0;  wr_cycle[20069] = 1'b0;  addr_rom[20069]='h00000000;  wr_data_rom[20069]='h00000000;
    rd_cycle[20070] = 1'b0;  wr_cycle[20070] = 1'b0;  addr_rom[20070]='h00000000;  wr_data_rom[20070]='h00000000;
    rd_cycle[20071] = 1'b0;  wr_cycle[20071] = 1'b0;  addr_rom[20071]='h00000000;  wr_data_rom[20071]='h00000000;
    rd_cycle[20072] = 1'b0;  wr_cycle[20072] = 1'b0;  addr_rom[20072]='h00000000;  wr_data_rom[20072]='h00000000;
    rd_cycle[20073] = 1'b0;  wr_cycle[20073] = 1'b0;  addr_rom[20073]='h00000000;  wr_data_rom[20073]='h00000000;
    rd_cycle[20074] = 1'b0;  wr_cycle[20074] = 1'b0;  addr_rom[20074]='h00000000;  wr_data_rom[20074]='h00000000;
    rd_cycle[20075] = 1'b0;  wr_cycle[20075] = 1'b0;  addr_rom[20075]='h00000000;  wr_data_rom[20075]='h00000000;
    rd_cycle[20076] = 1'b0;  wr_cycle[20076] = 1'b0;  addr_rom[20076]='h00000000;  wr_data_rom[20076]='h00000000;
    rd_cycle[20077] = 1'b0;  wr_cycle[20077] = 1'b0;  addr_rom[20077]='h00000000;  wr_data_rom[20077]='h00000000;
    rd_cycle[20078] = 1'b0;  wr_cycle[20078] = 1'b0;  addr_rom[20078]='h00000000;  wr_data_rom[20078]='h00000000;
    rd_cycle[20079] = 1'b0;  wr_cycle[20079] = 1'b0;  addr_rom[20079]='h00000000;  wr_data_rom[20079]='h00000000;
    rd_cycle[20080] = 1'b0;  wr_cycle[20080] = 1'b0;  addr_rom[20080]='h00000000;  wr_data_rom[20080]='h00000000;
    rd_cycle[20081] = 1'b0;  wr_cycle[20081] = 1'b0;  addr_rom[20081]='h00000000;  wr_data_rom[20081]='h00000000;
    rd_cycle[20082] = 1'b0;  wr_cycle[20082] = 1'b0;  addr_rom[20082]='h00000000;  wr_data_rom[20082]='h00000000;
    rd_cycle[20083] = 1'b0;  wr_cycle[20083] = 1'b0;  addr_rom[20083]='h00000000;  wr_data_rom[20083]='h00000000;
    rd_cycle[20084] = 1'b0;  wr_cycle[20084] = 1'b0;  addr_rom[20084]='h00000000;  wr_data_rom[20084]='h00000000;
    rd_cycle[20085] = 1'b0;  wr_cycle[20085] = 1'b0;  addr_rom[20085]='h00000000;  wr_data_rom[20085]='h00000000;
    rd_cycle[20086] = 1'b0;  wr_cycle[20086] = 1'b0;  addr_rom[20086]='h00000000;  wr_data_rom[20086]='h00000000;
    rd_cycle[20087] = 1'b0;  wr_cycle[20087] = 1'b0;  addr_rom[20087]='h00000000;  wr_data_rom[20087]='h00000000;
    rd_cycle[20088] = 1'b0;  wr_cycle[20088] = 1'b0;  addr_rom[20088]='h00000000;  wr_data_rom[20088]='h00000000;
    rd_cycle[20089] = 1'b0;  wr_cycle[20089] = 1'b0;  addr_rom[20089]='h00000000;  wr_data_rom[20089]='h00000000;
    rd_cycle[20090] = 1'b0;  wr_cycle[20090] = 1'b0;  addr_rom[20090]='h00000000;  wr_data_rom[20090]='h00000000;
    rd_cycle[20091] = 1'b0;  wr_cycle[20091] = 1'b0;  addr_rom[20091]='h00000000;  wr_data_rom[20091]='h00000000;
    rd_cycle[20092] = 1'b0;  wr_cycle[20092] = 1'b0;  addr_rom[20092]='h00000000;  wr_data_rom[20092]='h00000000;
    rd_cycle[20093] = 1'b0;  wr_cycle[20093] = 1'b0;  addr_rom[20093]='h00000000;  wr_data_rom[20093]='h00000000;
    rd_cycle[20094] = 1'b0;  wr_cycle[20094] = 1'b0;  addr_rom[20094]='h00000000;  wr_data_rom[20094]='h00000000;
    rd_cycle[20095] = 1'b0;  wr_cycle[20095] = 1'b0;  addr_rom[20095]='h00000000;  wr_data_rom[20095]='h00000000;
    rd_cycle[20096] = 1'b0;  wr_cycle[20096] = 1'b0;  addr_rom[20096]='h00000000;  wr_data_rom[20096]='h00000000;
    rd_cycle[20097] = 1'b0;  wr_cycle[20097] = 1'b0;  addr_rom[20097]='h00000000;  wr_data_rom[20097]='h00000000;
    rd_cycle[20098] = 1'b0;  wr_cycle[20098] = 1'b0;  addr_rom[20098]='h00000000;  wr_data_rom[20098]='h00000000;
    rd_cycle[20099] = 1'b0;  wr_cycle[20099] = 1'b0;  addr_rom[20099]='h00000000;  wr_data_rom[20099]='h00000000;
    rd_cycle[20100] = 1'b0;  wr_cycle[20100] = 1'b0;  addr_rom[20100]='h00000000;  wr_data_rom[20100]='h00000000;
    rd_cycle[20101] = 1'b0;  wr_cycle[20101] = 1'b0;  addr_rom[20101]='h00000000;  wr_data_rom[20101]='h00000000;
    rd_cycle[20102] = 1'b0;  wr_cycle[20102] = 1'b0;  addr_rom[20102]='h00000000;  wr_data_rom[20102]='h00000000;
    rd_cycle[20103] = 1'b0;  wr_cycle[20103] = 1'b0;  addr_rom[20103]='h00000000;  wr_data_rom[20103]='h00000000;
    rd_cycle[20104] = 1'b0;  wr_cycle[20104] = 1'b0;  addr_rom[20104]='h00000000;  wr_data_rom[20104]='h00000000;
    rd_cycle[20105] = 1'b0;  wr_cycle[20105] = 1'b0;  addr_rom[20105]='h00000000;  wr_data_rom[20105]='h00000000;
    rd_cycle[20106] = 1'b0;  wr_cycle[20106] = 1'b0;  addr_rom[20106]='h00000000;  wr_data_rom[20106]='h00000000;
    rd_cycle[20107] = 1'b0;  wr_cycle[20107] = 1'b0;  addr_rom[20107]='h00000000;  wr_data_rom[20107]='h00000000;
    rd_cycle[20108] = 1'b0;  wr_cycle[20108] = 1'b0;  addr_rom[20108]='h00000000;  wr_data_rom[20108]='h00000000;
    rd_cycle[20109] = 1'b0;  wr_cycle[20109] = 1'b0;  addr_rom[20109]='h00000000;  wr_data_rom[20109]='h00000000;
    rd_cycle[20110] = 1'b0;  wr_cycle[20110] = 1'b0;  addr_rom[20110]='h00000000;  wr_data_rom[20110]='h00000000;
    rd_cycle[20111] = 1'b0;  wr_cycle[20111] = 1'b0;  addr_rom[20111]='h00000000;  wr_data_rom[20111]='h00000000;
    rd_cycle[20112] = 1'b0;  wr_cycle[20112] = 1'b0;  addr_rom[20112]='h00000000;  wr_data_rom[20112]='h00000000;
    rd_cycle[20113] = 1'b0;  wr_cycle[20113] = 1'b0;  addr_rom[20113]='h00000000;  wr_data_rom[20113]='h00000000;
    rd_cycle[20114] = 1'b0;  wr_cycle[20114] = 1'b0;  addr_rom[20114]='h00000000;  wr_data_rom[20114]='h00000000;
    rd_cycle[20115] = 1'b0;  wr_cycle[20115] = 1'b0;  addr_rom[20115]='h00000000;  wr_data_rom[20115]='h00000000;
    rd_cycle[20116] = 1'b0;  wr_cycle[20116] = 1'b0;  addr_rom[20116]='h00000000;  wr_data_rom[20116]='h00000000;
    rd_cycle[20117] = 1'b0;  wr_cycle[20117] = 1'b0;  addr_rom[20117]='h00000000;  wr_data_rom[20117]='h00000000;
    rd_cycle[20118] = 1'b0;  wr_cycle[20118] = 1'b0;  addr_rom[20118]='h00000000;  wr_data_rom[20118]='h00000000;
    rd_cycle[20119] = 1'b0;  wr_cycle[20119] = 1'b0;  addr_rom[20119]='h00000000;  wr_data_rom[20119]='h00000000;
    rd_cycle[20120] = 1'b0;  wr_cycle[20120] = 1'b0;  addr_rom[20120]='h00000000;  wr_data_rom[20120]='h00000000;
    rd_cycle[20121] = 1'b0;  wr_cycle[20121] = 1'b0;  addr_rom[20121]='h00000000;  wr_data_rom[20121]='h00000000;
    rd_cycle[20122] = 1'b0;  wr_cycle[20122] = 1'b0;  addr_rom[20122]='h00000000;  wr_data_rom[20122]='h00000000;
    rd_cycle[20123] = 1'b0;  wr_cycle[20123] = 1'b0;  addr_rom[20123]='h00000000;  wr_data_rom[20123]='h00000000;
    rd_cycle[20124] = 1'b0;  wr_cycle[20124] = 1'b0;  addr_rom[20124]='h00000000;  wr_data_rom[20124]='h00000000;
    rd_cycle[20125] = 1'b0;  wr_cycle[20125] = 1'b0;  addr_rom[20125]='h00000000;  wr_data_rom[20125]='h00000000;
    rd_cycle[20126] = 1'b0;  wr_cycle[20126] = 1'b0;  addr_rom[20126]='h00000000;  wr_data_rom[20126]='h00000000;
    rd_cycle[20127] = 1'b0;  wr_cycle[20127] = 1'b0;  addr_rom[20127]='h00000000;  wr_data_rom[20127]='h00000000;
    rd_cycle[20128] = 1'b0;  wr_cycle[20128] = 1'b0;  addr_rom[20128]='h00000000;  wr_data_rom[20128]='h00000000;
    rd_cycle[20129] = 1'b0;  wr_cycle[20129] = 1'b0;  addr_rom[20129]='h00000000;  wr_data_rom[20129]='h00000000;
    rd_cycle[20130] = 1'b0;  wr_cycle[20130] = 1'b0;  addr_rom[20130]='h00000000;  wr_data_rom[20130]='h00000000;
    rd_cycle[20131] = 1'b0;  wr_cycle[20131] = 1'b0;  addr_rom[20131]='h00000000;  wr_data_rom[20131]='h00000000;
    rd_cycle[20132] = 1'b0;  wr_cycle[20132] = 1'b0;  addr_rom[20132]='h00000000;  wr_data_rom[20132]='h00000000;
    rd_cycle[20133] = 1'b0;  wr_cycle[20133] = 1'b0;  addr_rom[20133]='h00000000;  wr_data_rom[20133]='h00000000;
    rd_cycle[20134] = 1'b0;  wr_cycle[20134] = 1'b0;  addr_rom[20134]='h00000000;  wr_data_rom[20134]='h00000000;
    rd_cycle[20135] = 1'b0;  wr_cycle[20135] = 1'b0;  addr_rom[20135]='h00000000;  wr_data_rom[20135]='h00000000;
    rd_cycle[20136] = 1'b0;  wr_cycle[20136] = 1'b0;  addr_rom[20136]='h00000000;  wr_data_rom[20136]='h00000000;
    rd_cycle[20137] = 1'b0;  wr_cycle[20137] = 1'b0;  addr_rom[20137]='h00000000;  wr_data_rom[20137]='h00000000;
    rd_cycle[20138] = 1'b0;  wr_cycle[20138] = 1'b0;  addr_rom[20138]='h00000000;  wr_data_rom[20138]='h00000000;
    rd_cycle[20139] = 1'b0;  wr_cycle[20139] = 1'b0;  addr_rom[20139]='h00000000;  wr_data_rom[20139]='h00000000;
    rd_cycle[20140] = 1'b0;  wr_cycle[20140] = 1'b0;  addr_rom[20140]='h00000000;  wr_data_rom[20140]='h00000000;
    rd_cycle[20141] = 1'b0;  wr_cycle[20141] = 1'b0;  addr_rom[20141]='h00000000;  wr_data_rom[20141]='h00000000;
    rd_cycle[20142] = 1'b0;  wr_cycle[20142] = 1'b0;  addr_rom[20142]='h00000000;  wr_data_rom[20142]='h00000000;
    rd_cycle[20143] = 1'b0;  wr_cycle[20143] = 1'b0;  addr_rom[20143]='h00000000;  wr_data_rom[20143]='h00000000;
    rd_cycle[20144] = 1'b0;  wr_cycle[20144] = 1'b0;  addr_rom[20144]='h00000000;  wr_data_rom[20144]='h00000000;
    rd_cycle[20145] = 1'b0;  wr_cycle[20145] = 1'b0;  addr_rom[20145]='h00000000;  wr_data_rom[20145]='h00000000;
    rd_cycle[20146] = 1'b0;  wr_cycle[20146] = 1'b0;  addr_rom[20146]='h00000000;  wr_data_rom[20146]='h00000000;
    rd_cycle[20147] = 1'b0;  wr_cycle[20147] = 1'b0;  addr_rom[20147]='h00000000;  wr_data_rom[20147]='h00000000;
    rd_cycle[20148] = 1'b0;  wr_cycle[20148] = 1'b0;  addr_rom[20148]='h00000000;  wr_data_rom[20148]='h00000000;
    rd_cycle[20149] = 1'b0;  wr_cycle[20149] = 1'b0;  addr_rom[20149]='h00000000;  wr_data_rom[20149]='h00000000;
    rd_cycle[20150] = 1'b0;  wr_cycle[20150] = 1'b0;  addr_rom[20150]='h00000000;  wr_data_rom[20150]='h00000000;
    rd_cycle[20151] = 1'b0;  wr_cycle[20151] = 1'b0;  addr_rom[20151]='h00000000;  wr_data_rom[20151]='h00000000;
    rd_cycle[20152] = 1'b0;  wr_cycle[20152] = 1'b0;  addr_rom[20152]='h00000000;  wr_data_rom[20152]='h00000000;
    rd_cycle[20153] = 1'b0;  wr_cycle[20153] = 1'b0;  addr_rom[20153]='h00000000;  wr_data_rom[20153]='h00000000;
    rd_cycle[20154] = 1'b0;  wr_cycle[20154] = 1'b0;  addr_rom[20154]='h00000000;  wr_data_rom[20154]='h00000000;
    rd_cycle[20155] = 1'b0;  wr_cycle[20155] = 1'b0;  addr_rom[20155]='h00000000;  wr_data_rom[20155]='h00000000;
    rd_cycle[20156] = 1'b0;  wr_cycle[20156] = 1'b0;  addr_rom[20156]='h00000000;  wr_data_rom[20156]='h00000000;
    rd_cycle[20157] = 1'b0;  wr_cycle[20157] = 1'b0;  addr_rom[20157]='h00000000;  wr_data_rom[20157]='h00000000;
    rd_cycle[20158] = 1'b0;  wr_cycle[20158] = 1'b0;  addr_rom[20158]='h00000000;  wr_data_rom[20158]='h00000000;
    rd_cycle[20159] = 1'b0;  wr_cycle[20159] = 1'b0;  addr_rom[20159]='h00000000;  wr_data_rom[20159]='h00000000;
    rd_cycle[20160] = 1'b0;  wr_cycle[20160] = 1'b0;  addr_rom[20160]='h00000000;  wr_data_rom[20160]='h00000000;
    rd_cycle[20161] = 1'b0;  wr_cycle[20161] = 1'b0;  addr_rom[20161]='h00000000;  wr_data_rom[20161]='h00000000;
    rd_cycle[20162] = 1'b0;  wr_cycle[20162] = 1'b0;  addr_rom[20162]='h00000000;  wr_data_rom[20162]='h00000000;
    rd_cycle[20163] = 1'b0;  wr_cycle[20163] = 1'b0;  addr_rom[20163]='h00000000;  wr_data_rom[20163]='h00000000;
    rd_cycle[20164] = 1'b0;  wr_cycle[20164] = 1'b0;  addr_rom[20164]='h00000000;  wr_data_rom[20164]='h00000000;
    rd_cycle[20165] = 1'b0;  wr_cycle[20165] = 1'b0;  addr_rom[20165]='h00000000;  wr_data_rom[20165]='h00000000;
    rd_cycle[20166] = 1'b0;  wr_cycle[20166] = 1'b0;  addr_rom[20166]='h00000000;  wr_data_rom[20166]='h00000000;
    rd_cycle[20167] = 1'b0;  wr_cycle[20167] = 1'b0;  addr_rom[20167]='h00000000;  wr_data_rom[20167]='h00000000;
    rd_cycle[20168] = 1'b0;  wr_cycle[20168] = 1'b0;  addr_rom[20168]='h00000000;  wr_data_rom[20168]='h00000000;
    rd_cycle[20169] = 1'b0;  wr_cycle[20169] = 1'b0;  addr_rom[20169]='h00000000;  wr_data_rom[20169]='h00000000;
    rd_cycle[20170] = 1'b0;  wr_cycle[20170] = 1'b0;  addr_rom[20170]='h00000000;  wr_data_rom[20170]='h00000000;
    rd_cycle[20171] = 1'b0;  wr_cycle[20171] = 1'b0;  addr_rom[20171]='h00000000;  wr_data_rom[20171]='h00000000;
    rd_cycle[20172] = 1'b0;  wr_cycle[20172] = 1'b0;  addr_rom[20172]='h00000000;  wr_data_rom[20172]='h00000000;
    rd_cycle[20173] = 1'b0;  wr_cycle[20173] = 1'b0;  addr_rom[20173]='h00000000;  wr_data_rom[20173]='h00000000;
    rd_cycle[20174] = 1'b0;  wr_cycle[20174] = 1'b0;  addr_rom[20174]='h00000000;  wr_data_rom[20174]='h00000000;
    rd_cycle[20175] = 1'b0;  wr_cycle[20175] = 1'b0;  addr_rom[20175]='h00000000;  wr_data_rom[20175]='h00000000;
    rd_cycle[20176] = 1'b0;  wr_cycle[20176] = 1'b0;  addr_rom[20176]='h00000000;  wr_data_rom[20176]='h00000000;
    rd_cycle[20177] = 1'b0;  wr_cycle[20177] = 1'b0;  addr_rom[20177]='h00000000;  wr_data_rom[20177]='h00000000;
    rd_cycle[20178] = 1'b0;  wr_cycle[20178] = 1'b0;  addr_rom[20178]='h00000000;  wr_data_rom[20178]='h00000000;
    rd_cycle[20179] = 1'b0;  wr_cycle[20179] = 1'b0;  addr_rom[20179]='h00000000;  wr_data_rom[20179]='h00000000;
    rd_cycle[20180] = 1'b0;  wr_cycle[20180] = 1'b0;  addr_rom[20180]='h00000000;  wr_data_rom[20180]='h00000000;
    rd_cycle[20181] = 1'b0;  wr_cycle[20181] = 1'b0;  addr_rom[20181]='h00000000;  wr_data_rom[20181]='h00000000;
    rd_cycle[20182] = 1'b0;  wr_cycle[20182] = 1'b0;  addr_rom[20182]='h00000000;  wr_data_rom[20182]='h00000000;
    rd_cycle[20183] = 1'b0;  wr_cycle[20183] = 1'b0;  addr_rom[20183]='h00000000;  wr_data_rom[20183]='h00000000;
    rd_cycle[20184] = 1'b0;  wr_cycle[20184] = 1'b0;  addr_rom[20184]='h00000000;  wr_data_rom[20184]='h00000000;
    rd_cycle[20185] = 1'b0;  wr_cycle[20185] = 1'b0;  addr_rom[20185]='h00000000;  wr_data_rom[20185]='h00000000;
    rd_cycle[20186] = 1'b0;  wr_cycle[20186] = 1'b0;  addr_rom[20186]='h00000000;  wr_data_rom[20186]='h00000000;
    rd_cycle[20187] = 1'b0;  wr_cycle[20187] = 1'b0;  addr_rom[20187]='h00000000;  wr_data_rom[20187]='h00000000;
    rd_cycle[20188] = 1'b0;  wr_cycle[20188] = 1'b0;  addr_rom[20188]='h00000000;  wr_data_rom[20188]='h00000000;
    rd_cycle[20189] = 1'b0;  wr_cycle[20189] = 1'b0;  addr_rom[20189]='h00000000;  wr_data_rom[20189]='h00000000;
    rd_cycle[20190] = 1'b0;  wr_cycle[20190] = 1'b0;  addr_rom[20190]='h00000000;  wr_data_rom[20190]='h00000000;
    rd_cycle[20191] = 1'b0;  wr_cycle[20191] = 1'b0;  addr_rom[20191]='h00000000;  wr_data_rom[20191]='h00000000;
    rd_cycle[20192] = 1'b0;  wr_cycle[20192] = 1'b0;  addr_rom[20192]='h00000000;  wr_data_rom[20192]='h00000000;
    rd_cycle[20193] = 1'b0;  wr_cycle[20193] = 1'b0;  addr_rom[20193]='h00000000;  wr_data_rom[20193]='h00000000;
    rd_cycle[20194] = 1'b0;  wr_cycle[20194] = 1'b0;  addr_rom[20194]='h00000000;  wr_data_rom[20194]='h00000000;
    rd_cycle[20195] = 1'b0;  wr_cycle[20195] = 1'b0;  addr_rom[20195]='h00000000;  wr_data_rom[20195]='h00000000;
    rd_cycle[20196] = 1'b0;  wr_cycle[20196] = 1'b0;  addr_rom[20196]='h00000000;  wr_data_rom[20196]='h00000000;
    rd_cycle[20197] = 1'b0;  wr_cycle[20197] = 1'b0;  addr_rom[20197]='h00000000;  wr_data_rom[20197]='h00000000;
    rd_cycle[20198] = 1'b0;  wr_cycle[20198] = 1'b0;  addr_rom[20198]='h00000000;  wr_data_rom[20198]='h00000000;
    rd_cycle[20199] = 1'b0;  wr_cycle[20199] = 1'b0;  addr_rom[20199]='h00000000;  wr_data_rom[20199]='h00000000;
    rd_cycle[20200] = 1'b0;  wr_cycle[20200] = 1'b0;  addr_rom[20200]='h00000000;  wr_data_rom[20200]='h00000000;
    rd_cycle[20201] = 1'b0;  wr_cycle[20201] = 1'b0;  addr_rom[20201]='h00000000;  wr_data_rom[20201]='h00000000;
    rd_cycle[20202] = 1'b0;  wr_cycle[20202] = 1'b0;  addr_rom[20202]='h00000000;  wr_data_rom[20202]='h00000000;
    rd_cycle[20203] = 1'b0;  wr_cycle[20203] = 1'b0;  addr_rom[20203]='h00000000;  wr_data_rom[20203]='h00000000;
    rd_cycle[20204] = 1'b0;  wr_cycle[20204] = 1'b0;  addr_rom[20204]='h00000000;  wr_data_rom[20204]='h00000000;
    rd_cycle[20205] = 1'b0;  wr_cycle[20205] = 1'b0;  addr_rom[20205]='h00000000;  wr_data_rom[20205]='h00000000;
    rd_cycle[20206] = 1'b0;  wr_cycle[20206] = 1'b0;  addr_rom[20206]='h00000000;  wr_data_rom[20206]='h00000000;
    rd_cycle[20207] = 1'b0;  wr_cycle[20207] = 1'b0;  addr_rom[20207]='h00000000;  wr_data_rom[20207]='h00000000;
    rd_cycle[20208] = 1'b0;  wr_cycle[20208] = 1'b0;  addr_rom[20208]='h00000000;  wr_data_rom[20208]='h00000000;
    rd_cycle[20209] = 1'b0;  wr_cycle[20209] = 1'b0;  addr_rom[20209]='h00000000;  wr_data_rom[20209]='h00000000;
    rd_cycle[20210] = 1'b0;  wr_cycle[20210] = 1'b0;  addr_rom[20210]='h00000000;  wr_data_rom[20210]='h00000000;
    rd_cycle[20211] = 1'b0;  wr_cycle[20211] = 1'b0;  addr_rom[20211]='h00000000;  wr_data_rom[20211]='h00000000;
    rd_cycle[20212] = 1'b0;  wr_cycle[20212] = 1'b0;  addr_rom[20212]='h00000000;  wr_data_rom[20212]='h00000000;
    rd_cycle[20213] = 1'b0;  wr_cycle[20213] = 1'b0;  addr_rom[20213]='h00000000;  wr_data_rom[20213]='h00000000;
    rd_cycle[20214] = 1'b0;  wr_cycle[20214] = 1'b0;  addr_rom[20214]='h00000000;  wr_data_rom[20214]='h00000000;
    rd_cycle[20215] = 1'b0;  wr_cycle[20215] = 1'b0;  addr_rom[20215]='h00000000;  wr_data_rom[20215]='h00000000;
    rd_cycle[20216] = 1'b0;  wr_cycle[20216] = 1'b0;  addr_rom[20216]='h00000000;  wr_data_rom[20216]='h00000000;
    rd_cycle[20217] = 1'b0;  wr_cycle[20217] = 1'b0;  addr_rom[20217]='h00000000;  wr_data_rom[20217]='h00000000;
    rd_cycle[20218] = 1'b0;  wr_cycle[20218] = 1'b0;  addr_rom[20218]='h00000000;  wr_data_rom[20218]='h00000000;
    rd_cycle[20219] = 1'b0;  wr_cycle[20219] = 1'b0;  addr_rom[20219]='h00000000;  wr_data_rom[20219]='h00000000;
    rd_cycle[20220] = 1'b0;  wr_cycle[20220] = 1'b0;  addr_rom[20220]='h00000000;  wr_data_rom[20220]='h00000000;
    rd_cycle[20221] = 1'b0;  wr_cycle[20221] = 1'b0;  addr_rom[20221]='h00000000;  wr_data_rom[20221]='h00000000;
    rd_cycle[20222] = 1'b0;  wr_cycle[20222] = 1'b0;  addr_rom[20222]='h00000000;  wr_data_rom[20222]='h00000000;
    rd_cycle[20223] = 1'b0;  wr_cycle[20223] = 1'b0;  addr_rom[20223]='h00000000;  wr_data_rom[20223]='h00000000;
    rd_cycle[20224] = 1'b0;  wr_cycle[20224] = 1'b0;  addr_rom[20224]='h00000000;  wr_data_rom[20224]='h00000000;
    rd_cycle[20225] = 1'b0;  wr_cycle[20225] = 1'b0;  addr_rom[20225]='h00000000;  wr_data_rom[20225]='h00000000;
    rd_cycle[20226] = 1'b0;  wr_cycle[20226] = 1'b0;  addr_rom[20226]='h00000000;  wr_data_rom[20226]='h00000000;
    rd_cycle[20227] = 1'b0;  wr_cycle[20227] = 1'b0;  addr_rom[20227]='h00000000;  wr_data_rom[20227]='h00000000;
    rd_cycle[20228] = 1'b0;  wr_cycle[20228] = 1'b0;  addr_rom[20228]='h00000000;  wr_data_rom[20228]='h00000000;
    rd_cycle[20229] = 1'b0;  wr_cycle[20229] = 1'b0;  addr_rom[20229]='h00000000;  wr_data_rom[20229]='h00000000;
    rd_cycle[20230] = 1'b0;  wr_cycle[20230] = 1'b0;  addr_rom[20230]='h00000000;  wr_data_rom[20230]='h00000000;
    rd_cycle[20231] = 1'b0;  wr_cycle[20231] = 1'b0;  addr_rom[20231]='h00000000;  wr_data_rom[20231]='h00000000;
    rd_cycle[20232] = 1'b0;  wr_cycle[20232] = 1'b0;  addr_rom[20232]='h00000000;  wr_data_rom[20232]='h00000000;
    rd_cycle[20233] = 1'b0;  wr_cycle[20233] = 1'b0;  addr_rom[20233]='h00000000;  wr_data_rom[20233]='h00000000;
    rd_cycle[20234] = 1'b0;  wr_cycle[20234] = 1'b0;  addr_rom[20234]='h00000000;  wr_data_rom[20234]='h00000000;
    rd_cycle[20235] = 1'b0;  wr_cycle[20235] = 1'b0;  addr_rom[20235]='h00000000;  wr_data_rom[20235]='h00000000;
    rd_cycle[20236] = 1'b0;  wr_cycle[20236] = 1'b0;  addr_rom[20236]='h00000000;  wr_data_rom[20236]='h00000000;
    rd_cycle[20237] = 1'b0;  wr_cycle[20237] = 1'b0;  addr_rom[20237]='h00000000;  wr_data_rom[20237]='h00000000;
    rd_cycle[20238] = 1'b0;  wr_cycle[20238] = 1'b0;  addr_rom[20238]='h00000000;  wr_data_rom[20238]='h00000000;
    rd_cycle[20239] = 1'b0;  wr_cycle[20239] = 1'b0;  addr_rom[20239]='h00000000;  wr_data_rom[20239]='h00000000;
    rd_cycle[20240] = 1'b0;  wr_cycle[20240] = 1'b0;  addr_rom[20240]='h00000000;  wr_data_rom[20240]='h00000000;
    rd_cycle[20241] = 1'b0;  wr_cycle[20241] = 1'b0;  addr_rom[20241]='h00000000;  wr_data_rom[20241]='h00000000;
    rd_cycle[20242] = 1'b0;  wr_cycle[20242] = 1'b0;  addr_rom[20242]='h00000000;  wr_data_rom[20242]='h00000000;
    rd_cycle[20243] = 1'b0;  wr_cycle[20243] = 1'b0;  addr_rom[20243]='h00000000;  wr_data_rom[20243]='h00000000;
    rd_cycle[20244] = 1'b0;  wr_cycle[20244] = 1'b0;  addr_rom[20244]='h00000000;  wr_data_rom[20244]='h00000000;
    rd_cycle[20245] = 1'b0;  wr_cycle[20245] = 1'b0;  addr_rom[20245]='h00000000;  wr_data_rom[20245]='h00000000;
    rd_cycle[20246] = 1'b0;  wr_cycle[20246] = 1'b0;  addr_rom[20246]='h00000000;  wr_data_rom[20246]='h00000000;
    rd_cycle[20247] = 1'b0;  wr_cycle[20247] = 1'b0;  addr_rom[20247]='h00000000;  wr_data_rom[20247]='h00000000;
    rd_cycle[20248] = 1'b0;  wr_cycle[20248] = 1'b0;  addr_rom[20248]='h00000000;  wr_data_rom[20248]='h00000000;
    rd_cycle[20249] = 1'b0;  wr_cycle[20249] = 1'b0;  addr_rom[20249]='h00000000;  wr_data_rom[20249]='h00000000;
    rd_cycle[20250] = 1'b0;  wr_cycle[20250] = 1'b0;  addr_rom[20250]='h00000000;  wr_data_rom[20250]='h00000000;
    rd_cycle[20251] = 1'b0;  wr_cycle[20251] = 1'b0;  addr_rom[20251]='h00000000;  wr_data_rom[20251]='h00000000;
    rd_cycle[20252] = 1'b0;  wr_cycle[20252] = 1'b0;  addr_rom[20252]='h00000000;  wr_data_rom[20252]='h00000000;
    rd_cycle[20253] = 1'b0;  wr_cycle[20253] = 1'b0;  addr_rom[20253]='h00000000;  wr_data_rom[20253]='h00000000;
    rd_cycle[20254] = 1'b0;  wr_cycle[20254] = 1'b0;  addr_rom[20254]='h00000000;  wr_data_rom[20254]='h00000000;
    rd_cycle[20255] = 1'b0;  wr_cycle[20255] = 1'b0;  addr_rom[20255]='h00000000;  wr_data_rom[20255]='h00000000;
    rd_cycle[20256] = 1'b0;  wr_cycle[20256] = 1'b0;  addr_rom[20256]='h00000000;  wr_data_rom[20256]='h00000000;
    rd_cycle[20257] = 1'b0;  wr_cycle[20257] = 1'b0;  addr_rom[20257]='h00000000;  wr_data_rom[20257]='h00000000;
    rd_cycle[20258] = 1'b0;  wr_cycle[20258] = 1'b0;  addr_rom[20258]='h00000000;  wr_data_rom[20258]='h00000000;
    rd_cycle[20259] = 1'b0;  wr_cycle[20259] = 1'b0;  addr_rom[20259]='h00000000;  wr_data_rom[20259]='h00000000;
    rd_cycle[20260] = 1'b0;  wr_cycle[20260] = 1'b0;  addr_rom[20260]='h00000000;  wr_data_rom[20260]='h00000000;
    rd_cycle[20261] = 1'b0;  wr_cycle[20261] = 1'b0;  addr_rom[20261]='h00000000;  wr_data_rom[20261]='h00000000;
    rd_cycle[20262] = 1'b0;  wr_cycle[20262] = 1'b0;  addr_rom[20262]='h00000000;  wr_data_rom[20262]='h00000000;
    rd_cycle[20263] = 1'b0;  wr_cycle[20263] = 1'b0;  addr_rom[20263]='h00000000;  wr_data_rom[20263]='h00000000;
    rd_cycle[20264] = 1'b0;  wr_cycle[20264] = 1'b0;  addr_rom[20264]='h00000000;  wr_data_rom[20264]='h00000000;
    rd_cycle[20265] = 1'b0;  wr_cycle[20265] = 1'b0;  addr_rom[20265]='h00000000;  wr_data_rom[20265]='h00000000;
    rd_cycle[20266] = 1'b0;  wr_cycle[20266] = 1'b0;  addr_rom[20266]='h00000000;  wr_data_rom[20266]='h00000000;
    rd_cycle[20267] = 1'b0;  wr_cycle[20267] = 1'b0;  addr_rom[20267]='h00000000;  wr_data_rom[20267]='h00000000;
    rd_cycle[20268] = 1'b0;  wr_cycle[20268] = 1'b0;  addr_rom[20268]='h00000000;  wr_data_rom[20268]='h00000000;
    rd_cycle[20269] = 1'b0;  wr_cycle[20269] = 1'b0;  addr_rom[20269]='h00000000;  wr_data_rom[20269]='h00000000;
    rd_cycle[20270] = 1'b0;  wr_cycle[20270] = 1'b0;  addr_rom[20270]='h00000000;  wr_data_rom[20270]='h00000000;
    rd_cycle[20271] = 1'b0;  wr_cycle[20271] = 1'b0;  addr_rom[20271]='h00000000;  wr_data_rom[20271]='h00000000;
    rd_cycle[20272] = 1'b0;  wr_cycle[20272] = 1'b0;  addr_rom[20272]='h00000000;  wr_data_rom[20272]='h00000000;
    rd_cycle[20273] = 1'b0;  wr_cycle[20273] = 1'b0;  addr_rom[20273]='h00000000;  wr_data_rom[20273]='h00000000;
    rd_cycle[20274] = 1'b0;  wr_cycle[20274] = 1'b0;  addr_rom[20274]='h00000000;  wr_data_rom[20274]='h00000000;
    rd_cycle[20275] = 1'b0;  wr_cycle[20275] = 1'b0;  addr_rom[20275]='h00000000;  wr_data_rom[20275]='h00000000;
    rd_cycle[20276] = 1'b0;  wr_cycle[20276] = 1'b0;  addr_rom[20276]='h00000000;  wr_data_rom[20276]='h00000000;
    rd_cycle[20277] = 1'b0;  wr_cycle[20277] = 1'b0;  addr_rom[20277]='h00000000;  wr_data_rom[20277]='h00000000;
    rd_cycle[20278] = 1'b0;  wr_cycle[20278] = 1'b0;  addr_rom[20278]='h00000000;  wr_data_rom[20278]='h00000000;
    rd_cycle[20279] = 1'b0;  wr_cycle[20279] = 1'b0;  addr_rom[20279]='h00000000;  wr_data_rom[20279]='h00000000;
    rd_cycle[20280] = 1'b0;  wr_cycle[20280] = 1'b0;  addr_rom[20280]='h00000000;  wr_data_rom[20280]='h00000000;
    rd_cycle[20281] = 1'b0;  wr_cycle[20281] = 1'b0;  addr_rom[20281]='h00000000;  wr_data_rom[20281]='h00000000;
    rd_cycle[20282] = 1'b0;  wr_cycle[20282] = 1'b0;  addr_rom[20282]='h00000000;  wr_data_rom[20282]='h00000000;
    rd_cycle[20283] = 1'b0;  wr_cycle[20283] = 1'b0;  addr_rom[20283]='h00000000;  wr_data_rom[20283]='h00000000;
    rd_cycle[20284] = 1'b0;  wr_cycle[20284] = 1'b0;  addr_rom[20284]='h00000000;  wr_data_rom[20284]='h00000000;
    rd_cycle[20285] = 1'b0;  wr_cycle[20285] = 1'b0;  addr_rom[20285]='h00000000;  wr_data_rom[20285]='h00000000;
    rd_cycle[20286] = 1'b0;  wr_cycle[20286] = 1'b0;  addr_rom[20286]='h00000000;  wr_data_rom[20286]='h00000000;
    rd_cycle[20287] = 1'b0;  wr_cycle[20287] = 1'b0;  addr_rom[20287]='h00000000;  wr_data_rom[20287]='h00000000;
    rd_cycle[20288] = 1'b0;  wr_cycle[20288] = 1'b0;  addr_rom[20288]='h00000000;  wr_data_rom[20288]='h00000000;
    rd_cycle[20289] = 1'b0;  wr_cycle[20289] = 1'b0;  addr_rom[20289]='h00000000;  wr_data_rom[20289]='h00000000;
    rd_cycle[20290] = 1'b0;  wr_cycle[20290] = 1'b0;  addr_rom[20290]='h00000000;  wr_data_rom[20290]='h00000000;
    rd_cycle[20291] = 1'b0;  wr_cycle[20291] = 1'b0;  addr_rom[20291]='h00000000;  wr_data_rom[20291]='h00000000;
    rd_cycle[20292] = 1'b0;  wr_cycle[20292] = 1'b0;  addr_rom[20292]='h00000000;  wr_data_rom[20292]='h00000000;
    rd_cycle[20293] = 1'b0;  wr_cycle[20293] = 1'b0;  addr_rom[20293]='h00000000;  wr_data_rom[20293]='h00000000;
    rd_cycle[20294] = 1'b0;  wr_cycle[20294] = 1'b0;  addr_rom[20294]='h00000000;  wr_data_rom[20294]='h00000000;
    rd_cycle[20295] = 1'b0;  wr_cycle[20295] = 1'b0;  addr_rom[20295]='h00000000;  wr_data_rom[20295]='h00000000;
    rd_cycle[20296] = 1'b0;  wr_cycle[20296] = 1'b0;  addr_rom[20296]='h00000000;  wr_data_rom[20296]='h00000000;
    rd_cycle[20297] = 1'b0;  wr_cycle[20297] = 1'b0;  addr_rom[20297]='h00000000;  wr_data_rom[20297]='h00000000;
    rd_cycle[20298] = 1'b0;  wr_cycle[20298] = 1'b0;  addr_rom[20298]='h00000000;  wr_data_rom[20298]='h00000000;
    rd_cycle[20299] = 1'b0;  wr_cycle[20299] = 1'b0;  addr_rom[20299]='h00000000;  wr_data_rom[20299]='h00000000;
    rd_cycle[20300] = 1'b0;  wr_cycle[20300] = 1'b0;  addr_rom[20300]='h00000000;  wr_data_rom[20300]='h00000000;
    rd_cycle[20301] = 1'b0;  wr_cycle[20301] = 1'b0;  addr_rom[20301]='h00000000;  wr_data_rom[20301]='h00000000;
    rd_cycle[20302] = 1'b0;  wr_cycle[20302] = 1'b0;  addr_rom[20302]='h00000000;  wr_data_rom[20302]='h00000000;
    rd_cycle[20303] = 1'b0;  wr_cycle[20303] = 1'b0;  addr_rom[20303]='h00000000;  wr_data_rom[20303]='h00000000;
    rd_cycle[20304] = 1'b0;  wr_cycle[20304] = 1'b0;  addr_rom[20304]='h00000000;  wr_data_rom[20304]='h00000000;
    rd_cycle[20305] = 1'b0;  wr_cycle[20305] = 1'b0;  addr_rom[20305]='h00000000;  wr_data_rom[20305]='h00000000;
    rd_cycle[20306] = 1'b0;  wr_cycle[20306] = 1'b0;  addr_rom[20306]='h00000000;  wr_data_rom[20306]='h00000000;
    rd_cycle[20307] = 1'b0;  wr_cycle[20307] = 1'b0;  addr_rom[20307]='h00000000;  wr_data_rom[20307]='h00000000;
    rd_cycle[20308] = 1'b0;  wr_cycle[20308] = 1'b0;  addr_rom[20308]='h00000000;  wr_data_rom[20308]='h00000000;
    rd_cycle[20309] = 1'b0;  wr_cycle[20309] = 1'b0;  addr_rom[20309]='h00000000;  wr_data_rom[20309]='h00000000;
    rd_cycle[20310] = 1'b0;  wr_cycle[20310] = 1'b0;  addr_rom[20310]='h00000000;  wr_data_rom[20310]='h00000000;
    rd_cycle[20311] = 1'b0;  wr_cycle[20311] = 1'b0;  addr_rom[20311]='h00000000;  wr_data_rom[20311]='h00000000;
    rd_cycle[20312] = 1'b0;  wr_cycle[20312] = 1'b0;  addr_rom[20312]='h00000000;  wr_data_rom[20312]='h00000000;
    rd_cycle[20313] = 1'b0;  wr_cycle[20313] = 1'b0;  addr_rom[20313]='h00000000;  wr_data_rom[20313]='h00000000;
    rd_cycle[20314] = 1'b0;  wr_cycle[20314] = 1'b0;  addr_rom[20314]='h00000000;  wr_data_rom[20314]='h00000000;
    rd_cycle[20315] = 1'b0;  wr_cycle[20315] = 1'b0;  addr_rom[20315]='h00000000;  wr_data_rom[20315]='h00000000;
    rd_cycle[20316] = 1'b0;  wr_cycle[20316] = 1'b0;  addr_rom[20316]='h00000000;  wr_data_rom[20316]='h00000000;
    rd_cycle[20317] = 1'b0;  wr_cycle[20317] = 1'b0;  addr_rom[20317]='h00000000;  wr_data_rom[20317]='h00000000;
    rd_cycle[20318] = 1'b0;  wr_cycle[20318] = 1'b0;  addr_rom[20318]='h00000000;  wr_data_rom[20318]='h00000000;
    rd_cycle[20319] = 1'b0;  wr_cycle[20319] = 1'b0;  addr_rom[20319]='h00000000;  wr_data_rom[20319]='h00000000;
    rd_cycle[20320] = 1'b0;  wr_cycle[20320] = 1'b0;  addr_rom[20320]='h00000000;  wr_data_rom[20320]='h00000000;
    rd_cycle[20321] = 1'b0;  wr_cycle[20321] = 1'b0;  addr_rom[20321]='h00000000;  wr_data_rom[20321]='h00000000;
    rd_cycle[20322] = 1'b0;  wr_cycle[20322] = 1'b0;  addr_rom[20322]='h00000000;  wr_data_rom[20322]='h00000000;
    rd_cycle[20323] = 1'b0;  wr_cycle[20323] = 1'b0;  addr_rom[20323]='h00000000;  wr_data_rom[20323]='h00000000;
    rd_cycle[20324] = 1'b0;  wr_cycle[20324] = 1'b0;  addr_rom[20324]='h00000000;  wr_data_rom[20324]='h00000000;
    rd_cycle[20325] = 1'b0;  wr_cycle[20325] = 1'b0;  addr_rom[20325]='h00000000;  wr_data_rom[20325]='h00000000;
    rd_cycle[20326] = 1'b0;  wr_cycle[20326] = 1'b0;  addr_rom[20326]='h00000000;  wr_data_rom[20326]='h00000000;
    rd_cycle[20327] = 1'b0;  wr_cycle[20327] = 1'b0;  addr_rom[20327]='h00000000;  wr_data_rom[20327]='h00000000;
    rd_cycle[20328] = 1'b0;  wr_cycle[20328] = 1'b0;  addr_rom[20328]='h00000000;  wr_data_rom[20328]='h00000000;
    rd_cycle[20329] = 1'b0;  wr_cycle[20329] = 1'b0;  addr_rom[20329]='h00000000;  wr_data_rom[20329]='h00000000;
    rd_cycle[20330] = 1'b0;  wr_cycle[20330] = 1'b0;  addr_rom[20330]='h00000000;  wr_data_rom[20330]='h00000000;
    rd_cycle[20331] = 1'b0;  wr_cycle[20331] = 1'b0;  addr_rom[20331]='h00000000;  wr_data_rom[20331]='h00000000;
    rd_cycle[20332] = 1'b0;  wr_cycle[20332] = 1'b0;  addr_rom[20332]='h00000000;  wr_data_rom[20332]='h00000000;
    rd_cycle[20333] = 1'b0;  wr_cycle[20333] = 1'b0;  addr_rom[20333]='h00000000;  wr_data_rom[20333]='h00000000;
    rd_cycle[20334] = 1'b0;  wr_cycle[20334] = 1'b0;  addr_rom[20334]='h00000000;  wr_data_rom[20334]='h00000000;
    rd_cycle[20335] = 1'b0;  wr_cycle[20335] = 1'b0;  addr_rom[20335]='h00000000;  wr_data_rom[20335]='h00000000;
    rd_cycle[20336] = 1'b0;  wr_cycle[20336] = 1'b0;  addr_rom[20336]='h00000000;  wr_data_rom[20336]='h00000000;
    rd_cycle[20337] = 1'b0;  wr_cycle[20337] = 1'b0;  addr_rom[20337]='h00000000;  wr_data_rom[20337]='h00000000;
    rd_cycle[20338] = 1'b0;  wr_cycle[20338] = 1'b0;  addr_rom[20338]='h00000000;  wr_data_rom[20338]='h00000000;
    rd_cycle[20339] = 1'b0;  wr_cycle[20339] = 1'b0;  addr_rom[20339]='h00000000;  wr_data_rom[20339]='h00000000;
    rd_cycle[20340] = 1'b0;  wr_cycle[20340] = 1'b0;  addr_rom[20340]='h00000000;  wr_data_rom[20340]='h00000000;
    rd_cycle[20341] = 1'b0;  wr_cycle[20341] = 1'b0;  addr_rom[20341]='h00000000;  wr_data_rom[20341]='h00000000;
    rd_cycle[20342] = 1'b0;  wr_cycle[20342] = 1'b0;  addr_rom[20342]='h00000000;  wr_data_rom[20342]='h00000000;
    rd_cycle[20343] = 1'b0;  wr_cycle[20343] = 1'b0;  addr_rom[20343]='h00000000;  wr_data_rom[20343]='h00000000;
    rd_cycle[20344] = 1'b0;  wr_cycle[20344] = 1'b0;  addr_rom[20344]='h00000000;  wr_data_rom[20344]='h00000000;
    rd_cycle[20345] = 1'b0;  wr_cycle[20345] = 1'b0;  addr_rom[20345]='h00000000;  wr_data_rom[20345]='h00000000;
    rd_cycle[20346] = 1'b0;  wr_cycle[20346] = 1'b0;  addr_rom[20346]='h00000000;  wr_data_rom[20346]='h00000000;
    rd_cycle[20347] = 1'b0;  wr_cycle[20347] = 1'b0;  addr_rom[20347]='h00000000;  wr_data_rom[20347]='h00000000;
    rd_cycle[20348] = 1'b0;  wr_cycle[20348] = 1'b0;  addr_rom[20348]='h00000000;  wr_data_rom[20348]='h00000000;
    rd_cycle[20349] = 1'b0;  wr_cycle[20349] = 1'b0;  addr_rom[20349]='h00000000;  wr_data_rom[20349]='h00000000;
    rd_cycle[20350] = 1'b0;  wr_cycle[20350] = 1'b0;  addr_rom[20350]='h00000000;  wr_data_rom[20350]='h00000000;
    rd_cycle[20351] = 1'b0;  wr_cycle[20351] = 1'b0;  addr_rom[20351]='h00000000;  wr_data_rom[20351]='h00000000;
    rd_cycle[20352] = 1'b0;  wr_cycle[20352] = 1'b0;  addr_rom[20352]='h00000000;  wr_data_rom[20352]='h00000000;
    rd_cycle[20353] = 1'b0;  wr_cycle[20353] = 1'b0;  addr_rom[20353]='h00000000;  wr_data_rom[20353]='h00000000;
    rd_cycle[20354] = 1'b0;  wr_cycle[20354] = 1'b0;  addr_rom[20354]='h00000000;  wr_data_rom[20354]='h00000000;
    rd_cycle[20355] = 1'b0;  wr_cycle[20355] = 1'b0;  addr_rom[20355]='h00000000;  wr_data_rom[20355]='h00000000;
    rd_cycle[20356] = 1'b0;  wr_cycle[20356] = 1'b0;  addr_rom[20356]='h00000000;  wr_data_rom[20356]='h00000000;
    rd_cycle[20357] = 1'b0;  wr_cycle[20357] = 1'b0;  addr_rom[20357]='h00000000;  wr_data_rom[20357]='h00000000;
    rd_cycle[20358] = 1'b0;  wr_cycle[20358] = 1'b0;  addr_rom[20358]='h00000000;  wr_data_rom[20358]='h00000000;
    rd_cycle[20359] = 1'b0;  wr_cycle[20359] = 1'b0;  addr_rom[20359]='h00000000;  wr_data_rom[20359]='h00000000;
    rd_cycle[20360] = 1'b0;  wr_cycle[20360] = 1'b0;  addr_rom[20360]='h00000000;  wr_data_rom[20360]='h00000000;
    rd_cycle[20361] = 1'b0;  wr_cycle[20361] = 1'b0;  addr_rom[20361]='h00000000;  wr_data_rom[20361]='h00000000;
    rd_cycle[20362] = 1'b0;  wr_cycle[20362] = 1'b0;  addr_rom[20362]='h00000000;  wr_data_rom[20362]='h00000000;
    rd_cycle[20363] = 1'b0;  wr_cycle[20363] = 1'b0;  addr_rom[20363]='h00000000;  wr_data_rom[20363]='h00000000;
    rd_cycle[20364] = 1'b0;  wr_cycle[20364] = 1'b0;  addr_rom[20364]='h00000000;  wr_data_rom[20364]='h00000000;
    rd_cycle[20365] = 1'b0;  wr_cycle[20365] = 1'b0;  addr_rom[20365]='h00000000;  wr_data_rom[20365]='h00000000;
    rd_cycle[20366] = 1'b0;  wr_cycle[20366] = 1'b0;  addr_rom[20366]='h00000000;  wr_data_rom[20366]='h00000000;
    rd_cycle[20367] = 1'b0;  wr_cycle[20367] = 1'b0;  addr_rom[20367]='h00000000;  wr_data_rom[20367]='h00000000;
    rd_cycle[20368] = 1'b0;  wr_cycle[20368] = 1'b0;  addr_rom[20368]='h00000000;  wr_data_rom[20368]='h00000000;
    rd_cycle[20369] = 1'b0;  wr_cycle[20369] = 1'b0;  addr_rom[20369]='h00000000;  wr_data_rom[20369]='h00000000;
    rd_cycle[20370] = 1'b0;  wr_cycle[20370] = 1'b0;  addr_rom[20370]='h00000000;  wr_data_rom[20370]='h00000000;
    rd_cycle[20371] = 1'b0;  wr_cycle[20371] = 1'b0;  addr_rom[20371]='h00000000;  wr_data_rom[20371]='h00000000;
    rd_cycle[20372] = 1'b0;  wr_cycle[20372] = 1'b0;  addr_rom[20372]='h00000000;  wr_data_rom[20372]='h00000000;
    rd_cycle[20373] = 1'b0;  wr_cycle[20373] = 1'b0;  addr_rom[20373]='h00000000;  wr_data_rom[20373]='h00000000;
    rd_cycle[20374] = 1'b0;  wr_cycle[20374] = 1'b0;  addr_rom[20374]='h00000000;  wr_data_rom[20374]='h00000000;
    rd_cycle[20375] = 1'b0;  wr_cycle[20375] = 1'b0;  addr_rom[20375]='h00000000;  wr_data_rom[20375]='h00000000;
    rd_cycle[20376] = 1'b0;  wr_cycle[20376] = 1'b0;  addr_rom[20376]='h00000000;  wr_data_rom[20376]='h00000000;
    rd_cycle[20377] = 1'b0;  wr_cycle[20377] = 1'b0;  addr_rom[20377]='h00000000;  wr_data_rom[20377]='h00000000;
    rd_cycle[20378] = 1'b0;  wr_cycle[20378] = 1'b0;  addr_rom[20378]='h00000000;  wr_data_rom[20378]='h00000000;
    rd_cycle[20379] = 1'b0;  wr_cycle[20379] = 1'b0;  addr_rom[20379]='h00000000;  wr_data_rom[20379]='h00000000;
    rd_cycle[20380] = 1'b0;  wr_cycle[20380] = 1'b0;  addr_rom[20380]='h00000000;  wr_data_rom[20380]='h00000000;
    rd_cycle[20381] = 1'b0;  wr_cycle[20381] = 1'b0;  addr_rom[20381]='h00000000;  wr_data_rom[20381]='h00000000;
    rd_cycle[20382] = 1'b0;  wr_cycle[20382] = 1'b0;  addr_rom[20382]='h00000000;  wr_data_rom[20382]='h00000000;
    rd_cycle[20383] = 1'b0;  wr_cycle[20383] = 1'b0;  addr_rom[20383]='h00000000;  wr_data_rom[20383]='h00000000;
    rd_cycle[20384] = 1'b0;  wr_cycle[20384] = 1'b0;  addr_rom[20384]='h00000000;  wr_data_rom[20384]='h00000000;
    rd_cycle[20385] = 1'b0;  wr_cycle[20385] = 1'b0;  addr_rom[20385]='h00000000;  wr_data_rom[20385]='h00000000;
    rd_cycle[20386] = 1'b0;  wr_cycle[20386] = 1'b0;  addr_rom[20386]='h00000000;  wr_data_rom[20386]='h00000000;
    rd_cycle[20387] = 1'b0;  wr_cycle[20387] = 1'b0;  addr_rom[20387]='h00000000;  wr_data_rom[20387]='h00000000;
    rd_cycle[20388] = 1'b0;  wr_cycle[20388] = 1'b0;  addr_rom[20388]='h00000000;  wr_data_rom[20388]='h00000000;
    rd_cycle[20389] = 1'b0;  wr_cycle[20389] = 1'b0;  addr_rom[20389]='h00000000;  wr_data_rom[20389]='h00000000;
    rd_cycle[20390] = 1'b0;  wr_cycle[20390] = 1'b0;  addr_rom[20390]='h00000000;  wr_data_rom[20390]='h00000000;
    rd_cycle[20391] = 1'b0;  wr_cycle[20391] = 1'b0;  addr_rom[20391]='h00000000;  wr_data_rom[20391]='h00000000;
    rd_cycle[20392] = 1'b0;  wr_cycle[20392] = 1'b0;  addr_rom[20392]='h00000000;  wr_data_rom[20392]='h00000000;
    rd_cycle[20393] = 1'b0;  wr_cycle[20393] = 1'b0;  addr_rom[20393]='h00000000;  wr_data_rom[20393]='h00000000;
    rd_cycle[20394] = 1'b0;  wr_cycle[20394] = 1'b0;  addr_rom[20394]='h00000000;  wr_data_rom[20394]='h00000000;
    rd_cycle[20395] = 1'b0;  wr_cycle[20395] = 1'b0;  addr_rom[20395]='h00000000;  wr_data_rom[20395]='h00000000;
    rd_cycle[20396] = 1'b0;  wr_cycle[20396] = 1'b0;  addr_rom[20396]='h00000000;  wr_data_rom[20396]='h00000000;
    rd_cycle[20397] = 1'b0;  wr_cycle[20397] = 1'b0;  addr_rom[20397]='h00000000;  wr_data_rom[20397]='h00000000;
    rd_cycle[20398] = 1'b0;  wr_cycle[20398] = 1'b0;  addr_rom[20398]='h00000000;  wr_data_rom[20398]='h00000000;
    rd_cycle[20399] = 1'b0;  wr_cycle[20399] = 1'b0;  addr_rom[20399]='h00000000;  wr_data_rom[20399]='h00000000;
    rd_cycle[20400] = 1'b0;  wr_cycle[20400] = 1'b0;  addr_rom[20400]='h00000000;  wr_data_rom[20400]='h00000000;
    rd_cycle[20401] = 1'b0;  wr_cycle[20401] = 1'b0;  addr_rom[20401]='h00000000;  wr_data_rom[20401]='h00000000;
    rd_cycle[20402] = 1'b0;  wr_cycle[20402] = 1'b0;  addr_rom[20402]='h00000000;  wr_data_rom[20402]='h00000000;
    rd_cycle[20403] = 1'b0;  wr_cycle[20403] = 1'b0;  addr_rom[20403]='h00000000;  wr_data_rom[20403]='h00000000;
    rd_cycle[20404] = 1'b0;  wr_cycle[20404] = 1'b0;  addr_rom[20404]='h00000000;  wr_data_rom[20404]='h00000000;
    rd_cycle[20405] = 1'b0;  wr_cycle[20405] = 1'b0;  addr_rom[20405]='h00000000;  wr_data_rom[20405]='h00000000;
    rd_cycle[20406] = 1'b0;  wr_cycle[20406] = 1'b0;  addr_rom[20406]='h00000000;  wr_data_rom[20406]='h00000000;
    rd_cycle[20407] = 1'b0;  wr_cycle[20407] = 1'b0;  addr_rom[20407]='h00000000;  wr_data_rom[20407]='h00000000;
    rd_cycle[20408] = 1'b0;  wr_cycle[20408] = 1'b0;  addr_rom[20408]='h00000000;  wr_data_rom[20408]='h00000000;
    rd_cycle[20409] = 1'b0;  wr_cycle[20409] = 1'b0;  addr_rom[20409]='h00000000;  wr_data_rom[20409]='h00000000;
    rd_cycle[20410] = 1'b0;  wr_cycle[20410] = 1'b0;  addr_rom[20410]='h00000000;  wr_data_rom[20410]='h00000000;
    rd_cycle[20411] = 1'b0;  wr_cycle[20411] = 1'b0;  addr_rom[20411]='h00000000;  wr_data_rom[20411]='h00000000;
    rd_cycle[20412] = 1'b0;  wr_cycle[20412] = 1'b0;  addr_rom[20412]='h00000000;  wr_data_rom[20412]='h00000000;
    rd_cycle[20413] = 1'b0;  wr_cycle[20413] = 1'b0;  addr_rom[20413]='h00000000;  wr_data_rom[20413]='h00000000;
    rd_cycle[20414] = 1'b0;  wr_cycle[20414] = 1'b0;  addr_rom[20414]='h00000000;  wr_data_rom[20414]='h00000000;
    rd_cycle[20415] = 1'b0;  wr_cycle[20415] = 1'b0;  addr_rom[20415]='h00000000;  wr_data_rom[20415]='h00000000;
    rd_cycle[20416] = 1'b0;  wr_cycle[20416] = 1'b0;  addr_rom[20416]='h00000000;  wr_data_rom[20416]='h00000000;
    rd_cycle[20417] = 1'b0;  wr_cycle[20417] = 1'b0;  addr_rom[20417]='h00000000;  wr_data_rom[20417]='h00000000;
    rd_cycle[20418] = 1'b0;  wr_cycle[20418] = 1'b0;  addr_rom[20418]='h00000000;  wr_data_rom[20418]='h00000000;
    rd_cycle[20419] = 1'b0;  wr_cycle[20419] = 1'b0;  addr_rom[20419]='h00000000;  wr_data_rom[20419]='h00000000;
    rd_cycle[20420] = 1'b0;  wr_cycle[20420] = 1'b0;  addr_rom[20420]='h00000000;  wr_data_rom[20420]='h00000000;
    rd_cycle[20421] = 1'b0;  wr_cycle[20421] = 1'b0;  addr_rom[20421]='h00000000;  wr_data_rom[20421]='h00000000;
    rd_cycle[20422] = 1'b0;  wr_cycle[20422] = 1'b0;  addr_rom[20422]='h00000000;  wr_data_rom[20422]='h00000000;
    rd_cycle[20423] = 1'b0;  wr_cycle[20423] = 1'b0;  addr_rom[20423]='h00000000;  wr_data_rom[20423]='h00000000;
    rd_cycle[20424] = 1'b0;  wr_cycle[20424] = 1'b0;  addr_rom[20424]='h00000000;  wr_data_rom[20424]='h00000000;
    rd_cycle[20425] = 1'b0;  wr_cycle[20425] = 1'b0;  addr_rom[20425]='h00000000;  wr_data_rom[20425]='h00000000;
    rd_cycle[20426] = 1'b0;  wr_cycle[20426] = 1'b0;  addr_rom[20426]='h00000000;  wr_data_rom[20426]='h00000000;
    rd_cycle[20427] = 1'b0;  wr_cycle[20427] = 1'b0;  addr_rom[20427]='h00000000;  wr_data_rom[20427]='h00000000;
    rd_cycle[20428] = 1'b0;  wr_cycle[20428] = 1'b0;  addr_rom[20428]='h00000000;  wr_data_rom[20428]='h00000000;
    rd_cycle[20429] = 1'b0;  wr_cycle[20429] = 1'b0;  addr_rom[20429]='h00000000;  wr_data_rom[20429]='h00000000;
    rd_cycle[20430] = 1'b0;  wr_cycle[20430] = 1'b0;  addr_rom[20430]='h00000000;  wr_data_rom[20430]='h00000000;
    rd_cycle[20431] = 1'b0;  wr_cycle[20431] = 1'b0;  addr_rom[20431]='h00000000;  wr_data_rom[20431]='h00000000;
    rd_cycle[20432] = 1'b0;  wr_cycle[20432] = 1'b0;  addr_rom[20432]='h00000000;  wr_data_rom[20432]='h00000000;
    rd_cycle[20433] = 1'b0;  wr_cycle[20433] = 1'b0;  addr_rom[20433]='h00000000;  wr_data_rom[20433]='h00000000;
    rd_cycle[20434] = 1'b0;  wr_cycle[20434] = 1'b0;  addr_rom[20434]='h00000000;  wr_data_rom[20434]='h00000000;
    rd_cycle[20435] = 1'b0;  wr_cycle[20435] = 1'b0;  addr_rom[20435]='h00000000;  wr_data_rom[20435]='h00000000;
    rd_cycle[20436] = 1'b0;  wr_cycle[20436] = 1'b0;  addr_rom[20436]='h00000000;  wr_data_rom[20436]='h00000000;
    rd_cycle[20437] = 1'b0;  wr_cycle[20437] = 1'b0;  addr_rom[20437]='h00000000;  wr_data_rom[20437]='h00000000;
    rd_cycle[20438] = 1'b0;  wr_cycle[20438] = 1'b0;  addr_rom[20438]='h00000000;  wr_data_rom[20438]='h00000000;
    rd_cycle[20439] = 1'b0;  wr_cycle[20439] = 1'b0;  addr_rom[20439]='h00000000;  wr_data_rom[20439]='h00000000;
    rd_cycle[20440] = 1'b0;  wr_cycle[20440] = 1'b0;  addr_rom[20440]='h00000000;  wr_data_rom[20440]='h00000000;
    rd_cycle[20441] = 1'b0;  wr_cycle[20441] = 1'b0;  addr_rom[20441]='h00000000;  wr_data_rom[20441]='h00000000;
    rd_cycle[20442] = 1'b0;  wr_cycle[20442] = 1'b0;  addr_rom[20442]='h00000000;  wr_data_rom[20442]='h00000000;
    rd_cycle[20443] = 1'b0;  wr_cycle[20443] = 1'b0;  addr_rom[20443]='h00000000;  wr_data_rom[20443]='h00000000;
    rd_cycle[20444] = 1'b0;  wr_cycle[20444] = 1'b0;  addr_rom[20444]='h00000000;  wr_data_rom[20444]='h00000000;
    rd_cycle[20445] = 1'b0;  wr_cycle[20445] = 1'b0;  addr_rom[20445]='h00000000;  wr_data_rom[20445]='h00000000;
    rd_cycle[20446] = 1'b0;  wr_cycle[20446] = 1'b0;  addr_rom[20446]='h00000000;  wr_data_rom[20446]='h00000000;
    rd_cycle[20447] = 1'b0;  wr_cycle[20447] = 1'b0;  addr_rom[20447]='h00000000;  wr_data_rom[20447]='h00000000;
    rd_cycle[20448] = 1'b0;  wr_cycle[20448] = 1'b0;  addr_rom[20448]='h00000000;  wr_data_rom[20448]='h00000000;
    rd_cycle[20449] = 1'b0;  wr_cycle[20449] = 1'b0;  addr_rom[20449]='h00000000;  wr_data_rom[20449]='h00000000;
    rd_cycle[20450] = 1'b0;  wr_cycle[20450] = 1'b0;  addr_rom[20450]='h00000000;  wr_data_rom[20450]='h00000000;
    rd_cycle[20451] = 1'b0;  wr_cycle[20451] = 1'b0;  addr_rom[20451]='h00000000;  wr_data_rom[20451]='h00000000;
    rd_cycle[20452] = 1'b0;  wr_cycle[20452] = 1'b0;  addr_rom[20452]='h00000000;  wr_data_rom[20452]='h00000000;
    rd_cycle[20453] = 1'b0;  wr_cycle[20453] = 1'b0;  addr_rom[20453]='h00000000;  wr_data_rom[20453]='h00000000;
    rd_cycle[20454] = 1'b0;  wr_cycle[20454] = 1'b0;  addr_rom[20454]='h00000000;  wr_data_rom[20454]='h00000000;
    rd_cycle[20455] = 1'b0;  wr_cycle[20455] = 1'b0;  addr_rom[20455]='h00000000;  wr_data_rom[20455]='h00000000;
    rd_cycle[20456] = 1'b0;  wr_cycle[20456] = 1'b0;  addr_rom[20456]='h00000000;  wr_data_rom[20456]='h00000000;
    rd_cycle[20457] = 1'b0;  wr_cycle[20457] = 1'b0;  addr_rom[20457]='h00000000;  wr_data_rom[20457]='h00000000;
    rd_cycle[20458] = 1'b0;  wr_cycle[20458] = 1'b0;  addr_rom[20458]='h00000000;  wr_data_rom[20458]='h00000000;
    rd_cycle[20459] = 1'b0;  wr_cycle[20459] = 1'b0;  addr_rom[20459]='h00000000;  wr_data_rom[20459]='h00000000;
    rd_cycle[20460] = 1'b0;  wr_cycle[20460] = 1'b0;  addr_rom[20460]='h00000000;  wr_data_rom[20460]='h00000000;
    rd_cycle[20461] = 1'b0;  wr_cycle[20461] = 1'b0;  addr_rom[20461]='h00000000;  wr_data_rom[20461]='h00000000;
    rd_cycle[20462] = 1'b0;  wr_cycle[20462] = 1'b0;  addr_rom[20462]='h00000000;  wr_data_rom[20462]='h00000000;
    rd_cycle[20463] = 1'b0;  wr_cycle[20463] = 1'b0;  addr_rom[20463]='h00000000;  wr_data_rom[20463]='h00000000;
    rd_cycle[20464] = 1'b0;  wr_cycle[20464] = 1'b0;  addr_rom[20464]='h00000000;  wr_data_rom[20464]='h00000000;
    rd_cycle[20465] = 1'b0;  wr_cycle[20465] = 1'b0;  addr_rom[20465]='h00000000;  wr_data_rom[20465]='h00000000;
    rd_cycle[20466] = 1'b0;  wr_cycle[20466] = 1'b0;  addr_rom[20466]='h00000000;  wr_data_rom[20466]='h00000000;
    rd_cycle[20467] = 1'b0;  wr_cycle[20467] = 1'b0;  addr_rom[20467]='h00000000;  wr_data_rom[20467]='h00000000;
    rd_cycle[20468] = 1'b0;  wr_cycle[20468] = 1'b0;  addr_rom[20468]='h00000000;  wr_data_rom[20468]='h00000000;
    rd_cycle[20469] = 1'b0;  wr_cycle[20469] = 1'b0;  addr_rom[20469]='h00000000;  wr_data_rom[20469]='h00000000;
    rd_cycle[20470] = 1'b0;  wr_cycle[20470] = 1'b0;  addr_rom[20470]='h00000000;  wr_data_rom[20470]='h00000000;
    rd_cycle[20471] = 1'b0;  wr_cycle[20471] = 1'b0;  addr_rom[20471]='h00000000;  wr_data_rom[20471]='h00000000;
    rd_cycle[20472] = 1'b0;  wr_cycle[20472] = 1'b0;  addr_rom[20472]='h00000000;  wr_data_rom[20472]='h00000000;
    rd_cycle[20473] = 1'b0;  wr_cycle[20473] = 1'b0;  addr_rom[20473]='h00000000;  wr_data_rom[20473]='h00000000;
    rd_cycle[20474] = 1'b0;  wr_cycle[20474] = 1'b0;  addr_rom[20474]='h00000000;  wr_data_rom[20474]='h00000000;
    rd_cycle[20475] = 1'b0;  wr_cycle[20475] = 1'b0;  addr_rom[20475]='h00000000;  wr_data_rom[20475]='h00000000;
    rd_cycle[20476] = 1'b0;  wr_cycle[20476] = 1'b0;  addr_rom[20476]='h00000000;  wr_data_rom[20476]='h00000000;
    rd_cycle[20477] = 1'b0;  wr_cycle[20477] = 1'b0;  addr_rom[20477]='h00000000;  wr_data_rom[20477]='h00000000;
    rd_cycle[20478] = 1'b0;  wr_cycle[20478] = 1'b0;  addr_rom[20478]='h00000000;  wr_data_rom[20478]='h00000000;
    rd_cycle[20479] = 1'b0;  wr_cycle[20479] = 1'b0;  addr_rom[20479]='h00000000;  wr_data_rom[20479]='h00000000;
    // 4096 sequence read cycles
    rd_cycle[20480] = 1'b1;  wr_cycle[20480] = 1'b0;  addr_rom[20480]='h00000000;  wr_data_rom[20480]='h00000000;
    rd_cycle[20481] = 1'b1;  wr_cycle[20481] = 1'b0;  addr_rom[20481]='h00000004;  wr_data_rom[20481]='h00000000;
    rd_cycle[20482] = 1'b1;  wr_cycle[20482] = 1'b0;  addr_rom[20482]='h00000008;  wr_data_rom[20482]='h00000000;
    rd_cycle[20483] = 1'b1;  wr_cycle[20483] = 1'b0;  addr_rom[20483]='h0000000c;  wr_data_rom[20483]='h00000000;
    rd_cycle[20484] = 1'b1;  wr_cycle[20484] = 1'b0;  addr_rom[20484]='h00000010;  wr_data_rom[20484]='h00000000;
    rd_cycle[20485] = 1'b1;  wr_cycle[20485] = 1'b0;  addr_rom[20485]='h00000014;  wr_data_rom[20485]='h00000000;
    rd_cycle[20486] = 1'b1;  wr_cycle[20486] = 1'b0;  addr_rom[20486]='h00000018;  wr_data_rom[20486]='h00000000;
    rd_cycle[20487] = 1'b1;  wr_cycle[20487] = 1'b0;  addr_rom[20487]='h0000001c;  wr_data_rom[20487]='h00000000;
    rd_cycle[20488] = 1'b1;  wr_cycle[20488] = 1'b0;  addr_rom[20488]='h00000020;  wr_data_rom[20488]='h00000000;
    rd_cycle[20489] = 1'b1;  wr_cycle[20489] = 1'b0;  addr_rom[20489]='h00000024;  wr_data_rom[20489]='h00000000;
    rd_cycle[20490] = 1'b1;  wr_cycle[20490] = 1'b0;  addr_rom[20490]='h00000028;  wr_data_rom[20490]='h00000000;
    rd_cycle[20491] = 1'b1;  wr_cycle[20491] = 1'b0;  addr_rom[20491]='h0000002c;  wr_data_rom[20491]='h00000000;
    rd_cycle[20492] = 1'b1;  wr_cycle[20492] = 1'b0;  addr_rom[20492]='h00000030;  wr_data_rom[20492]='h00000000;
    rd_cycle[20493] = 1'b1;  wr_cycle[20493] = 1'b0;  addr_rom[20493]='h00000034;  wr_data_rom[20493]='h00000000;
    rd_cycle[20494] = 1'b1;  wr_cycle[20494] = 1'b0;  addr_rom[20494]='h00000038;  wr_data_rom[20494]='h00000000;
    rd_cycle[20495] = 1'b1;  wr_cycle[20495] = 1'b0;  addr_rom[20495]='h0000003c;  wr_data_rom[20495]='h00000000;
    rd_cycle[20496] = 1'b1;  wr_cycle[20496] = 1'b0;  addr_rom[20496]='h00000040;  wr_data_rom[20496]='h00000000;
    rd_cycle[20497] = 1'b1;  wr_cycle[20497] = 1'b0;  addr_rom[20497]='h00000044;  wr_data_rom[20497]='h00000000;
    rd_cycle[20498] = 1'b1;  wr_cycle[20498] = 1'b0;  addr_rom[20498]='h00000048;  wr_data_rom[20498]='h00000000;
    rd_cycle[20499] = 1'b1;  wr_cycle[20499] = 1'b0;  addr_rom[20499]='h0000004c;  wr_data_rom[20499]='h00000000;
    rd_cycle[20500] = 1'b1;  wr_cycle[20500] = 1'b0;  addr_rom[20500]='h00000050;  wr_data_rom[20500]='h00000000;
    rd_cycle[20501] = 1'b1;  wr_cycle[20501] = 1'b0;  addr_rom[20501]='h00000054;  wr_data_rom[20501]='h00000000;
    rd_cycle[20502] = 1'b1;  wr_cycle[20502] = 1'b0;  addr_rom[20502]='h00000058;  wr_data_rom[20502]='h00000000;
    rd_cycle[20503] = 1'b1;  wr_cycle[20503] = 1'b0;  addr_rom[20503]='h0000005c;  wr_data_rom[20503]='h00000000;
    rd_cycle[20504] = 1'b1;  wr_cycle[20504] = 1'b0;  addr_rom[20504]='h00000060;  wr_data_rom[20504]='h00000000;
    rd_cycle[20505] = 1'b1;  wr_cycle[20505] = 1'b0;  addr_rom[20505]='h00000064;  wr_data_rom[20505]='h00000000;
    rd_cycle[20506] = 1'b1;  wr_cycle[20506] = 1'b0;  addr_rom[20506]='h00000068;  wr_data_rom[20506]='h00000000;
    rd_cycle[20507] = 1'b1;  wr_cycle[20507] = 1'b0;  addr_rom[20507]='h0000006c;  wr_data_rom[20507]='h00000000;
    rd_cycle[20508] = 1'b1;  wr_cycle[20508] = 1'b0;  addr_rom[20508]='h00000070;  wr_data_rom[20508]='h00000000;
    rd_cycle[20509] = 1'b1;  wr_cycle[20509] = 1'b0;  addr_rom[20509]='h00000074;  wr_data_rom[20509]='h00000000;
    rd_cycle[20510] = 1'b1;  wr_cycle[20510] = 1'b0;  addr_rom[20510]='h00000078;  wr_data_rom[20510]='h00000000;
    rd_cycle[20511] = 1'b1;  wr_cycle[20511] = 1'b0;  addr_rom[20511]='h0000007c;  wr_data_rom[20511]='h00000000;
    rd_cycle[20512] = 1'b1;  wr_cycle[20512] = 1'b0;  addr_rom[20512]='h00000080;  wr_data_rom[20512]='h00000000;
    rd_cycle[20513] = 1'b1;  wr_cycle[20513] = 1'b0;  addr_rom[20513]='h00000084;  wr_data_rom[20513]='h00000000;
    rd_cycle[20514] = 1'b1;  wr_cycle[20514] = 1'b0;  addr_rom[20514]='h00000088;  wr_data_rom[20514]='h00000000;
    rd_cycle[20515] = 1'b1;  wr_cycle[20515] = 1'b0;  addr_rom[20515]='h0000008c;  wr_data_rom[20515]='h00000000;
    rd_cycle[20516] = 1'b1;  wr_cycle[20516] = 1'b0;  addr_rom[20516]='h00000090;  wr_data_rom[20516]='h00000000;
    rd_cycle[20517] = 1'b1;  wr_cycle[20517] = 1'b0;  addr_rom[20517]='h00000094;  wr_data_rom[20517]='h00000000;
    rd_cycle[20518] = 1'b1;  wr_cycle[20518] = 1'b0;  addr_rom[20518]='h00000098;  wr_data_rom[20518]='h00000000;
    rd_cycle[20519] = 1'b1;  wr_cycle[20519] = 1'b0;  addr_rom[20519]='h0000009c;  wr_data_rom[20519]='h00000000;
    rd_cycle[20520] = 1'b1;  wr_cycle[20520] = 1'b0;  addr_rom[20520]='h000000a0;  wr_data_rom[20520]='h00000000;
    rd_cycle[20521] = 1'b1;  wr_cycle[20521] = 1'b0;  addr_rom[20521]='h000000a4;  wr_data_rom[20521]='h00000000;
    rd_cycle[20522] = 1'b1;  wr_cycle[20522] = 1'b0;  addr_rom[20522]='h000000a8;  wr_data_rom[20522]='h00000000;
    rd_cycle[20523] = 1'b1;  wr_cycle[20523] = 1'b0;  addr_rom[20523]='h000000ac;  wr_data_rom[20523]='h00000000;
    rd_cycle[20524] = 1'b1;  wr_cycle[20524] = 1'b0;  addr_rom[20524]='h000000b0;  wr_data_rom[20524]='h00000000;
    rd_cycle[20525] = 1'b1;  wr_cycle[20525] = 1'b0;  addr_rom[20525]='h000000b4;  wr_data_rom[20525]='h00000000;
    rd_cycle[20526] = 1'b1;  wr_cycle[20526] = 1'b0;  addr_rom[20526]='h000000b8;  wr_data_rom[20526]='h00000000;
    rd_cycle[20527] = 1'b1;  wr_cycle[20527] = 1'b0;  addr_rom[20527]='h000000bc;  wr_data_rom[20527]='h00000000;
    rd_cycle[20528] = 1'b1;  wr_cycle[20528] = 1'b0;  addr_rom[20528]='h000000c0;  wr_data_rom[20528]='h00000000;
    rd_cycle[20529] = 1'b1;  wr_cycle[20529] = 1'b0;  addr_rom[20529]='h000000c4;  wr_data_rom[20529]='h00000000;
    rd_cycle[20530] = 1'b1;  wr_cycle[20530] = 1'b0;  addr_rom[20530]='h000000c8;  wr_data_rom[20530]='h00000000;
    rd_cycle[20531] = 1'b1;  wr_cycle[20531] = 1'b0;  addr_rom[20531]='h000000cc;  wr_data_rom[20531]='h00000000;
    rd_cycle[20532] = 1'b1;  wr_cycle[20532] = 1'b0;  addr_rom[20532]='h000000d0;  wr_data_rom[20532]='h00000000;
    rd_cycle[20533] = 1'b1;  wr_cycle[20533] = 1'b0;  addr_rom[20533]='h000000d4;  wr_data_rom[20533]='h00000000;
    rd_cycle[20534] = 1'b1;  wr_cycle[20534] = 1'b0;  addr_rom[20534]='h000000d8;  wr_data_rom[20534]='h00000000;
    rd_cycle[20535] = 1'b1;  wr_cycle[20535] = 1'b0;  addr_rom[20535]='h000000dc;  wr_data_rom[20535]='h00000000;
    rd_cycle[20536] = 1'b1;  wr_cycle[20536] = 1'b0;  addr_rom[20536]='h000000e0;  wr_data_rom[20536]='h00000000;
    rd_cycle[20537] = 1'b1;  wr_cycle[20537] = 1'b0;  addr_rom[20537]='h000000e4;  wr_data_rom[20537]='h00000000;
    rd_cycle[20538] = 1'b1;  wr_cycle[20538] = 1'b0;  addr_rom[20538]='h000000e8;  wr_data_rom[20538]='h00000000;
    rd_cycle[20539] = 1'b1;  wr_cycle[20539] = 1'b0;  addr_rom[20539]='h000000ec;  wr_data_rom[20539]='h00000000;
    rd_cycle[20540] = 1'b1;  wr_cycle[20540] = 1'b0;  addr_rom[20540]='h000000f0;  wr_data_rom[20540]='h00000000;
    rd_cycle[20541] = 1'b1;  wr_cycle[20541] = 1'b0;  addr_rom[20541]='h000000f4;  wr_data_rom[20541]='h00000000;
    rd_cycle[20542] = 1'b1;  wr_cycle[20542] = 1'b0;  addr_rom[20542]='h000000f8;  wr_data_rom[20542]='h00000000;
    rd_cycle[20543] = 1'b1;  wr_cycle[20543] = 1'b0;  addr_rom[20543]='h000000fc;  wr_data_rom[20543]='h00000000;
    rd_cycle[20544] = 1'b1;  wr_cycle[20544] = 1'b0;  addr_rom[20544]='h00000100;  wr_data_rom[20544]='h00000000;
    rd_cycle[20545] = 1'b1;  wr_cycle[20545] = 1'b0;  addr_rom[20545]='h00000104;  wr_data_rom[20545]='h00000000;
    rd_cycle[20546] = 1'b1;  wr_cycle[20546] = 1'b0;  addr_rom[20546]='h00000108;  wr_data_rom[20546]='h00000000;
    rd_cycle[20547] = 1'b1;  wr_cycle[20547] = 1'b0;  addr_rom[20547]='h0000010c;  wr_data_rom[20547]='h00000000;
    rd_cycle[20548] = 1'b1;  wr_cycle[20548] = 1'b0;  addr_rom[20548]='h00000110;  wr_data_rom[20548]='h00000000;
    rd_cycle[20549] = 1'b1;  wr_cycle[20549] = 1'b0;  addr_rom[20549]='h00000114;  wr_data_rom[20549]='h00000000;
    rd_cycle[20550] = 1'b1;  wr_cycle[20550] = 1'b0;  addr_rom[20550]='h00000118;  wr_data_rom[20550]='h00000000;
    rd_cycle[20551] = 1'b1;  wr_cycle[20551] = 1'b0;  addr_rom[20551]='h0000011c;  wr_data_rom[20551]='h00000000;
    rd_cycle[20552] = 1'b1;  wr_cycle[20552] = 1'b0;  addr_rom[20552]='h00000120;  wr_data_rom[20552]='h00000000;
    rd_cycle[20553] = 1'b1;  wr_cycle[20553] = 1'b0;  addr_rom[20553]='h00000124;  wr_data_rom[20553]='h00000000;
    rd_cycle[20554] = 1'b1;  wr_cycle[20554] = 1'b0;  addr_rom[20554]='h00000128;  wr_data_rom[20554]='h00000000;
    rd_cycle[20555] = 1'b1;  wr_cycle[20555] = 1'b0;  addr_rom[20555]='h0000012c;  wr_data_rom[20555]='h00000000;
    rd_cycle[20556] = 1'b1;  wr_cycle[20556] = 1'b0;  addr_rom[20556]='h00000130;  wr_data_rom[20556]='h00000000;
    rd_cycle[20557] = 1'b1;  wr_cycle[20557] = 1'b0;  addr_rom[20557]='h00000134;  wr_data_rom[20557]='h00000000;
    rd_cycle[20558] = 1'b1;  wr_cycle[20558] = 1'b0;  addr_rom[20558]='h00000138;  wr_data_rom[20558]='h00000000;
    rd_cycle[20559] = 1'b1;  wr_cycle[20559] = 1'b0;  addr_rom[20559]='h0000013c;  wr_data_rom[20559]='h00000000;
    rd_cycle[20560] = 1'b1;  wr_cycle[20560] = 1'b0;  addr_rom[20560]='h00000140;  wr_data_rom[20560]='h00000000;
    rd_cycle[20561] = 1'b1;  wr_cycle[20561] = 1'b0;  addr_rom[20561]='h00000144;  wr_data_rom[20561]='h00000000;
    rd_cycle[20562] = 1'b1;  wr_cycle[20562] = 1'b0;  addr_rom[20562]='h00000148;  wr_data_rom[20562]='h00000000;
    rd_cycle[20563] = 1'b1;  wr_cycle[20563] = 1'b0;  addr_rom[20563]='h0000014c;  wr_data_rom[20563]='h00000000;
    rd_cycle[20564] = 1'b1;  wr_cycle[20564] = 1'b0;  addr_rom[20564]='h00000150;  wr_data_rom[20564]='h00000000;
    rd_cycle[20565] = 1'b1;  wr_cycle[20565] = 1'b0;  addr_rom[20565]='h00000154;  wr_data_rom[20565]='h00000000;
    rd_cycle[20566] = 1'b1;  wr_cycle[20566] = 1'b0;  addr_rom[20566]='h00000158;  wr_data_rom[20566]='h00000000;
    rd_cycle[20567] = 1'b1;  wr_cycle[20567] = 1'b0;  addr_rom[20567]='h0000015c;  wr_data_rom[20567]='h00000000;
    rd_cycle[20568] = 1'b1;  wr_cycle[20568] = 1'b0;  addr_rom[20568]='h00000160;  wr_data_rom[20568]='h00000000;
    rd_cycle[20569] = 1'b1;  wr_cycle[20569] = 1'b0;  addr_rom[20569]='h00000164;  wr_data_rom[20569]='h00000000;
    rd_cycle[20570] = 1'b1;  wr_cycle[20570] = 1'b0;  addr_rom[20570]='h00000168;  wr_data_rom[20570]='h00000000;
    rd_cycle[20571] = 1'b1;  wr_cycle[20571] = 1'b0;  addr_rom[20571]='h0000016c;  wr_data_rom[20571]='h00000000;
    rd_cycle[20572] = 1'b1;  wr_cycle[20572] = 1'b0;  addr_rom[20572]='h00000170;  wr_data_rom[20572]='h00000000;
    rd_cycle[20573] = 1'b1;  wr_cycle[20573] = 1'b0;  addr_rom[20573]='h00000174;  wr_data_rom[20573]='h00000000;
    rd_cycle[20574] = 1'b1;  wr_cycle[20574] = 1'b0;  addr_rom[20574]='h00000178;  wr_data_rom[20574]='h00000000;
    rd_cycle[20575] = 1'b1;  wr_cycle[20575] = 1'b0;  addr_rom[20575]='h0000017c;  wr_data_rom[20575]='h00000000;
    rd_cycle[20576] = 1'b1;  wr_cycle[20576] = 1'b0;  addr_rom[20576]='h00000180;  wr_data_rom[20576]='h00000000;
    rd_cycle[20577] = 1'b1;  wr_cycle[20577] = 1'b0;  addr_rom[20577]='h00000184;  wr_data_rom[20577]='h00000000;
    rd_cycle[20578] = 1'b1;  wr_cycle[20578] = 1'b0;  addr_rom[20578]='h00000188;  wr_data_rom[20578]='h00000000;
    rd_cycle[20579] = 1'b1;  wr_cycle[20579] = 1'b0;  addr_rom[20579]='h0000018c;  wr_data_rom[20579]='h00000000;
    rd_cycle[20580] = 1'b1;  wr_cycle[20580] = 1'b0;  addr_rom[20580]='h00000190;  wr_data_rom[20580]='h00000000;
    rd_cycle[20581] = 1'b1;  wr_cycle[20581] = 1'b0;  addr_rom[20581]='h00000194;  wr_data_rom[20581]='h00000000;
    rd_cycle[20582] = 1'b1;  wr_cycle[20582] = 1'b0;  addr_rom[20582]='h00000198;  wr_data_rom[20582]='h00000000;
    rd_cycle[20583] = 1'b1;  wr_cycle[20583] = 1'b0;  addr_rom[20583]='h0000019c;  wr_data_rom[20583]='h00000000;
    rd_cycle[20584] = 1'b1;  wr_cycle[20584] = 1'b0;  addr_rom[20584]='h000001a0;  wr_data_rom[20584]='h00000000;
    rd_cycle[20585] = 1'b1;  wr_cycle[20585] = 1'b0;  addr_rom[20585]='h000001a4;  wr_data_rom[20585]='h00000000;
    rd_cycle[20586] = 1'b1;  wr_cycle[20586] = 1'b0;  addr_rom[20586]='h000001a8;  wr_data_rom[20586]='h00000000;
    rd_cycle[20587] = 1'b1;  wr_cycle[20587] = 1'b0;  addr_rom[20587]='h000001ac;  wr_data_rom[20587]='h00000000;
    rd_cycle[20588] = 1'b1;  wr_cycle[20588] = 1'b0;  addr_rom[20588]='h000001b0;  wr_data_rom[20588]='h00000000;
    rd_cycle[20589] = 1'b1;  wr_cycle[20589] = 1'b0;  addr_rom[20589]='h000001b4;  wr_data_rom[20589]='h00000000;
    rd_cycle[20590] = 1'b1;  wr_cycle[20590] = 1'b0;  addr_rom[20590]='h000001b8;  wr_data_rom[20590]='h00000000;
    rd_cycle[20591] = 1'b1;  wr_cycle[20591] = 1'b0;  addr_rom[20591]='h000001bc;  wr_data_rom[20591]='h00000000;
    rd_cycle[20592] = 1'b1;  wr_cycle[20592] = 1'b0;  addr_rom[20592]='h000001c0;  wr_data_rom[20592]='h00000000;
    rd_cycle[20593] = 1'b1;  wr_cycle[20593] = 1'b0;  addr_rom[20593]='h000001c4;  wr_data_rom[20593]='h00000000;
    rd_cycle[20594] = 1'b1;  wr_cycle[20594] = 1'b0;  addr_rom[20594]='h000001c8;  wr_data_rom[20594]='h00000000;
    rd_cycle[20595] = 1'b1;  wr_cycle[20595] = 1'b0;  addr_rom[20595]='h000001cc;  wr_data_rom[20595]='h00000000;
    rd_cycle[20596] = 1'b1;  wr_cycle[20596] = 1'b0;  addr_rom[20596]='h000001d0;  wr_data_rom[20596]='h00000000;
    rd_cycle[20597] = 1'b1;  wr_cycle[20597] = 1'b0;  addr_rom[20597]='h000001d4;  wr_data_rom[20597]='h00000000;
    rd_cycle[20598] = 1'b1;  wr_cycle[20598] = 1'b0;  addr_rom[20598]='h000001d8;  wr_data_rom[20598]='h00000000;
    rd_cycle[20599] = 1'b1;  wr_cycle[20599] = 1'b0;  addr_rom[20599]='h000001dc;  wr_data_rom[20599]='h00000000;
    rd_cycle[20600] = 1'b1;  wr_cycle[20600] = 1'b0;  addr_rom[20600]='h000001e0;  wr_data_rom[20600]='h00000000;
    rd_cycle[20601] = 1'b1;  wr_cycle[20601] = 1'b0;  addr_rom[20601]='h000001e4;  wr_data_rom[20601]='h00000000;
    rd_cycle[20602] = 1'b1;  wr_cycle[20602] = 1'b0;  addr_rom[20602]='h000001e8;  wr_data_rom[20602]='h00000000;
    rd_cycle[20603] = 1'b1;  wr_cycle[20603] = 1'b0;  addr_rom[20603]='h000001ec;  wr_data_rom[20603]='h00000000;
    rd_cycle[20604] = 1'b1;  wr_cycle[20604] = 1'b0;  addr_rom[20604]='h000001f0;  wr_data_rom[20604]='h00000000;
    rd_cycle[20605] = 1'b1;  wr_cycle[20605] = 1'b0;  addr_rom[20605]='h000001f4;  wr_data_rom[20605]='h00000000;
    rd_cycle[20606] = 1'b1;  wr_cycle[20606] = 1'b0;  addr_rom[20606]='h000001f8;  wr_data_rom[20606]='h00000000;
    rd_cycle[20607] = 1'b1;  wr_cycle[20607] = 1'b0;  addr_rom[20607]='h000001fc;  wr_data_rom[20607]='h00000000;
    rd_cycle[20608] = 1'b1;  wr_cycle[20608] = 1'b0;  addr_rom[20608]='h00000200;  wr_data_rom[20608]='h00000000;
    rd_cycle[20609] = 1'b1;  wr_cycle[20609] = 1'b0;  addr_rom[20609]='h00000204;  wr_data_rom[20609]='h00000000;
    rd_cycle[20610] = 1'b1;  wr_cycle[20610] = 1'b0;  addr_rom[20610]='h00000208;  wr_data_rom[20610]='h00000000;
    rd_cycle[20611] = 1'b1;  wr_cycle[20611] = 1'b0;  addr_rom[20611]='h0000020c;  wr_data_rom[20611]='h00000000;
    rd_cycle[20612] = 1'b1;  wr_cycle[20612] = 1'b0;  addr_rom[20612]='h00000210;  wr_data_rom[20612]='h00000000;
    rd_cycle[20613] = 1'b1;  wr_cycle[20613] = 1'b0;  addr_rom[20613]='h00000214;  wr_data_rom[20613]='h00000000;
    rd_cycle[20614] = 1'b1;  wr_cycle[20614] = 1'b0;  addr_rom[20614]='h00000218;  wr_data_rom[20614]='h00000000;
    rd_cycle[20615] = 1'b1;  wr_cycle[20615] = 1'b0;  addr_rom[20615]='h0000021c;  wr_data_rom[20615]='h00000000;
    rd_cycle[20616] = 1'b1;  wr_cycle[20616] = 1'b0;  addr_rom[20616]='h00000220;  wr_data_rom[20616]='h00000000;
    rd_cycle[20617] = 1'b1;  wr_cycle[20617] = 1'b0;  addr_rom[20617]='h00000224;  wr_data_rom[20617]='h00000000;
    rd_cycle[20618] = 1'b1;  wr_cycle[20618] = 1'b0;  addr_rom[20618]='h00000228;  wr_data_rom[20618]='h00000000;
    rd_cycle[20619] = 1'b1;  wr_cycle[20619] = 1'b0;  addr_rom[20619]='h0000022c;  wr_data_rom[20619]='h00000000;
    rd_cycle[20620] = 1'b1;  wr_cycle[20620] = 1'b0;  addr_rom[20620]='h00000230;  wr_data_rom[20620]='h00000000;
    rd_cycle[20621] = 1'b1;  wr_cycle[20621] = 1'b0;  addr_rom[20621]='h00000234;  wr_data_rom[20621]='h00000000;
    rd_cycle[20622] = 1'b1;  wr_cycle[20622] = 1'b0;  addr_rom[20622]='h00000238;  wr_data_rom[20622]='h00000000;
    rd_cycle[20623] = 1'b1;  wr_cycle[20623] = 1'b0;  addr_rom[20623]='h0000023c;  wr_data_rom[20623]='h00000000;
    rd_cycle[20624] = 1'b1;  wr_cycle[20624] = 1'b0;  addr_rom[20624]='h00000240;  wr_data_rom[20624]='h00000000;
    rd_cycle[20625] = 1'b1;  wr_cycle[20625] = 1'b0;  addr_rom[20625]='h00000244;  wr_data_rom[20625]='h00000000;
    rd_cycle[20626] = 1'b1;  wr_cycle[20626] = 1'b0;  addr_rom[20626]='h00000248;  wr_data_rom[20626]='h00000000;
    rd_cycle[20627] = 1'b1;  wr_cycle[20627] = 1'b0;  addr_rom[20627]='h0000024c;  wr_data_rom[20627]='h00000000;
    rd_cycle[20628] = 1'b1;  wr_cycle[20628] = 1'b0;  addr_rom[20628]='h00000250;  wr_data_rom[20628]='h00000000;
    rd_cycle[20629] = 1'b1;  wr_cycle[20629] = 1'b0;  addr_rom[20629]='h00000254;  wr_data_rom[20629]='h00000000;
    rd_cycle[20630] = 1'b1;  wr_cycle[20630] = 1'b0;  addr_rom[20630]='h00000258;  wr_data_rom[20630]='h00000000;
    rd_cycle[20631] = 1'b1;  wr_cycle[20631] = 1'b0;  addr_rom[20631]='h0000025c;  wr_data_rom[20631]='h00000000;
    rd_cycle[20632] = 1'b1;  wr_cycle[20632] = 1'b0;  addr_rom[20632]='h00000260;  wr_data_rom[20632]='h00000000;
    rd_cycle[20633] = 1'b1;  wr_cycle[20633] = 1'b0;  addr_rom[20633]='h00000264;  wr_data_rom[20633]='h00000000;
    rd_cycle[20634] = 1'b1;  wr_cycle[20634] = 1'b0;  addr_rom[20634]='h00000268;  wr_data_rom[20634]='h00000000;
    rd_cycle[20635] = 1'b1;  wr_cycle[20635] = 1'b0;  addr_rom[20635]='h0000026c;  wr_data_rom[20635]='h00000000;
    rd_cycle[20636] = 1'b1;  wr_cycle[20636] = 1'b0;  addr_rom[20636]='h00000270;  wr_data_rom[20636]='h00000000;
    rd_cycle[20637] = 1'b1;  wr_cycle[20637] = 1'b0;  addr_rom[20637]='h00000274;  wr_data_rom[20637]='h00000000;
    rd_cycle[20638] = 1'b1;  wr_cycle[20638] = 1'b0;  addr_rom[20638]='h00000278;  wr_data_rom[20638]='h00000000;
    rd_cycle[20639] = 1'b1;  wr_cycle[20639] = 1'b0;  addr_rom[20639]='h0000027c;  wr_data_rom[20639]='h00000000;
    rd_cycle[20640] = 1'b1;  wr_cycle[20640] = 1'b0;  addr_rom[20640]='h00000280;  wr_data_rom[20640]='h00000000;
    rd_cycle[20641] = 1'b1;  wr_cycle[20641] = 1'b0;  addr_rom[20641]='h00000284;  wr_data_rom[20641]='h00000000;
    rd_cycle[20642] = 1'b1;  wr_cycle[20642] = 1'b0;  addr_rom[20642]='h00000288;  wr_data_rom[20642]='h00000000;
    rd_cycle[20643] = 1'b1;  wr_cycle[20643] = 1'b0;  addr_rom[20643]='h0000028c;  wr_data_rom[20643]='h00000000;
    rd_cycle[20644] = 1'b1;  wr_cycle[20644] = 1'b0;  addr_rom[20644]='h00000290;  wr_data_rom[20644]='h00000000;
    rd_cycle[20645] = 1'b1;  wr_cycle[20645] = 1'b0;  addr_rom[20645]='h00000294;  wr_data_rom[20645]='h00000000;
    rd_cycle[20646] = 1'b1;  wr_cycle[20646] = 1'b0;  addr_rom[20646]='h00000298;  wr_data_rom[20646]='h00000000;
    rd_cycle[20647] = 1'b1;  wr_cycle[20647] = 1'b0;  addr_rom[20647]='h0000029c;  wr_data_rom[20647]='h00000000;
    rd_cycle[20648] = 1'b1;  wr_cycle[20648] = 1'b0;  addr_rom[20648]='h000002a0;  wr_data_rom[20648]='h00000000;
    rd_cycle[20649] = 1'b1;  wr_cycle[20649] = 1'b0;  addr_rom[20649]='h000002a4;  wr_data_rom[20649]='h00000000;
    rd_cycle[20650] = 1'b1;  wr_cycle[20650] = 1'b0;  addr_rom[20650]='h000002a8;  wr_data_rom[20650]='h00000000;
    rd_cycle[20651] = 1'b1;  wr_cycle[20651] = 1'b0;  addr_rom[20651]='h000002ac;  wr_data_rom[20651]='h00000000;
    rd_cycle[20652] = 1'b1;  wr_cycle[20652] = 1'b0;  addr_rom[20652]='h000002b0;  wr_data_rom[20652]='h00000000;
    rd_cycle[20653] = 1'b1;  wr_cycle[20653] = 1'b0;  addr_rom[20653]='h000002b4;  wr_data_rom[20653]='h00000000;
    rd_cycle[20654] = 1'b1;  wr_cycle[20654] = 1'b0;  addr_rom[20654]='h000002b8;  wr_data_rom[20654]='h00000000;
    rd_cycle[20655] = 1'b1;  wr_cycle[20655] = 1'b0;  addr_rom[20655]='h000002bc;  wr_data_rom[20655]='h00000000;
    rd_cycle[20656] = 1'b1;  wr_cycle[20656] = 1'b0;  addr_rom[20656]='h000002c0;  wr_data_rom[20656]='h00000000;
    rd_cycle[20657] = 1'b1;  wr_cycle[20657] = 1'b0;  addr_rom[20657]='h000002c4;  wr_data_rom[20657]='h00000000;
    rd_cycle[20658] = 1'b1;  wr_cycle[20658] = 1'b0;  addr_rom[20658]='h000002c8;  wr_data_rom[20658]='h00000000;
    rd_cycle[20659] = 1'b1;  wr_cycle[20659] = 1'b0;  addr_rom[20659]='h000002cc;  wr_data_rom[20659]='h00000000;
    rd_cycle[20660] = 1'b1;  wr_cycle[20660] = 1'b0;  addr_rom[20660]='h000002d0;  wr_data_rom[20660]='h00000000;
    rd_cycle[20661] = 1'b1;  wr_cycle[20661] = 1'b0;  addr_rom[20661]='h000002d4;  wr_data_rom[20661]='h00000000;
    rd_cycle[20662] = 1'b1;  wr_cycle[20662] = 1'b0;  addr_rom[20662]='h000002d8;  wr_data_rom[20662]='h00000000;
    rd_cycle[20663] = 1'b1;  wr_cycle[20663] = 1'b0;  addr_rom[20663]='h000002dc;  wr_data_rom[20663]='h00000000;
    rd_cycle[20664] = 1'b1;  wr_cycle[20664] = 1'b0;  addr_rom[20664]='h000002e0;  wr_data_rom[20664]='h00000000;
    rd_cycle[20665] = 1'b1;  wr_cycle[20665] = 1'b0;  addr_rom[20665]='h000002e4;  wr_data_rom[20665]='h00000000;
    rd_cycle[20666] = 1'b1;  wr_cycle[20666] = 1'b0;  addr_rom[20666]='h000002e8;  wr_data_rom[20666]='h00000000;
    rd_cycle[20667] = 1'b1;  wr_cycle[20667] = 1'b0;  addr_rom[20667]='h000002ec;  wr_data_rom[20667]='h00000000;
    rd_cycle[20668] = 1'b1;  wr_cycle[20668] = 1'b0;  addr_rom[20668]='h000002f0;  wr_data_rom[20668]='h00000000;
    rd_cycle[20669] = 1'b1;  wr_cycle[20669] = 1'b0;  addr_rom[20669]='h000002f4;  wr_data_rom[20669]='h00000000;
    rd_cycle[20670] = 1'b1;  wr_cycle[20670] = 1'b0;  addr_rom[20670]='h000002f8;  wr_data_rom[20670]='h00000000;
    rd_cycle[20671] = 1'b1;  wr_cycle[20671] = 1'b0;  addr_rom[20671]='h000002fc;  wr_data_rom[20671]='h00000000;
    rd_cycle[20672] = 1'b1;  wr_cycle[20672] = 1'b0;  addr_rom[20672]='h00000300;  wr_data_rom[20672]='h00000000;
    rd_cycle[20673] = 1'b1;  wr_cycle[20673] = 1'b0;  addr_rom[20673]='h00000304;  wr_data_rom[20673]='h00000000;
    rd_cycle[20674] = 1'b1;  wr_cycle[20674] = 1'b0;  addr_rom[20674]='h00000308;  wr_data_rom[20674]='h00000000;
    rd_cycle[20675] = 1'b1;  wr_cycle[20675] = 1'b0;  addr_rom[20675]='h0000030c;  wr_data_rom[20675]='h00000000;
    rd_cycle[20676] = 1'b1;  wr_cycle[20676] = 1'b0;  addr_rom[20676]='h00000310;  wr_data_rom[20676]='h00000000;
    rd_cycle[20677] = 1'b1;  wr_cycle[20677] = 1'b0;  addr_rom[20677]='h00000314;  wr_data_rom[20677]='h00000000;
    rd_cycle[20678] = 1'b1;  wr_cycle[20678] = 1'b0;  addr_rom[20678]='h00000318;  wr_data_rom[20678]='h00000000;
    rd_cycle[20679] = 1'b1;  wr_cycle[20679] = 1'b0;  addr_rom[20679]='h0000031c;  wr_data_rom[20679]='h00000000;
    rd_cycle[20680] = 1'b1;  wr_cycle[20680] = 1'b0;  addr_rom[20680]='h00000320;  wr_data_rom[20680]='h00000000;
    rd_cycle[20681] = 1'b1;  wr_cycle[20681] = 1'b0;  addr_rom[20681]='h00000324;  wr_data_rom[20681]='h00000000;
    rd_cycle[20682] = 1'b1;  wr_cycle[20682] = 1'b0;  addr_rom[20682]='h00000328;  wr_data_rom[20682]='h00000000;
    rd_cycle[20683] = 1'b1;  wr_cycle[20683] = 1'b0;  addr_rom[20683]='h0000032c;  wr_data_rom[20683]='h00000000;
    rd_cycle[20684] = 1'b1;  wr_cycle[20684] = 1'b0;  addr_rom[20684]='h00000330;  wr_data_rom[20684]='h00000000;
    rd_cycle[20685] = 1'b1;  wr_cycle[20685] = 1'b0;  addr_rom[20685]='h00000334;  wr_data_rom[20685]='h00000000;
    rd_cycle[20686] = 1'b1;  wr_cycle[20686] = 1'b0;  addr_rom[20686]='h00000338;  wr_data_rom[20686]='h00000000;
    rd_cycle[20687] = 1'b1;  wr_cycle[20687] = 1'b0;  addr_rom[20687]='h0000033c;  wr_data_rom[20687]='h00000000;
    rd_cycle[20688] = 1'b1;  wr_cycle[20688] = 1'b0;  addr_rom[20688]='h00000340;  wr_data_rom[20688]='h00000000;
    rd_cycle[20689] = 1'b1;  wr_cycle[20689] = 1'b0;  addr_rom[20689]='h00000344;  wr_data_rom[20689]='h00000000;
    rd_cycle[20690] = 1'b1;  wr_cycle[20690] = 1'b0;  addr_rom[20690]='h00000348;  wr_data_rom[20690]='h00000000;
    rd_cycle[20691] = 1'b1;  wr_cycle[20691] = 1'b0;  addr_rom[20691]='h0000034c;  wr_data_rom[20691]='h00000000;
    rd_cycle[20692] = 1'b1;  wr_cycle[20692] = 1'b0;  addr_rom[20692]='h00000350;  wr_data_rom[20692]='h00000000;
    rd_cycle[20693] = 1'b1;  wr_cycle[20693] = 1'b0;  addr_rom[20693]='h00000354;  wr_data_rom[20693]='h00000000;
    rd_cycle[20694] = 1'b1;  wr_cycle[20694] = 1'b0;  addr_rom[20694]='h00000358;  wr_data_rom[20694]='h00000000;
    rd_cycle[20695] = 1'b1;  wr_cycle[20695] = 1'b0;  addr_rom[20695]='h0000035c;  wr_data_rom[20695]='h00000000;
    rd_cycle[20696] = 1'b1;  wr_cycle[20696] = 1'b0;  addr_rom[20696]='h00000360;  wr_data_rom[20696]='h00000000;
    rd_cycle[20697] = 1'b1;  wr_cycle[20697] = 1'b0;  addr_rom[20697]='h00000364;  wr_data_rom[20697]='h00000000;
    rd_cycle[20698] = 1'b1;  wr_cycle[20698] = 1'b0;  addr_rom[20698]='h00000368;  wr_data_rom[20698]='h00000000;
    rd_cycle[20699] = 1'b1;  wr_cycle[20699] = 1'b0;  addr_rom[20699]='h0000036c;  wr_data_rom[20699]='h00000000;
    rd_cycle[20700] = 1'b1;  wr_cycle[20700] = 1'b0;  addr_rom[20700]='h00000370;  wr_data_rom[20700]='h00000000;
    rd_cycle[20701] = 1'b1;  wr_cycle[20701] = 1'b0;  addr_rom[20701]='h00000374;  wr_data_rom[20701]='h00000000;
    rd_cycle[20702] = 1'b1;  wr_cycle[20702] = 1'b0;  addr_rom[20702]='h00000378;  wr_data_rom[20702]='h00000000;
    rd_cycle[20703] = 1'b1;  wr_cycle[20703] = 1'b0;  addr_rom[20703]='h0000037c;  wr_data_rom[20703]='h00000000;
    rd_cycle[20704] = 1'b1;  wr_cycle[20704] = 1'b0;  addr_rom[20704]='h00000380;  wr_data_rom[20704]='h00000000;
    rd_cycle[20705] = 1'b1;  wr_cycle[20705] = 1'b0;  addr_rom[20705]='h00000384;  wr_data_rom[20705]='h00000000;
    rd_cycle[20706] = 1'b1;  wr_cycle[20706] = 1'b0;  addr_rom[20706]='h00000388;  wr_data_rom[20706]='h00000000;
    rd_cycle[20707] = 1'b1;  wr_cycle[20707] = 1'b0;  addr_rom[20707]='h0000038c;  wr_data_rom[20707]='h00000000;
    rd_cycle[20708] = 1'b1;  wr_cycle[20708] = 1'b0;  addr_rom[20708]='h00000390;  wr_data_rom[20708]='h00000000;
    rd_cycle[20709] = 1'b1;  wr_cycle[20709] = 1'b0;  addr_rom[20709]='h00000394;  wr_data_rom[20709]='h00000000;
    rd_cycle[20710] = 1'b1;  wr_cycle[20710] = 1'b0;  addr_rom[20710]='h00000398;  wr_data_rom[20710]='h00000000;
    rd_cycle[20711] = 1'b1;  wr_cycle[20711] = 1'b0;  addr_rom[20711]='h0000039c;  wr_data_rom[20711]='h00000000;
    rd_cycle[20712] = 1'b1;  wr_cycle[20712] = 1'b0;  addr_rom[20712]='h000003a0;  wr_data_rom[20712]='h00000000;
    rd_cycle[20713] = 1'b1;  wr_cycle[20713] = 1'b0;  addr_rom[20713]='h000003a4;  wr_data_rom[20713]='h00000000;
    rd_cycle[20714] = 1'b1;  wr_cycle[20714] = 1'b0;  addr_rom[20714]='h000003a8;  wr_data_rom[20714]='h00000000;
    rd_cycle[20715] = 1'b1;  wr_cycle[20715] = 1'b0;  addr_rom[20715]='h000003ac;  wr_data_rom[20715]='h00000000;
    rd_cycle[20716] = 1'b1;  wr_cycle[20716] = 1'b0;  addr_rom[20716]='h000003b0;  wr_data_rom[20716]='h00000000;
    rd_cycle[20717] = 1'b1;  wr_cycle[20717] = 1'b0;  addr_rom[20717]='h000003b4;  wr_data_rom[20717]='h00000000;
    rd_cycle[20718] = 1'b1;  wr_cycle[20718] = 1'b0;  addr_rom[20718]='h000003b8;  wr_data_rom[20718]='h00000000;
    rd_cycle[20719] = 1'b1;  wr_cycle[20719] = 1'b0;  addr_rom[20719]='h000003bc;  wr_data_rom[20719]='h00000000;
    rd_cycle[20720] = 1'b1;  wr_cycle[20720] = 1'b0;  addr_rom[20720]='h000003c0;  wr_data_rom[20720]='h00000000;
    rd_cycle[20721] = 1'b1;  wr_cycle[20721] = 1'b0;  addr_rom[20721]='h000003c4;  wr_data_rom[20721]='h00000000;
    rd_cycle[20722] = 1'b1;  wr_cycle[20722] = 1'b0;  addr_rom[20722]='h000003c8;  wr_data_rom[20722]='h00000000;
    rd_cycle[20723] = 1'b1;  wr_cycle[20723] = 1'b0;  addr_rom[20723]='h000003cc;  wr_data_rom[20723]='h00000000;
    rd_cycle[20724] = 1'b1;  wr_cycle[20724] = 1'b0;  addr_rom[20724]='h000003d0;  wr_data_rom[20724]='h00000000;
    rd_cycle[20725] = 1'b1;  wr_cycle[20725] = 1'b0;  addr_rom[20725]='h000003d4;  wr_data_rom[20725]='h00000000;
    rd_cycle[20726] = 1'b1;  wr_cycle[20726] = 1'b0;  addr_rom[20726]='h000003d8;  wr_data_rom[20726]='h00000000;
    rd_cycle[20727] = 1'b1;  wr_cycle[20727] = 1'b0;  addr_rom[20727]='h000003dc;  wr_data_rom[20727]='h00000000;
    rd_cycle[20728] = 1'b1;  wr_cycle[20728] = 1'b0;  addr_rom[20728]='h000003e0;  wr_data_rom[20728]='h00000000;
    rd_cycle[20729] = 1'b1;  wr_cycle[20729] = 1'b0;  addr_rom[20729]='h000003e4;  wr_data_rom[20729]='h00000000;
    rd_cycle[20730] = 1'b1;  wr_cycle[20730] = 1'b0;  addr_rom[20730]='h000003e8;  wr_data_rom[20730]='h00000000;
    rd_cycle[20731] = 1'b1;  wr_cycle[20731] = 1'b0;  addr_rom[20731]='h000003ec;  wr_data_rom[20731]='h00000000;
    rd_cycle[20732] = 1'b1;  wr_cycle[20732] = 1'b0;  addr_rom[20732]='h000003f0;  wr_data_rom[20732]='h00000000;
    rd_cycle[20733] = 1'b1;  wr_cycle[20733] = 1'b0;  addr_rom[20733]='h000003f4;  wr_data_rom[20733]='h00000000;
    rd_cycle[20734] = 1'b1;  wr_cycle[20734] = 1'b0;  addr_rom[20734]='h000003f8;  wr_data_rom[20734]='h00000000;
    rd_cycle[20735] = 1'b1;  wr_cycle[20735] = 1'b0;  addr_rom[20735]='h000003fc;  wr_data_rom[20735]='h00000000;
    rd_cycle[20736] = 1'b1;  wr_cycle[20736] = 1'b0;  addr_rom[20736]='h00000400;  wr_data_rom[20736]='h00000000;
    rd_cycle[20737] = 1'b1;  wr_cycle[20737] = 1'b0;  addr_rom[20737]='h00000404;  wr_data_rom[20737]='h00000000;
    rd_cycle[20738] = 1'b1;  wr_cycle[20738] = 1'b0;  addr_rom[20738]='h00000408;  wr_data_rom[20738]='h00000000;
    rd_cycle[20739] = 1'b1;  wr_cycle[20739] = 1'b0;  addr_rom[20739]='h0000040c;  wr_data_rom[20739]='h00000000;
    rd_cycle[20740] = 1'b1;  wr_cycle[20740] = 1'b0;  addr_rom[20740]='h00000410;  wr_data_rom[20740]='h00000000;
    rd_cycle[20741] = 1'b1;  wr_cycle[20741] = 1'b0;  addr_rom[20741]='h00000414;  wr_data_rom[20741]='h00000000;
    rd_cycle[20742] = 1'b1;  wr_cycle[20742] = 1'b0;  addr_rom[20742]='h00000418;  wr_data_rom[20742]='h00000000;
    rd_cycle[20743] = 1'b1;  wr_cycle[20743] = 1'b0;  addr_rom[20743]='h0000041c;  wr_data_rom[20743]='h00000000;
    rd_cycle[20744] = 1'b1;  wr_cycle[20744] = 1'b0;  addr_rom[20744]='h00000420;  wr_data_rom[20744]='h00000000;
    rd_cycle[20745] = 1'b1;  wr_cycle[20745] = 1'b0;  addr_rom[20745]='h00000424;  wr_data_rom[20745]='h00000000;
    rd_cycle[20746] = 1'b1;  wr_cycle[20746] = 1'b0;  addr_rom[20746]='h00000428;  wr_data_rom[20746]='h00000000;
    rd_cycle[20747] = 1'b1;  wr_cycle[20747] = 1'b0;  addr_rom[20747]='h0000042c;  wr_data_rom[20747]='h00000000;
    rd_cycle[20748] = 1'b1;  wr_cycle[20748] = 1'b0;  addr_rom[20748]='h00000430;  wr_data_rom[20748]='h00000000;
    rd_cycle[20749] = 1'b1;  wr_cycle[20749] = 1'b0;  addr_rom[20749]='h00000434;  wr_data_rom[20749]='h00000000;
    rd_cycle[20750] = 1'b1;  wr_cycle[20750] = 1'b0;  addr_rom[20750]='h00000438;  wr_data_rom[20750]='h00000000;
    rd_cycle[20751] = 1'b1;  wr_cycle[20751] = 1'b0;  addr_rom[20751]='h0000043c;  wr_data_rom[20751]='h00000000;
    rd_cycle[20752] = 1'b1;  wr_cycle[20752] = 1'b0;  addr_rom[20752]='h00000440;  wr_data_rom[20752]='h00000000;
    rd_cycle[20753] = 1'b1;  wr_cycle[20753] = 1'b0;  addr_rom[20753]='h00000444;  wr_data_rom[20753]='h00000000;
    rd_cycle[20754] = 1'b1;  wr_cycle[20754] = 1'b0;  addr_rom[20754]='h00000448;  wr_data_rom[20754]='h00000000;
    rd_cycle[20755] = 1'b1;  wr_cycle[20755] = 1'b0;  addr_rom[20755]='h0000044c;  wr_data_rom[20755]='h00000000;
    rd_cycle[20756] = 1'b1;  wr_cycle[20756] = 1'b0;  addr_rom[20756]='h00000450;  wr_data_rom[20756]='h00000000;
    rd_cycle[20757] = 1'b1;  wr_cycle[20757] = 1'b0;  addr_rom[20757]='h00000454;  wr_data_rom[20757]='h00000000;
    rd_cycle[20758] = 1'b1;  wr_cycle[20758] = 1'b0;  addr_rom[20758]='h00000458;  wr_data_rom[20758]='h00000000;
    rd_cycle[20759] = 1'b1;  wr_cycle[20759] = 1'b0;  addr_rom[20759]='h0000045c;  wr_data_rom[20759]='h00000000;
    rd_cycle[20760] = 1'b1;  wr_cycle[20760] = 1'b0;  addr_rom[20760]='h00000460;  wr_data_rom[20760]='h00000000;
    rd_cycle[20761] = 1'b1;  wr_cycle[20761] = 1'b0;  addr_rom[20761]='h00000464;  wr_data_rom[20761]='h00000000;
    rd_cycle[20762] = 1'b1;  wr_cycle[20762] = 1'b0;  addr_rom[20762]='h00000468;  wr_data_rom[20762]='h00000000;
    rd_cycle[20763] = 1'b1;  wr_cycle[20763] = 1'b0;  addr_rom[20763]='h0000046c;  wr_data_rom[20763]='h00000000;
    rd_cycle[20764] = 1'b1;  wr_cycle[20764] = 1'b0;  addr_rom[20764]='h00000470;  wr_data_rom[20764]='h00000000;
    rd_cycle[20765] = 1'b1;  wr_cycle[20765] = 1'b0;  addr_rom[20765]='h00000474;  wr_data_rom[20765]='h00000000;
    rd_cycle[20766] = 1'b1;  wr_cycle[20766] = 1'b0;  addr_rom[20766]='h00000478;  wr_data_rom[20766]='h00000000;
    rd_cycle[20767] = 1'b1;  wr_cycle[20767] = 1'b0;  addr_rom[20767]='h0000047c;  wr_data_rom[20767]='h00000000;
    rd_cycle[20768] = 1'b1;  wr_cycle[20768] = 1'b0;  addr_rom[20768]='h00000480;  wr_data_rom[20768]='h00000000;
    rd_cycle[20769] = 1'b1;  wr_cycle[20769] = 1'b0;  addr_rom[20769]='h00000484;  wr_data_rom[20769]='h00000000;
    rd_cycle[20770] = 1'b1;  wr_cycle[20770] = 1'b0;  addr_rom[20770]='h00000488;  wr_data_rom[20770]='h00000000;
    rd_cycle[20771] = 1'b1;  wr_cycle[20771] = 1'b0;  addr_rom[20771]='h0000048c;  wr_data_rom[20771]='h00000000;
    rd_cycle[20772] = 1'b1;  wr_cycle[20772] = 1'b0;  addr_rom[20772]='h00000490;  wr_data_rom[20772]='h00000000;
    rd_cycle[20773] = 1'b1;  wr_cycle[20773] = 1'b0;  addr_rom[20773]='h00000494;  wr_data_rom[20773]='h00000000;
    rd_cycle[20774] = 1'b1;  wr_cycle[20774] = 1'b0;  addr_rom[20774]='h00000498;  wr_data_rom[20774]='h00000000;
    rd_cycle[20775] = 1'b1;  wr_cycle[20775] = 1'b0;  addr_rom[20775]='h0000049c;  wr_data_rom[20775]='h00000000;
    rd_cycle[20776] = 1'b1;  wr_cycle[20776] = 1'b0;  addr_rom[20776]='h000004a0;  wr_data_rom[20776]='h00000000;
    rd_cycle[20777] = 1'b1;  wr_cycle[20777] = 1'b0;  addr_rom[20777]='h000004a4;  wr_data_rom[20777]='h00000000;
    rd_cycle[20778] = 1'b1;  wr_cycle[20778] = 1'b0;  addr_rom[20778]='h000004a8;  wr_data_rom[20778]='h00000000;
    rd_cycle[20779] = 1'b1;  wr_cycle[20779] = 1'b0;  addr_rom[20779]='h000004ac;  wr_data_rom[20779]='h00000000;
    rd_cycle[20780] = 1'b1;  wr_cycle[20780] = 1'b0;  addr_rom[20780]='h000004b0;  wr_data_rom[20780]='h00000000;
    rd_cycle[20781] = 1'b1;  wr_cycle[20781] = 1'b0;  addr_rom[20781]='h000004b4;  wr_data_rom[20781]='h00000000;
    rd_cycle[20782] = 1'b1;  wr_cycle[20782] = 1'b0;  addr_rom[20782]='h000004b8;  wr_data_rom[20782]='h00000000;
    rd_cycle[20783] = 1'b1;  wr_cycle[20783] = 1'b0;  addr_rom[20783]='h000004bc;  wr_data_rom[20783]='h00000000;
    rd_cycle[20784] = 1'b1;  wr_cycle[20784] = 1'b0;  addr_rom[20784]='h000004c0;  wr_data_rom[20784]='h00000000;
    rd_cycle[20785] = 1'b1;  wr_cycle[20785] = 1'b0;  addr_rom[20785]='h000004c4;  wr_data_rom[20785]='h00000000;
    rd_cycle[20786] = 1'b1;  wr_cycle[20786] = 1'b0;  addr_rom[20786]='h000004c8;  wr_data_rom[20786]='h00000000;
    rd_cycle[20787] = 1'b1;  wr_cycle[20787] = 1'b0;  addr_rom[20787]='h000004cc;  wr_data_rom[20787]='h00000000;
    rd_cycle[20788] = 1'b1;  wr_cycle[20788] = 1'b0;  addr_rom[20788]='h000004d0;  wr_data_rom[20788]='h00000000;
    rd_cycle[20789] = 1'b1;  wr_cycle[20789] = 1'b0;  addr_rom[20789]='h000004d4;  wr_data_rom[20789]='h00000000;
    rd_cycle[20790] = 1'b1;  wr_cycle[20790] = 1'b0;  addr_rom[20790]='h000004d8;  wr_data_rom[20790]='h00000000;
    rd_cycle[20791] = 1'b1;  wr_cycle[20791] = 1'b0;  addr_rom[20791]='h000004dc;  wr_data_rom[20791]='h00000000;
    rd_cycle[20792] = 1'b1;  wr_cycle[20792] = 1'b0;  addr_rom[20792]='h000004e0;  wr_data_rom[20792]='h00000000;
    rd_cycle[20793] = 1'b1;  wr_cycle[20793] = 1'b0;  addr_rom[20793]='h000004e4;  wr_data_rom[20793]='h00000000;
    rd_cycle[20794] = 1'b1;  wr_cycle[20794] = 1'b0;  addr_rom[20794]='h000004e8;  wr_data_rom[20794]='h00000000;
    rd_cycle[20795] = 1'b1;  wr_cycle[20795] = 1'b0;  addr_rom[20795]='h000004ec;  wr_data_rom[20795]='h00000000;
    rd_cycle[20796] = 1'b1;  wr_cycle[20796] = 1'b0;  addr_rom[20796]='h000004f0;  wr_data_rom[20796]='h00000000;
    rd_cycle[20797] = 1'b1;  wr_cycle[20797] = 1'b0;  addr_rom[20797]='h000004f4;  wr_data_rom[20797]='h00000000;
    rd_cycle[20798] = 1'b1;  wr_cycle[20798] = 1'b0;  addr_rom[20798]='h000004f8;  wr_data_rom[20798]='h00000000;
    rd_cycle[20799] = 1'b1;  wr_cycle[20799] = 1'b0;  addr_rom[20799]='h000004fc;  wr_data_rom[20799]='h00000000;
    rd_cycle[20800] = 1'b1;  wr_cycle[20800] = 1'b0;  addr_rom[20800]='h00000500;  wr_data_rom[20800]='h00000000;
    rd_cycle[20801] = 1'b1;  wr_cycle[20801] = 1'b0;  addr_rom[20801]='h00000504;  wr_data_rom[20801]='h00000000;
    rd_cycle[20802] = 1'b1;  wr_cycle[20802] = 1'b0;  addr_rom[20802]='h00000508;  wr_data_rom[20802]='h00000000;
    rd_cycle[20803] = 1'b1;  wr_cycle[20803] = 1'b0;  addr_rom[20803]='h0000050c;  wr_data_rom[20803]='h00000000;
    rd_cycle[20804] = 1'b1;  wr_cycle[20804] = 1'b0;  addr_rom[20804]='h00000510;  wr_data_rom[20804]='h00000000;
    rd_cycle[20805] = 1'b1;  wr_cycle[20805] = 1'b0;  addr_rom[20805]='h00000514;  wr_data_rom[20805]='h00000000;
    rd_cycle[20806] = 1'b1;  wr_cycle[20806] = 1'b0;  addr_rom[20806]='h00000518;  wr_data_rom[20806]='h00000000;
    rd_cycle[20807] = 1'b1;  wr_cycle[20807] = 1'b0;  addr_rom[20807]='h0000051c;  wr_data_rom[20807]='h00000000;
    rd_cycle[20808] = 1'b1;  wr_cycle[20808] = 1'b0;  addr_rom[20808]='h00000520;  wr_data_rom[20808]='h00000000;
    rd_cycle[20809] = 1'b1;  wr_cycle[20809] = 1'b0;  addr_rom[20809]='h00000524;  wr_data_rom[20809]='h00000000;
    rd_cycle[20810] = 1'b1;  wr_cycle[20810] = 1'b0;  addr_rom[20810]='h00000528;  wr_data_rom[20810]='h00000000;
    rd_cycle[20811] = 1'b1;  wr_cycle[20811] = 1'b0;  addr_rom[20811]='h0000052c;  wr_data_rom[20811]='h00000000;
    rd_cycle[20812] = 1'b1;  wr_cycle[20812] = 1'b0;  addr_rom[20812]='h00000530;  wr_data_rom[20812]='h00000000;
    rd_cycle[20813] = 1'b1;  wr_cycle[20813] = 1'b0;  addr_rom[20813]='h00000534;  wr_data_rom[20813]='h00000000;
    rd_cycle[20814] = 1'b1;  wr_cycle[20814] = 1'b0;  addr_rom[20814]='h00000538;  wr_data_rom[20814]='h00000000;
    rd_cycle[20815] = 1'b1;  wr_cycle[20815] = 1'b0;  addr_rom[20815]='h0000053c;  wr_data_rom[20815]='h00000000;
    rd_cycle[20816] = 1'b1;  wr_cycle[20816] = 1'b0;  addr_rom[20816]='h00000540;  wr_data_rom[20816]='h00000000;
    rd_cycle[20817] = 1'b1;  wr_cycle[20817] = 1'b0;  addr_rom[20817]='h00000544;  wr_data_rom[20817]='h00000000;
    rd_cycle[20818] = 1'b1;  wr_cycle[20818] = 1'b0;  addr_rom[20818]='h00000548;  wr_data_rom[20818]='h00000000;
    rd_cycle[20819] = 1'b1;  wr_cycle[20819] = 1'b0;  addr_rom[20819]='h0000054c;  wr_data_rom[20819]='h00000000;
    rd_cycle[20820] = 1'b1;  wr_cycle[20820] = 1'b0;  addr_rom[20820]='h00000550;  wr_data_rom[20820]='h00000000;
    rd_cycle[20821] = 1'b1;  wr_cycle[20821] = 1'b0;  addr_rom[20821]='h00000554;  wr_data_rom[20821]='h00000000;
    rd_cycle[20822] = 1'b1;  wr_cycle[20822] = 1'b0;  addr_rom[20822]='h00000558;  wr_data_rom[20822]='h00000000;
    rd_cycle[20823] = 1'b1;  wr_cycle[20823] = 1'b0;  addr_rom[20823]='h0000055c;  wr_data_rom[20823]='h00000000;
    rd_cycle[20824] = 1'b1;  wr_cycle[20824] = 1'b0;  addr_rom[20824]='h00000560;  wr_data_rom[20824]='h00000000;
    rd_cycle[20825] = 1'b1;  wr_cycle[20825] = 1'b0;  addr_rom[20825]='h00000564;  wr_data_rom[20825]='h00000000;
    rd_cycle[20826] = 1'b1;  wr_cycle[20826] = 1'b0;  addr_rom[20826]='h00000568;  wr_data_rom[20826]='h00000000;
    rd_cycle[20827] = 1'b1;  wr_cycle[20827] = 1'b0;  addr_rom[20827]='h0000056c;  wr_data_rom[20827]='h00000000;
    rd_cycle[20828] = 1'b1;  wr_cycle[20828] = 1'b0;  addr_rom[20828]='h00000570;  wr_data_rom[20828]='h00000000;
    rd_cycle[20829] = 1'b1;  wr_cycle[20829] = 1'b0;  addr_rom[20829]='h00000574;  wr_data_rom[20829]='h00000000;
    rd_cycle[20830] = 1'b1;  wr_cycle[20830] = 1'b0;  addr_rom[20830]='h00000578;  wr_data_rom[20830]='h00000000;
    rd_cycle[20831] = 1'b1;  wr_cycle[20831] = 1'b0;  addr_rom[20831]='h0000057c;  wr_data_rom[20831]='h00000000;
    rd_cycle[20832] = 1'b1;  wr_cycle[20832] = 1'b0;  addr_rom[20832]='h00000580;  wr_data_rom[20832]='h00000000;
    rd_cycle[20833] = 1'b1;  wr_cycle[20833] = 1'b0;  addr_rom[20833]='h00000584;  wr_data_rom[20833]='h00000000;
    rd_cycle[20834] = 1'b1;  wr_cycle[20834] = 1'b0;  addr_rom[20834]='h00000588;  wr_data_rom[20834]='h00000000;
    rd_cycle[20835] = 1'b1;  wr_cycle[20835] = 1'b0;  addr_rom[20835]='h0000058c;  wr_data_rom[20835]='h00000000;
    rd_cycle[20836] = 1'b1;  wr_cycle[20836] = 1'b0;  addr_rom[20836]='h00000590;  wr_data_rom[20836]='h00000000;
    rd_cycle[20837] = 1'b1;  wr_cycle[20837] = 1'b0;  addr_rom[20837]='h00000594;  wr_data_rom[20837]='h00000000;
    rd_cycle[20838] = 1'b1;  wr_cycle[20838] = 1'b0;  addr_rom[20838]='h00000598;  wr_data_rom[20838]='h00000000;
    rd_cycle[20839] = 1'b1;  wr_cycle[20839] = 1'b0;  addr_rom[20839]='h0000059c;  wr_data_rom[20839]='h00000000;
    rd_cycle[20840] = 1'b1;  wr_cycle[20840] = 1'b0;  addr_rom[20840]='h000005a0;  wr_data_rom[20840]='h00000000;
    rd_cycle[20841] = 1'b1;  wr_cycle[20841] = 1'b0;  addr_rom[20841]='h000005a4;  wr_data_rom[20841]='h00000000;
    rd_cycle[20842] = 1'b1;  wr_cycle[20842] = 1'b0;  addr_rom[20842]='h000005a8;  wr_data_rom[20842]='h00000000;
    rd_cycle[20843] = 1'b1;  wr_cycle[20843] = 1'b0;  addr_rom[20843]='h000005ac;  wr_data_rom[20843]='h00000000;
    rd_cycle[20844] = 1'b1;  wr_cycle[20844] = 1'b0;  addr_rom[20844]='h000005b0;  wr_data_rom[20844]='h00000000;
    rd_cycle[20845] = 1'b1;  wr_cycle[20845] = 1'b0;  addr_rom[20845]='h000005b4;  wr_data_rom[20845]='h00000000;
    rd_cycle[20846] = 1'b1;  wr_cycle[20846] = 1'b0;  addr_rom[20846]='h000005b8;  wr_data_rom[20846]='h00000000;
    rd_cycle[20847] = 1'b1;  wr_cycle[20847] = 1'b0;  addr_rom[20847]='h000005bc;  wr_data_rom[20847]='h00000000;
    rd_cycle[20848] = 1'b1;  wr_cycle[20848] = 1'b0;  addr_rom[20848]='h000005c0;  wr_data_rom[20848]='h00000000;
    rd_cycle[20849] = 1'b1;  wr_cycle[20849] = 1'b0;  addr_rom[20849]='h000005c4;  wr_data_rom[20849]='h00000000;
    rd_cycle[20850] = 1'b1;  wr_cycle[20850] = 1'b0;  addr_rom[20850]='h000005c8;  wr_data_rom[20850]='h00000000;
    rd_cycle[20851] = 1'b1;  wr_cycle[20851] = 1'b0;  addr_rom[20851]='h000005cc;  wr_data_rom[20851]='h00000000;
    rd_cycle[20852] = 1'b1;  wr_cycle[20852] = 1'b0;  addr_rom[20852]='h000005d0;  wr_data_rom[20852]='h00000000;
    rd_cycle[20853] = 1'b1;  wr_cycle[20853] = 1'b0;  addr_rom[20853]='h000005d4;  wr_data_rom[20853]='h00000000;
    rd_cycle[20854] = 1'b1;  wr_cycle[20854] = 1'b0;  addr_rom[20854]='h000005d8;  wr_data_rom[20854]='h00000000;
    rd_cycle[20855] = 1'b1;  wr_cycle[20855] = 1'b0;  addr_rom[20855]='h000005dc;  wr_data_rom[20855]='h00000000;
    rd_cycle[20856] = 1'b1;  wr_cycle[20856] = 1'b0;  addr_rom[20856]='h000005e0;  wr_data_rom[20856]='h00000000;
    rd_cycle[20857] = 1'b1;  wr_cycle[20857] = 1'b0;  addr_rom[20857]='h000005e4;  wr_data_rom[20857]='h00000000;
    rd_cycle[20858] = 1'b1;  wr_cycle[20858] = 1'b0;  addr_rom[20858]='h000005e8;  wr_data_rom[20858]='h00000000;
    rd_cycle[20859] = 1'b1;  wr_cycle[20859] = 1'b0;  addr_rom[20859]='h000005ec;  wr_data_rom[20859]='h00000000;
    rd_cycle[20860] = 1'b1;  wr_cycle[20860] = 1'b0;  addr_rom[20860]='h000005f0;  wr_data_rom[20860]='h00000000;
    rd_cycle[20861] = 1'b1;  wr_cycle[20861] = 1'b0;  addr_rom[20861]='h000005f4;  wr_data_rom[20861]='h00000000;
    rd_cycle[20862] = 1'b1;  wr_cycle[20862] = 1'b0;  addr_rom[20862]='h000005f8;  wr_data_rom[20862]='h00000000;
    rd_cycle[20863] = 1'b1;  wr_cycle[20863] = 1'b0;  addr_rom[20863]='h000005fc;  wr_data_rom[20863]='h00000000;
    rd_cycle[20864] = 1'b1;  wr_cycle[20864] = 1'b0;  addr_rom[20864]='h00000600;  wr_data_rom[20864]='h00000000;
    rd_cycle[20865] = 1'b1;  wr_cycle[20865] = 1'b0;  addr_rom[20865]='h00000604;  wr_data_rom[20865]='h00000000;
    rd_cycle[20866] = 1'b1;  wr_cycle[20866] = 1'b0;  addr_rom[20866]='h00000608;  wr_data_rom[20866]='h00000000;
    rd_cycle[20867] = 1'b1;  wr_cycle[20867] = 1'b0;  addr_rom[20867]='h0000060c;  wr_data_rom[20867]='h00000000;
    rd_cycle[20868] = 1'b1;  wr_cycle[20868] = 1'b0;  addr_rom[20868]='h00000610;  wr_data_rom[20868]='h00000000;
    rd_cycle[20869] = 1'b1;  wr_cycle[20869] = 1'b0;  addr_rom[20869]='h00000614;  wr_data_rom[20869]='h00000000;
    rd_cycle[20870] = 1'b1;  wr_cycle[20870] = 1'b0;  addr_rom[20870]='h00000618;  wr_data_rom[20870]='h00000000;
    rd_cycle[20871] = 1'b1;  wr_cycle[20871] = 1'b0;  addr_rom[20871]='h0000061c;  wr_data_rom[20871]='h00000000;
    rd_cycle[20872] = 1'b1;  wr_cycle[20872] = 1'b0;  addr_rom[20872]='h00000620;  wr_data_rom[20872]='h00000000;
    rd_cycle[20873] = 1'b1;  wr_cycle[20873] = 1'b0;  addr_rom[20873]='h00000624;  wr_data_rom[20873]='h00000000;
    rd_cycle[20874] = 1'b1;  wr_cycle[20874] = 1'b0;  addr_rom[20874]='h00000628;  wr_data_rom[20874]='h00000000;
    rd_cycle[20875] = 1'b1;  wr_cycle[20875] = 1'b0;  addr_rom[20875]='h0000062c;  wr_data_rom[20875]='h00000000;
    rd_cycle[20876] = 1'b1;  wr_cycle[20876] = 1'b0;  addr_rom[20876]='h00000630;  wr_data_rom[20876]='h00000000;
    rd_cycle[20877] = 1'b1;  wr_cycle[20877] = 1'b0;  addr_rom[20877]='h00000634;  wr_data_rom[20877]='h00000000;
    rd_cycle[20878] = 1'b1;  wr_cycle[20878] = 1'b0;  addr_rom[20878]='h00000638;  wr_data_rom[20878]='h00000000;
    rd_cycle[20879] = 1'b1;  wr_cycle[20879] = 1'b0;  addr_rom[20879]='h0000063c;  wr_data_rom[20879]='h00000000;
    rd_cycle[20880] = 1'b1;  wr_cycle[20880] = 1'b0;  addr_rom[20880]='h00000640;  wr_data_rom[20880]='h00000000;
    rd_cycle[20881] = 1'b1;  wr_cycle[20881] = 1'b0;  addr_rom[20881]='h00000644;  wr_data_rom[20881]='h00000000;
    rd_cycle[20882] = 1'b1;  wr_cycle[20882] = 1'b0;  addr_rom[20882]='h00000648;  wr_data_rom[20882]='h00000000;
    rd_cycle[20883] = 1'b1;  wr_cycle[20883] = 1'b0;  addr_rom[20883]='h0000064c;  wr_data_rom[20883]='h00000000;
    rd_cycle[20884] = 1'b1;  wr_cycle[20884] = 1'b0;  addr_rom[20884]='h00000650;  wr_data_rom[20884]='h00000000;
    rd_cycle[20885] = 1'b1;  wr_cycle[20885] = 1'b0;  addr_rom[20885]='h00000654;  wr_data_rom[20885]='h00000000;
    rd_cycle[20886] = 1'b1;  wr_cycle[20886] = 1'b0;  addr_rom[20886]='h00000658;  wr_data_rom[20886]='h00000000;
    rd_cycle[20887] = 1'b1;  wr_cycle[20887] = 1'b0;  addr_rom[20887]='h0000065c;  wr_data_rom[20887]='h00000000;
    rd_cycle[20888] = 1'b1;  wr_cycle[20888] = 1'b0;  addr_rom[20888]='h00000660;  wr_data_rom[20888]='h00000000;
    rd_cycle[20889] = 1'b1;  wr_cycle[20889] = 1'b0;  addr_rom[20889]='h00000664;  wr_data_rom[20889]='h00000000;
    rd_cycle[20890] = 1'b1;  wr_cycle[20890] = 1'b0;  addr_rom[20890]='h00000668;  wr_data_rom[20890]='h00000000;
    rd_cycle[20891] = 1'b1;  wr_cycle[20891] = 1'b0;  addr_rom[20891]='h0000066c;  wr_data_rom[20891]='h00000000;
    rd_cycle[20892] = 1'b1;  wr_cycle[20892] = 1'b0;  addr_rom[20892]='h00000670;  wr_data_rom[20892]='h00000000;
    rd_cycle[20893] = 1'b1;  wr_cycle[20893] = 1'b0;  addr_rom[20893]='h00000674;  wr_data_rom[20893]='h00000000;
    rd_cycle[20894] = 1'b1;  wr_cycle[20894] = 1'b0;  addr_rom[20894]='h00000678;  wr_data_rom[20894]='h00000000;
    rd_cycle[20895] = 1'b1;  wr_cycle[20895] = 1'b0;  addr_rom[20895]='h0000067c;  wr_data_rom[20895]='h00000000;
    rd_cycle[20896] = 1'b1;  wr_cycle[20896] = 1'b0;  addr_rom[20896]='h00000680;  wr_data_rom[20896]='h00000000;
    rd_cycle[20897] = 1'b1;  wr_cycle[20897] = 1'b0;  addr_rom[20897]='h00000684;  wr_data_rom[20897]='h00000000;
    rd_cycle[20898] = 1'b1;  wr_cycle[20898] = 1'b0;  addr_rom[20898]='h00000688;  wr_data_rom[20898]='h00000000;
    rd_cycle[20899] = 1'b1;  wr_cycle[20899] = 1'b0;  addr_rom[20899]='h0000068c;  wr_data_rom[20899]='h00000000;
    rd_cycle[20900] = 1'b1;  wr_cycle[20900] = 1'b0;  addr_rom[20900]='h00000690;  wr_data_rom[20900]='h00000000;
    rd_cycle[20901] = 1'b1;  wr_cycle[20901] = 1'b0;  addr_rom[20901]='h00000694;  wr_data_rom[20901]='h00000000;
    rd_cycle[20902] = 1'b1;  wr_cycle[20902] = 1'b0;  addr_rom[20902]='h00000698;  wr_data_rom[20902]='h00000000;
    rd_cycle[20903] = 1'b1;  wr_cycle[20903] = 1'b0;  addr_rom[20903]='h0000069c;  wr_data_rom[20903]='h00000000;
    rd_cycle[20904] = 1'b1;  wr_cycle[20904] = 1'b0;  addr_rom[20904]='h000006a0;  wr_data_rom[20904]='h00000000;
    rd_cycle[20905] = 1'b1;  wr_cycle[20905] = 1'b0;  addr_rom[20905]='h000006a4;  wr_data_rom[20905]='h00000000;
    rd_cycle[20906] = 1'b1;  wr_cycle[20906] = 1'b0;  addr_rom[20906]='h000006a8;  wr_data_rom[20906]='h00000000;
    rd_cycle[20907] = 1'b1;  wr_cycle[20907] = 1'b0;  addr_rom[20907]='h000006ac;  wr_data_rom[20907]='h00000000;
    rd_cycle[20908] = 1'b1;  wr_cycle[20908] = 1'b0;  addr_rom[20908]='h000006b0;  wr_data_rom[20908]='h00000000;
    rd_cycle[20909] = 1'b1;  wr_cycle[20909] = 1'b0;  addr_rom[20909]='h000006b4;  wr_data_rom[20909]='h00000000;
    rd_cycle[20910] = 1'b1;  wr_cycle[20910] = 1'b0;  addr_rom[20910]='h000006b8;  wr_data_rom[20910]='h00000000;
    rd_cycle[20911] = 1'b1;  wr_cycle[20911] = 1'b0;  addr_rom[20911]='h000006bc;  wr_data_rom[20911]='h00000000;
    rd_cycle[20912] = 1'b1;  wr_cycle[20912] = 1'b0;  addr_rom[20912]='h000006c0;  wr_data_rom[20912]='h00000000;
    rd_cycle[20913] = 1'b1;  wr_cycle[20913] = 1'b0;  addr_rom[20913]='h000006c4;  wr_data_rom[20913]='h00000000;
    rd_cycle[20914] = 1'b1;  wr_cycle[20914] = 1'b0;  addr_rom[20914]='h000006c8;  wr_data_rom[20914]='h00000000;
    rd_cycle[20915] = 1'b1;  wr_cycle[20915] = 1'b0;  addr_rom[20915]='h000006cc;  wr_data_rom[20915]='h00000000;
    rd_cycle[20916] = 1'b1;  wr_cycle[20916] = 1'b0;  addr_rom[20916]='h000006d0;  wr_data_rom[20916]='h00000000;
    rd_cycle[20917] = 1'b1;  wr_cycle[20917] = 1'b0;  addr_rom[20917]='h000006d4;  wr_data_rom[20917]='h00000000;
    rd_cycle[20918] = 1'b1;  wr_cycle[20918] = 1'b0;  addr_rom[20918]='h000006d8;  wr_data_rom[20918]='h00000000;
    rd_cycle[20919] = 1'b1;  wr_cycle[20919] = 1'b0;  addr_rom[20919]='h000006dc;  wr_data_rom[20919]='h00000000;
    rd_cycle[20920] = 1'b1;  wr_cycle[20920] = 1'b0;  addr_rom[20920]='h000006e0;  wr_data_rom[20920]='h00000000;
    rd_cycle[20921] = 1'b1;  wr_cycle[20921] = 1'b0;  addr_rom[20921]='h000006e4;  wr_data_rom[20921]='h00000000;
    rd_cycle[20922] = 1'b1;  wr_cycle[20922] = 1'b0;  addr_rom[20922]='h000006e8;  wr_data_rom[20922]='h00000000;
    rd_cycle[20923] = 1'b1;  wr_cycle[20923] = 1'b0;  addr_rom[20923]='h000006ec;  wr_data_rom[20923]='h00000000;
    rd_cycle[20924] = 1'b1;  wr_cycle[20924] = 1'b0;  addr_rom[20924]='h000006f0;  wr_data_rom[20924]='h00000000;
    rd_cycle[20925] = 1'b1;  wr_cycle[20925] = 1'b0;  addr_rom[20925]='h000006f4;  wr_data_rom[20925]='h00000000;
    rd_cycle[20926] = 1'b1;  wr_cycle[20926] = 1'b0;  addr_rom[20926]='h000006f8;  wr_data_rom[20926]='h00000000;
    rd_cycle[20927] = 1'b1;  wr_cycle[20927] = 1'b0;  addr_rom[20927]='h000006fc;  wr_data_rom[20927]='h00000000;
    rd_cycle[20928] = 1'b1;  wr_cycle[20928] = 1'b0;  addr_rom[20928]='h00000700;  wr_data_rom[20928]='h00000000;
    rd_cycle[20929] = 1'b1;  wr_cycle[20929] = 1'b0;  addr_rom[20929]='h00000704;  wr_data_rom[20929]='h00000000;
    rd_cycle[20930] = 1'b1;  wr_cycle[20930] = 1'b0;  addr_rom[20930]='h00000708;  wr_data_rom[20930]='h00000000;
    rd_cycle[20931] = 1'b1;  wr_cycle[20931] = 1'b0;  addr_rom[20931]='h0000070c;  wr_data_rom[20931]='h00000000;
    rd_cycle[20932] = 1'b1;  wr_cycle[20932] = 1'b0;  addr_rom[20932]='h00000710;  wr_data_rom[20932]='h00000000;
    rd_cycle[20933] = 1'b1;  wr_cycle[20933] = 1'b0;  addr_rom[20933]='h00000714;  wr_data_rom[20933]='h00000000;
    rd_cycle[20934] = 1'b1;  wr_cycle[20934] = 1'b0;  addr_rom[20934]='h00000718;  wr_data_rom[20934]='h00000000;
    rd_cycle[20935] = 1'b1;  wr_cycle[20935] = 1'b0;  addr_rom[20935]='h0000071c;  wr_data_rom[20935]='h00000000;
    rd_cycle[20936] = 1'b1;  wr_cycle[20936] = 1'b0;  addr_rom[20936]='h00000720;  wr_data_rom[20936]='h00000000;
    rd_cycle[20937] = 1'b1;  wr_cycle[20937] = 1'b0;  addr_rom[20937]='h00000724;  wr_data_rom[20937]='h00000000;
    rd_cycle[20938] = 1'b1;  wr_cycle[20938] = 1'b0;  addr_rom[20938]='h00000728;  wr_data_rom[20938]='h00000000;
    rd_cycle[20939] = 1'b1;  wr_cycle[20939] = 1'b0;  addr_rom[20939]='h0000072c;  wr_data_rom[20939]='h00000000;
    rd_cycle[20940] = 1'b1;  wr_cycle[20940] = 1'b0;  addr_rom[20940]='h00000730;  wr_data_rom[20940]='h00000000;
    rd_cycle[20941] = 1'b1;  wr_cycle[20941] = 1'b0;  addr_rom[20941]='h00000734;  wr_data_rom[20941]='h00000000;
    rd_cycle[20942] = 1'b1;  wr_cycle[20942] = 1'b0;  addr_rom[20942]='h00000738;  wr_data_rom[20942]='h00000000;
    rd_cycle[20943] = 1'b1;  wr_cycle[20943] = 1'b0;  addr_rom[20943]='h0000073c;  wr_data_rom[20943]='h00000000;
    rd_cycle[20944] = 1'b1;  wr_cycle[20944] = 1'b0;  addr_rom[20944]='h00000740;  wr_data_rom[20944]='h00000000;
    rd_cycle[20945] = 1'b1;  wr_cycle[20945] = 1'b0;  addr_rom[20945]='h00000744;  wr_data_rom[20945]='h00000000;
    rd_cycle[20946] = 1'b1;  wr_cycle[20946] = 1'b0;  addr_rom[20946]='h00000748;  wr_data_rom[20946]='h00000000;
    rd_cycle[20947] = 1'b1;  wr_cycle[20947] = 1'b0;  addr_rom[20947]='h0000074c;  wr_data_rom[20947]='h00000000;
    rd_cycle[20948] = 1'b1;  wr_cycle[20948] = 1'b0;  addr_rom[20948]='h00000750;  wr_data_rom[20948]='h00000000;
    rd_cycle[20949] = 1'b1;  wr_cycle[20949] = 1'b0;  addr_rom[20949]='h00000754;  wr_data_rom[20949]='h00000000;
    rd_cycle[20950] = 1'b1;  wr_cycle[20950] = 1'b0;  addr_rom[20950]='h00000758;  wr_data_rom[20950]='h00000000;
    rd_cycle[20951] = 1'b1;  wr_cycle[20951] = 1'b0;  addr_rom[20951]='h0000075c;  wr_data_rom[20951]='h00000000;
    rd_cycle[20952] = 1'b1;  wr_cycle[20952] = 1'b0;  addr_rom[20952]='h00000760;  wr_data_rom[20952]='h00000000;
    rd_cycle[20953] = 1'b1;  wr_cycle[20953] = 1'b0;  addr_rom[20953]='h00000764;  wr_data_rom[20953]='h00000000;
    rd_cycle[20954] = 1'b1;  wr_cycle[20954] = 1'b0;  addr_rom[20954]='h00000768;  wr_data_rom[20954]='h00000000;
    rd_cycle[20955] = 1'b1;  wr_cycle[20955] = 1'b0;  addr_rom[20955]='h0000076c;  wr_data_rom[20955]='h00000000;
    rd_cycle[20956] = 1'b1;  wr_cycle[20956] = 1'b0;  addr_rom[20956]='h00000770;  wr_data_rom[20956]='h00000000;
    rd_cycle[20957] = 1'b1;  wr_cycle[20957] = 1'b0;  addr_rom[20957]='h00000774;  wr_data_rom[20957]='h00000000;
    rd_cycle[20958] = 1'b1;  wr_cycle[20958] = 1'b0;  addr_rom[20958]='h00000778;  wr_data_rom[20958]='h00000000;
    rd_cycle[20959] = 1'b1;  wr_cycle[20959] = 1'b0;  addr_rom[20959]='h0000077c;  wr_data_rom[20959]='h00000000;
    rd_cycle[20960] = 1'b1;  wr_cycle[20960] = 1'b0;  addr_rom[20960]='h00000780;  wr_data_rom[20960]='h00000000;
    rd_cycle[20961] = 1'b1;  wr_cycle[20961] = 1'b0;  addr_rom[20961]='h00000784;  wr_data_rom[20961]='h00000000;
    rd_cycle[20962] = 1'b1;  wr_cycle[20962] = 1'b0;  addr_rom[20962]='h00000788;  wr_data_rom[20962]='h00000000;
    rd_cycle[20963] = 1'b1;  wr_cycle[20963] = 1'b0;  addr_rom[20963]='h0000078c;  wr_data_rom[20963]='h00000000;
    rd_cycle[20964] = 1'b1;  wr_cycle[20964] = 1'b0;  addr_rom[20964]='h00000790;  wr_data_rom[20964]='h00000000;
    rd_cycle[20965] = 1'b1;  wr_cycle[20965] = 1'b0;  addr_rom[20965]='h00000794;  wr_data_rom[20965]='h00000000;
    rd_cycle[20966] = 1'b1;  wr_cycle[20966] = 1'b0;  addr_rom[20966]='h00000798;  wr_data_rom[20966]='h00000000;
    rd_cycle[20967] = 1'b1;  wr_cycle[20967] = 1'b0;  addr_rom[20967]='h0000079c;  wr_data_rom[20967]='h00000000;
    rd_cycle[20968] = 1'b1;  wr_cycle[20968] = 1'b0;  addr_rom[20968]='h000007a0;  wr_data_rom[20968]='h00000000;
    rd_cycle[20969] = 1'b1;  wr_cycle[20969] = 1'b0;  addr_rom[20969]='h000007a4;  wr_data_rom[20969]='h00000000;
    rd_cycle[20970] = 1'b1;  wr_cycle[20970] = 1'b0;  addr_rom[20970]='h000007a8;  wr_data_rom[20970]='h00000000;
    rd_cycle[20971] = 1'b1;  wr_cycle[20971] = 1'b0;  addr_rom[20971]='h000007ac;  wr_data_rom[20971]='h00000000;
    rd_cycle[20972] = 1'b1;  wr_cycle[20972] = 1'b0;  addr_rom[20972]='h000007b0;  wr_data_rom[20972]='h00000000;
    rd_cycle[20973] = 1'b1;  wr_cycle[20973] = 1'b0;  addr_rom[20973]='h000007b4;  wr_data_rom[20973]='h00000000;
    rd_cycle[20974] = 1'b1;  wr_cycle[20974] = 1'b0;  addr_rom[20974]='h000007b8;  wr_data_rom[20974]='h00000000;
    rd_cycle[20975] = 1'b1;  wr_cycle[20975] = 1'b0;  addr_rom[20975]='h000007bc;  wr_data_rom[20975]='h00000000;
    rd_cycle[20976] = 1'b1;  wr_cycle[20976] = 1'b0;  addr_rom[20976]='h000007c0;  wr_data_rom[20976]='h00000000;
    rd_cycle[20977] = 1'b1;  wr_cycle[20977] = 1'b0;  addr_rom[20977]='h000007c4;  wr_data_rom[20977]='h00000000;
    rd_cycle[20978] = 1'b1;  wr_cycle[20978] = 1'b0;  addr_rom[20978]='h000007c8;  wr_data_rom[20978]='h00000000;
    rd_cycle[20979] = 1'b1;  wr_cycle[20979] = 1'b0;  addr_rom[20979]='h000007cc;  wr_data_rom[20979]='h00000000;
    rd_cycle[20980] = 1'b1;  wr_cycle[20980] = 1'b0;  addr_rom[20980]='h000007d0;  wr_data_rom[20980]='h00000000;
    rd_cycle[20981] = 1'b1;  wr_cycle[20981] = 1'b0;  addr_rom[20981]='h000007d4;  wr_data_rom[20981]='h00000000;
    rd_cycle[20982] = 1'b1;  wr_cycle[20982] = 1'b0;  addr_rom[20982]='h000007d8;  wr_data_rom[20982]='h00000000;
    rd_cycle[20983] = 1'b1;  wr_cycle[20983] = 1'b0;  addr_rom[20983]='h000007dc;  wr_data_rom[20983]='h00000000;
    rd_cycle[20984] = 1'b1;  wr_cycle[20984] = 1'b0;  addr_rom[20984]='h000007e0;  wr_data_rom[20984]='h00000000;
    rd_cycle[20985] = 1'b1;  wr_cycle[20985] = 1'b0;  addr_rom[20985]='h000007e4;  wr_data_rom[20985]='h00000000;
    rd_cycle[20986] = 1'b1;  wr_cycle[20986] = 1'b0;  addr_rom[20986]='h000007e8;  wr_data_rom[20986]='h00000000;
    rd_cycle[20987] = 1'b1;  wr_cycle[20987] = 1'b0;  addr_rom[20987]='h000007ec;  wr_data_rom[20987]='h00000000;
    rd_cycle[20988] = 1'b1;  wr_cycle[20988] = 1'b0;  addr_rom[20988]='h000007f0;  wr_data_rom[20988]='h00000000;
    rd_cycle[20989] = 1'b1;  wr_cycle[20989] = 1'b0;  addr_rom[20989]='h000007f4;  wr_data_rom[20989]='h00000000;
    rd_cycle[20990] = 1'b1;  wr_cycle[20990] = 1'b0;  addr_rom[20990]='h000007f8;  wr_data_rom[20990]='h00000000;
    rd_cycle[20991] = 1'b1;  wr_cycle[20991] = 1'b0;  addr_rom[20991]='h000007fc;  wr_data_rom[20991]='h00000000;
    rd_cycle[20992] = 1'b1;  wr_cycle[20992] = 1'b0;  addr_rom[20992]='h00000800;  wr_data_rom[20992]='h00000000;
    rd_cycle[20993] = 1'b1;  wr_cycle[20993] = 1'b0;  addr_rom[20993]='h00000804;  wr_data_rom[20993]='h00000000;
    rd_cycle[20994] = 1'b1;  wr_cycle[20994] = 1'b0;  addr_rom[20994]='h00000808;  wr_data_rom[20994]='h00000000;
    rd_cycle[20995] = 1'b1;  wr_cycle[20995] = 1'b0;  addr_rom[20995]='h0000080c;  wr_data_rom[20995]='h00000000;
    rd_cycle[20996] = 1'b1;  wr_cycle[20996] = 1'b0;  addr_rom[20996]='h00000810;  wr_data_rom[20996]='h00000000;
    rd_cycle[20997] = 1'b1;  wr_cycle[20997] = 1'b0;  addr_rom[20997]='h00000814;  wr_data_rom[20997]='h00000000;
    rd_cycle[20998] = 1'b1;  wr_cycle[20998] = 1'b0;  addr_rom[20998]='h00000818;  wr_data_rom[20998]='h00000000;
    rd_cycle[20999] = 1'b1;  wr_cycle[20999] = 1'b0;  addr_rom[20999]='h0000081c;  wr_data_rom[20999]='h00000000;
    rd_cycle[21000] = 1'b1;  wr_cycle[21000] = 1'b0;  addr_rom[21000]='h00000820;  wr_data_rom[21000]='h00000000;
    rd_cycle[21001] = 1'b1;  wr_cycle[21001] = 1'b0;  addr_rom[21001]='h00000824;  wr_data_rom[21001]='h00000000;
    rd_cycle[21002] = 1'b1;  wr_cycle[21002] = 1'b0;  addr_rom[21002]='h00000828;  wr_data_rom[21002]='h00000000;
    rd_cycle[21003] = 1'b1;  wr_cycle[21003] = 1'b0;  addr_rom[21003]='h0000082c;  wr_data_rom[21003]='h00000000;
    rd_cycle[21004] = 1'b1;  wr_cycle[21004] = 1'b0;  addr_rom[21004]='h00000830;  wr_data_rom[21004]='h00000000;
    rd_cycle[21005] = 1'b1;  wr_cycle[21005] = 1'b0;  addr_rom[21005]='h00000834;  wr_data_rom[21005]='h00000000;
    rd_cycle[21006] = 1'b1;  wr_cycle[21006] = 1'b0;  addr_rom[21006]='h00000838;  wr_data_rom[21006]='h00000000;
    rd_cycle[21007] = 1'b1;  wr_cycle[21007] = 1'b0;  addr_rom[21007]='h0000083c;  wr_data_rom[21007]='h00000000;
    rd_cycle[21008] = 1'b1;  wr_cycle[21008] = 1'b0;  addr_rom[21008]='h00000840;  wr_data_rom[21008]='h00000000;
    rd_cycle[21009] = 1'b1;  wr_cycle[21009] = 1'b0;  addr_rom[21009]='h00000844;  wr_data_rom[21009]='h00000000;
    rd_cycle[21010] = 1'b1;  wr_cycle[21010] = 1'b0;  addr_rom[21010]='h00000848;  wr_data_rom[21010]='h00000000;
    rd_cycle[21011] = 1'b1;  wr_cycle[21011] = 1'b0;  addr_rom[21011]='h0000084c;  wr_data_rom[21011]='h00000000;
    rd_cycle[21012] = 1'b1;  wr_cycle[21012] = 1'b0;  addr_rom[21012]='h00000850;  wr_data_rom[21012]='h00000000;
    rd_cycle[21013] = 1'b1;  wr_cycle[21013] = 1'b0;  addr_rom[21013]='h00000854;  wr_data_rom[21013]='h00000000;
    rd_cycle[21014] = 1'b1;  wr_cycle[21014] = 1'b0;  addr_rom[21014]='h00000858;  wr_data_rom[21014]='h00000000;
    rd_cycle[21015] = 1'b1;  wr_cycle[21015] = 1'b0;  addr_rom[21015]='h0000085c;  wr_data_rom[21015]='h00000000;
    rd_cycle[21016] = 1'b1;  wr_cycle[21016] = 1'b0;  addr_rom[21016]='h00000860;  wr_data_rom[21016]='h00000000;
    rd_cycle[21017] = 1'b1;  wr_cycle[21017] = 1'b0;  addr_rom[21017]='h00000864;  wr_data_rom[21017]='h00000000;
    rd_cycle[21018] = 1'b1;  wr_cycle[21018] = 1'b0;  addr_rom[21018]='h00000868;  wr_data_rom[21018]='h00000000;
    rd_cycle[21019] = 1'b1;  wr_cycle[21019] = 1'b0;  addr_rom[21019]='h0000086c;  wr_data_rom[21019]='h00000000;
    rd_cycle[21020] = 1'b1;  wr_cycle[21020] = 1'b0;  addr_rom[21020]='h00000870;  wr_data_rom[21020]='h00000000;
    rd_cycle[21021] = 1'b1;  wr_cycle[21021] = 1'b0;  addr_rom[21021]='h00000874;  wr_data_rom[21021]='h00000000;
    rd_cycle[21022] = 1'b1;  wr_cycle[21022] = 1'b0;  addr_rom[21022]='h00000878;  wr_data_rom[21022]='h00000000;
    rd_cycle[21023] = 1'b1;  wr_cycle[21023] = 1'b0;  addr_rom[21023]='h0000087c;  wr_data_rom[21023]='h00000000;
    rd_cycle[21024] = 1'b1;  wr_cycle[21024] = 1'b0;  addr_rom[21024]='h00000880;  wr_data_rom[21024]='h00000000;
    rd_cycle[21025] = 1'b1;  wr_cycle[21025] = 1'b0;  addr_rom[21025]='h00000884;  wr_data_rom[21025]='h00000000;
    rd_cycle[21026] = 1'b1;  wr_cycle[21026] = 1'b0;  addr_rom[21026]='h00000888;  wr_data_rom[21026]='h00000000;
    rd_cycle[21027] = 1'b1;  wr_cycle[21027] = 1'b0;  addr_rom[21027]='h0000088c;  wr_data_rom[21027]='h00000000;
    rd_cycle[21028] = 1'b1;  wr_cycle[21028] = 1'b0;  addr_rom[21028]='h00000890;  wr_data_rom[21028]='h00000000;
    rd_cycle[21029] = 1'b1;  wr_cycle[21029] = 1'b0;  addr_rom[21029]='h00000894;  wr_data_rom[21029]='h00000000;
    rd_cycle[21030] = 1'b1;  wr_cycle[21030] = 1'b0;  addr_rom[21030]='h00000898;  wr_data_rom[21030]='h00000000;
    rd_cycle[21031] = 1'b1;  wr_cycle[21031] = 1'b0;  addr_rom[21031]='h0000089c;  wr_data_rom[21031]='h00000000;
    rd_cycle[21032] = 1'b1;  wr_cycle[21032] = 1'b0;  addr_rom[21032]='h000008a0;  wr_data_rom[21032]='h00000000;
    rd_cycle[21033] = 1'b1;  wr_cycle[21033] = 1'b0;  addr_rom[21033]='h000008a4;  wr_data_rom[21033]='h00000000;
    rd_cycle[21034] = 1'b1;  wr_cycle[21034] = 1'b0;  addr_rom[21034]='h000008a8;  wr_data_rom[21034]='h00000000;
    rd_cycle[21035] = 1'b1;  wr_cycle[21035] = 1'b0;  addr_rom[21035]='h000008ac;  wr_data_rom[21035]='h00000000;
    rd_cycle[21036] = 1'b1;  wr_cycle[21036] = 1'b0;  addr_rom[21036]='h000008b0;  wr_data_rom[21036]='h00000000;
    rd_cycle[21037] = 1'b1;  wr_cycle[21037] = 1'b0;  addr_rom[21037]='h000008b4;  wr_data_rom[21037]='h00000000;
    rd_cycle[21038] = 1'b1;  wr_cycle[21038] = 1'b0;  addr_rom[21038]='h000008b8;  wr_data_rom[21038]='h00000000;
    rd_cycle[21039] = 1'b1;  wr_cycle[21039] = 1'b0;  addr_rom[21039]='h000008bc;  wr_data_rom[21039]='h00000000;
    rd_cycle[21040] = 1'b1;  wr_cycle[21040] = 1'b0;  addr_rom[21040]='h000008c0;  wr_data_rom[21040]='h00000000;
    rd_cycle[21041] = 1'b1;  wr_cycle[21041] = 1'b0;  addr_rom[21041]='h000008c4;  wr_data_rom[21041]='h00000000;
    rd_cycle[21042] = 1'b1;  wr_cycle[21042] = 1'b0;  addr_rom[21042]='h000008c8;  wr_data_rom[21042]='h00000000;
    rd_cycle[21043] = 1'b1;  wr_cycle[21043] = 1'b0;  addr_rom[21043]='h000008cc;  wr_data_rom[21043]='h00000000;
    rd_cycle[21044] = 1'b1;  wr_cycle[21044] = 1'b0;  addr_rom[21044]='h000008d0;  wr_data_rom[21044]='h00000000;
    rd_cycle[21045] = 1'b1;  wr_cycle[21045] = 1'b0;  addr_rom[21045]='h000008d4;  wr_data_rom[21045]='h00000000;
    rd_cycle[21046] = 1'b1;  wr_cycle[21046] = 1'b0;  addr_rom[21046]='h000008d8;  wr_data_rom[21046]='h00000000;
    rd_cycle[21047] = 1'b1;  wr_cycle[21047] = 1'b0;  addr_rom[21047]='h000008dc;  wr_data_rom[21047]='h00000000;
    rd_cycle[21048] = 1'b1;  wr_cycle[21048] = 1'b0;  addr_rom[21048]='h000008e0;  wr_data_rom[21048]='h00000000;
    rd_cycle[21049] = 1'b1;  wr_cycle[21049] = 1'b0;  addr_rom[21049]='h000008e4;  wr_data_rom[21049]='h00000000;
    rd_cycle[21050] = 1'b1;  wr_cycle[21050] = 1'b0;  addr_rom[21050]='h000008e8;  wr_data_rom[21050]='h00000000;
    rd_cycle[21051] = 1'b1;  wr_cycle[21051] = 1'b0;  addr_rom[21051]='h000008ec;  wr_data_rom[21051]='h00000000;
    rd_cycle[21052] = 1'b1;  wr_cycle[21052] = 1'b0;  addr_rom[21052]='h000008f0;  wr_data_rom[21052]='h00000000;
    rd_cycle[21053] = 1'b1;  wr_cycle[21053] = 1'b0;  addr_rom[21053]='h000008f4;  wr_data_rom[21053]='h00000000;
    rd_cycle[21054] = 1'b1;  wr_cycle[21054] = 1'b0;  addr_rom[21054]='h000008f8;  wr_data_rom[21054]='h00000000;
    rd_cycle[21055] = 1'b1;  wr_cycle[21055] = 1'b0;  addr_rom[21055]='h000008fc;  wr_data_rom[21055]='h00000000;
    rd_cycle[21056] = 1'b1;  wr_cycle[21056] = 1'b0;  addr_rom[21056]='h00000900;  wr_data_rom[21056]='h00000000;
    rd_cycle[21057] = 1'b1;  wr_cycle[21057] = 1'b0;  addr_rom[21057]='h00000904;  wr_data_rom[21057]='h00000000;
    rd_cycle[21058] = 1'b1;  wr_cycle[21058] = 1'b0;  addr_rom[21058]='h00000908;  wr_data_rom[21058]='h00000000;
    rd_cycle[21059] = 1'b1;  wr_cycle[21059] = 1'b0;  addr_rom[21059]='h0000090c;  wr_data_rom[21059]='h00000000;
    rd_cycle[21060] = 1'b1;  wr_cycle[21060] = 1'b0;  addr_rom[21060]='h00000910;  wr_data_rom[21060]='h00000000;
    rd_cycle[21061] = 1'b1;  wr_cycle[21061] = 1'b0;  addr_rom[21061]='h00000914;  wr_data_rom[21061]='h00000000;
    rd_cycle[21062] = 1'b1;  wr_cycle[21062] = 1'b0;  addr_rom[21062]='h00000918;  wr_data_rom[21062]='h00000000;
    rd_cycle[21063] = 1'b1;  wr_cycle[21063] = 1'b0;  addr_rom[21063]='h0000091c;  wr_data_rom[21063]='h00000000;
    rd_cycle[21064] = 1'b1;  wr_cycle[21064] = 1'b0;  addr_rom[21064]='h00000920;  wr_data_rom[21064]='h00000000;
    rd_cycle[21065] = 1'b1;  wr_cycle[21065] = 1'b0;  addr_rom[21065]='h00000924;  wr_data_rom[21065]='h00000000;
    rd_cycle[21066] = 1'b1;  wr_cycle[21066] = 1'b0;  addr_rom[21066]='h00000928;  wr_data_rom[21066]='h00000000;
    rd_cycle[21067] = 1'b1;  wr_cycle[21067] = 1'b0;  addr_rom[21067]='h0000092c;  wr_data_rom[21067]='h00000000;
    rd_cycle[21068] = 1'b1;  wr_cycle[21068] = 1'b0;  addr_rom[21068]='h00000930;  wr_data_rom[21068]='h00000000;
    rd_cycle[21069] = 1'b1;  wr_cycle[21069] = 1'b0;  addr_rom[21069]='h00000934;  wr_data_rom[21069]='h00000000;
    rd_cycle[21070] = 1'b1;  wr_cycle[21070] = 1'b0;  addr_rom[21070]='h00000938;  wr_data_rom[21070]='h00000000;
    rd_cycle[21071] = 1'b1;  wr_cycle[21071] = 1'b0;  addr_rom[21071]='h0000093c;  wr_data_rom[21071]='h00000000;
    rd_cycle[21072] = 1'b1;  wr_cycle[21072] = 1'b0;  addr_rom[21072]='h00000940;  wr_data_rom[21072]='h00000000;
    rd_cycle[21073] = 1'b1;  wr_cycle[21073] = 1'b0;  addr_rom[21073]='h00000944;  wr_data_rom[21073]='h00000000;
    rd_cycle[21074] = 1'b1;  wr_cycle[21074] = 1'b0;  addr_rom[21074]='h00000948;  wr_data_rom[21074]='h00000000;
    rd_cycle[21075] = 1'b1;  wr_cycle[21075] = 1'b0;  addr_rom[21075]='h0000094c;  wr_data_rom[21075]='h00000000;
    rd_cycle[21076] = 1'b1;  wr_cycle[21076] = 1'b0;  addr_rom[21076]='h00000950;  wr_data_rom[21076]='h00000000;
    rd_cycle[21077] = 1'b1;  wr_cycle[21077] = 1'b0;  addr_rom[21077]='h00000954;  wr_data_rom[21077]='h00000000;
    rd_cycle[21078] = 1'b1;  wr_cycle[21078] = 1'b0;  addr_rom[21078]='h00000958;  wr_data_rom[21078]='h00000000;
    rd_cycle[21079] = 1'b1;  wr_cycle[21079] = 1'b0;  addr_rom[21079]='h0000095c;  wr_data_rom[21079]='h00000000;
    rd_cycle[21080] = 1'b1;  wr_cycle[21080] = 1'b0;  addr_rom[21080]='h00000960;  wr_data_rom[21080]='h00000000;
    rd_cycle[21081] = 1'b1;  wr_cycle[21081] = 1'b0;  addr_rom[21081]='h00000964;  wr_data_rom[21081]='h00000000;
    rd_cycle[21082] = 1'b1;  wr_cycle[21082] = 1'b0;  addr_rom[21082]='h00000968;  wr_data_rom[21082]='h00000000;
    rd_cycle[21083] = 1'b1;  wr_cycle[21083] = 1'b0;  addr_rom[21083]='h0000096c;  wr_data_rom[21083]='h00000000;
    rd_cycle[21084] = 1'b1;  wr_cycle[21084] = 1'b0;  addr_rom[21084]='h00000970;  wr_data_rom[21084]='h00000000;
    rd_cycle[21085] = 1'b1;  wr_cycle[21085] = 1'b0;  addr_rom[21085]='h00000974;  wr_data_rom[21085]='h00000000;
    rd_cycle[21086] = 1'b1;  wr_cycle[21086] = 1'b0;  addr_rom[21086]='h00000978;  wr_data_rom[21086]='h00000000;
    rd_cycle[21087] = 1'b1;  wr_cycle[21087] = 1'b0;  addr_rom[21087]='h0000097c;  wr_data_rom[21087]='h00000000;
    rd_cycle[21088] = 1'b1;  wr_cycle[21088] = 1'b0;  addr_rom[21088]='h00000980;  wr_data_rom[21088]='h00000000;
    rd_cycle[21089] = 1'b1;  wr_cycle[21089] = 1'b0;  addr_rom[21089]='h00000984;  wr_data_rom[21089]='h00000000;
    rd_cycle[21090] = 1'b1;  wr_cycle[21090] = 1'b0;  addr_rom[21090]='h00000988;  wr_data_rom[21090]='h00000000;
    rd_cycle[21091] = 1'b1;  wr_cycle[21091] = 1'b0;  addr_rom[21091]='h0000098c;  wr_data_rom[21091]='h00000000;
    rd_cycle[21092] = 1'b1;  wr_cycle[21092] = 1'b0;  addr_rom[21092]='h00000990;  wr_data_rom[21092]='h00000000;
    rd_cycle[21093] = 1'b1;  wr_cycle[21093] = 1'b0;  addr_rom[21093]='h00000994;  wr_data_rom[21093]='h00000000;
    rd_cycle[21094] = 1'b1;  wr_cycle[21094] = 1'b0;  addr_rom[21094]='h00000998;  wr_data_rom[21094]='h00000000;
    rd_cycle[21095] = 1'b1;  wr_cycle[21095] = 1'b0;  addr_rom[21095]='h0000099c;  wr_data_rom[21095]='h00000000;
    rd_cycle[21096] = 1'b1;  wr_cycle[21096] = 1'b0;  addr_rom[21096]='h000009a0;  wr_data_rom[21096]='h00000000;
    rd_cycle[21097] = 1'b1;  wr_cycle[21097] = 1'b0;  addr_rom[21097]='h000009a4;  wr_data_rom[21097]='h00000000;
    rd_cycle[21098] = 1'b1;  wr_cycle[21098] = 1'b0;  addr_rom[21098]='h000009a8;  wr_data_rom[21098]='h00000000;
    rd_cycle[21099] = 1'b1;  wr_cycle[21099] = 1'b0;  addr_rom[21099]='h000009ac;  wr_data_rom[21099]='h00000000;
    rd_cycle[21100] = 1'b1;  wr_cycle[21100] = 1'b0;  addr_rom[21100]='h000009b0;  wr_data_rom[21100]='h00000000;
    rd_cycle[21101] = 1'b1;  wr_cycle[21101] = 1'b0;  addr_rom[21101]='h000009b4;  wr_data_rom[21101]='h00000000;
    rd_cycle[21102] = 1'b1;  wr_cycle[21102] = 1'b0;  addr_rom[21102]='h000009b8;  wr_data_rom[21102]='h00000000;
    rd_cycle[21103] = 1'b1;  wr_cycle[21103] = 1'b0;  addr_rom[21103]='h000009bc;  wr_data_rom[21103]='h00000000;
    rd_cycle[21104] = 1'b1;  wr_cycle[21104] = 1'b0;  addr_rom[21104]='h000009c0;  wr_data_rom[21104]='h00000000;
    rd_cycle[21105] = 1'b1;  wr_cycle[21105] = 1'b0;  addr_rom[21105]='h000009c4;  wr_data_rom[21105]='h00000000;
    rd_cycle[21106] = 1'b1;  wr_cycle[21106] = 1'b0;  addr_rom[21106]='h000009c8;  wr_data_rom[21106]='h00000000;
    rd_cycle[21107] = 1'b1;  wr_cycle[21107] = 1'b0;  addr_rom[21107]='h000009cc;  wr_data_rom[21107]='h00000000;
    rd_cycle[21108] = 1'b1;  wr_cycle[21108] = 1'b0;  addr_rom[21108]='h000009d0;  wr_data_rom[21108]='h00000000;
    rd_cycle[21109] = 1'b1;  wr_cycle[21109] = 1'b0;  addr_rom[21109]='h000009d4;  wr_data_rom[21109]='h00000000;
    rd_cycle[21110] = 1'b1;  wr_cycle[21110] = 1'b0;  addr_rom[21110]='h000009d8;  wr_data_rom[21110]='h00000000;
    rd_cycle[21111] = 1'b1;  wr_cycle[21111] = 1'b0;  addr_rom[21111]='h000009dc;  wr_data_rom[21111]='h00000000;
    rd_cycle[21112] = 1'b1;  wr_cycle[21112] = 1'b0;  addr_rom[21112]='h000009e0;  wr_data_rom[21112]='h00000000;
    rd_cycle[21113] = 1'b1;  wr_cycle[21113] = 1'b0;  addr_rom[21113]='h000009e4;  wr_data_rom[21113]='h00000000;
    rd_cycle[21114] = 1'b1;  wr_cycle[21114] = 1'b0;  addr_rom[21114]='h000009e8;  wr_data_rom[21114]='h00000000;
    rd_cycle[21115] = 1'b1;  wr_cycle[21115] = 1'b0;  addr_rom[21115]='h000009ec;  wr_data_rom[21115]='h00000000;
    rd_cycle[21116] = 1'b1;  wr_cycle[21116] = 1'b0;  addr_rom[21116]='h000009f0;  wr_data_rom[21116]='h00000000;
    rd_cycle[21117] = 1'b1;  wr_cycle[21117] = 1'b0;  addr_rom[21117]='h000009f4;  wr_data_rom[21117]='h00000000;
    rd_cycle[21118] = 1'b1;  wr_cycle[21118] = 1'b0;  addr_rom[21118]='h000009f8;  wr_data_rom[21118]='h00000000;
    rd_cycle[21119] = 1'b1;  wr_cycle[21119] = 1'b0;  addr_rom[21119]='h000009fc;  wr_data_rom[21119]='h00000000;
    rd_cycle[21120] = 1'b1;  wr_cycle[21120] = 1'b0;  addr_rom[21120]='h00000a00;  wr_data_rom[21120]='h00000000;
    rd_cycle[21121] = 1'b1;  wr_cycle[21121] = 1'b0;  addr_rom[21121]='h00000a04;  wr_data_rom[21121]='h00000000;
    rd_cycle[21122] = 1'b1;  wr_cycle[21122] = 1'b0;  addr_rom[21122]='h00000a08;  wr_data_rom[21122]='h00000000;
    rd_cycle[21123] = 1'b1;  wr_cycle[21123] = 1'b0;  addr_rom[21123]='h00000a0c;  wr_data_rom[21123]='h00000000;
    rd_cycle[21124] = 1'b1;  wr_cycle[21124] = 1'b0;  addr_rom[21124]='h00000a10;  wr_data_rom[21124]='h00000000;
    rd_cycle[21125] = 1'b1;  wr_cycle[21125] = 1'b0;  addr_rom[21125]='h00000a14;  wr_data_rom[21125]='h00000000;
    rd_cycle[21126] = 1'b1;  wr_cycle[21126] = 1'b0;  addr_rom[21126]='h00000a18;  wr_data_rom[21126]='h00000000;
    rd_cycle[21127] = 1'b1;  wr_cycle[21127] = 1'b0;  addr_rom[21127]='h00000a1c;  wr_data_rom[21127]='h00000000;
    rd_cycle[21128] = 1'b1;  wr_cycle[21128] = 1'b0;  addr_rom[21128]='h00000a20;  wr_data_rom[21128]='h00000000;
    rd_cycle[21129] = 1'b1;  wr_cycle[21129] = 1'b0;  addr_rom[21129]='h00000a24;  wr_data_rom[21129]='h00000000;
    rd_cycle[21130] = 1'b1;  wr_cycle[21130] = 1'b0;  addr_rom[21130]='h00000a28;  wr_data_rom[21130]='h00000000;
    rd_cycle[21131] = 1'b1;  wr_cycle[21131] = 1'b0;  addr_rom[21131]='h00000a2c;  wr_data_rom[21131]='h00000000;
    rd_cycle[21132] = 1'b1;  wr_cycle[21132] = 1'b0;  addr_rom[21132]='h00000a30;  wr_data_rom[21132]='h00000000;
    rd_cycle[21133] = 1'b1;  wr_cycle[21133] = 1'b0;  addr_rom[21133]='h00000a34;  wr_data_rom[21133]='h00000000;
    rd_cycle[21134] = 1'b1;  wr_cycle[21134] = 1'b0;  addr_rom[21134]='h00000a38;  wr_data_rom[21134]='h00000000;
    rd_cycle[21135] = 1'b1;  wr_cycle[21135] = 1'b0;  addr_rom[21135]='h00000a3c;  wr_data_rom[21135]='h00000000;
    rd_cycle[21136] = 1'b1;  wr_cycle[21136] = 1'b0;  addr_rom[21136]='h00000a40;  wr_data_rom[21136]='h00000000;
    rd_cycle[21137] = 1'b1;  wr_cycle[21137] = 1'b0;  addr_rom[21137]='h00000a44;  wr_data_rom[21137]='h00000000;
    rd_cycle[21138] = 1'b1;  wr_cycle[21138] = 1'b0;  addr_rom[21138]='h00000a48;  wr_data_rom[21138]='h00000000;
    rd_cycle[21139] = 1'b1;  wr_cycle[21139] = 1'b0;  addr_rom[21139]='h00000a4c;  wr_data_rom[21139]='h00000000;
    rd_cycle[21140] = 1'b1;  wr_cycle[21140] = 1'b0;  addr_rom[21140]='h00000a50;  wr_data_rom[21140]='h00000000;
    rd_cycle[21141] = 1'b1;  wr_cycle[21141] = 1'b0;  addr_rom[21141]='h00000a54;  wr_data_rom[21141]='h00000000;
    rd_cycle[21142] = 1'b1;  wr_cycle[21142] = 1'b0;  addr_rom[21142]='h00000a58;  wr_data_rom[21142]='h00000000;
    rd_cycle[21143] = 1'b1;  wr_cycle[21143] = 1'b0;  addr_rom[21143]='h00000a5c;  wr_data_rom[21143]='h00000000;
    rd_cycle[21144] = 1'b1;  wr_cycle[21144] = 1'b0;  addr_rom[21144]='h00000a60;  wr_data_rom[21144]='h00000000;
    rd_cycle[21145] = 1'b1;  wr_cycle[21145] = 1'b0;  addr_rom[21145]='h00000a64;  wr_data_rom[21145]='h00000000;
    rd_cycle[21146] = 1'b1;  wr_cycle[21146] = 1'b0;  addr_rom[21146]='h00000a68;  wr_data_rom[21146]='h00000000;
    rd_cycle[21147] = 1'b1;  wr_cycle[21147] = 1'b0;  addr_rom[21147]='h00000a6c;  wr_data_rom[21147]='h00000000;
    rd_cycle[21148] = 1'b1;  wr_cycle[21148] = 1'b0;  addr_rom[21148]='h00000a70;  wr_data_rom[21148]='h00000000;
    rd_cycle[21149] = 1'b1;  wr_cycle[21149] = 1'b0;  addr_rom[21149]='h00000a74;  wr_data_rom[21149]='h00000000;
    rd_cycle[21150] = 1'b1;  wr_cycle[21150] = 1'b0;  addr_rom[21150]='h00000a78;  wr_data_rom[21150]='h00000000;
    rd_cycle[21151] = 1'b1;  wr_cycle[21151] = 1'b0;  addr_rom[21151]='h00000a7c;  wr_data_rom[21151]='h00000000;
    rd_cycle[21152] = 1'b1;  wr_cycle[21152] = 1'b0;  addr_rom[21152]='h00000a80;  wr_data_rom[21152]='h00000000;
    rd_cycle[21153] = 1'b1;  wr_cycle[21153] = 1'b0;  addr_rom[21153]='h00000a84;  wr_data_rom[21153]='h00000000;
    rd_cycle[21154] = 1'b1;  wr_cycle[21154] = 1'b0;  addr_rom[21154]='h00000a88;  wr_data_rom[21154]='h00000000;
    rd_cycle[21155] = 1'b1;  wr_cycle[21155] = 1'b0;  addr_rom[21155]='h00000a8c;  wr_data_rom[21155]='h00000000;
    rd_cycle[21156] = 1'b1;  wr_cycle[21156] = 1'b0;  addr_rom[21156]='h00000a90;  wr_data_rom[21156]='h00000000;
    rd_cycle[21157] = 1'b1;  wr_cycle[21157] = 1'b0;  addr_rom[21157]='h00000a94;  wr_data_rom[21157]='h00000000;
    rd_cycle[21158] = 1'b1;  wr_cycle[21158] = 1'b0;  addr_rom[21158]='h00000a98;  wr_data_rom[21158]='h00000000;
    rd_cycle[21159] = 1'b1;  wr_cycle[21159] = 1'b0;  addr_rom[21159]='h00000a9c;  wr_data_rom[21159]='h00000000;
    rd_cycle[21160] = 1'b1;  wr_cycle[21160] = 1'b0;  addr_rom[21160]='h00000aa0;  wr_data_rom[21160]='h00000000;
    rd_cycle[21161] = 1'b1;  wr_cycle[21161] = 1'b0;  addr_rom[21161]='h00000aa4;  wr_data_rom[21161]='h00000000;
    rd_cycle[21162] = 1'b1;  wr_cycle[21162] = 1'b0;  addr_rom[21162]='h00000aa8;  wr_data_rom[21162]='h00000000;
    rd_cycle[21163] = 1'b1;  wr_cycle[21163] = 1'b0;  addr_rom[21163]='h00000aac;  wr_data_rom[21163]='h00000000;
    rd_cycle[21164] = 1'b1;  wr_cycle[21164] = 1'b0;  addr_rom[21164]='h00000ab0;  wr_data_rom[21164]='h00000000;
    rd_cycle[21165] = 1'b1;  wr_cycle[21165] = 1'b0;  addr_rom[21165]='h00000ab4;  wr_data_rom[21165]='h00000000;
    rd_cycle[21166] = 1'b1;  wr_cycle[21166] = 1'b0;  addr_rom[21166]='h00000ab8;  wr_data_rom[21166]='h00000000;
    rd_cycle[21167] = 1'b1;  wr_cycle[21167] = 1'b0;  addr_rom[21167]='h00000abc;  wr_data_rom[21167]='h00000000;
    rd_cycle[21168] = 1'b1;  wr_cycle[21168] = 1'b0;  addr_rom[21168]='h00000ac0;  wr_data_rom[21168]='h00000000;
    rd_cycle[21169] = 1'b1;  wr_cycle[21169] = 1'b0;  addr_rom[21169]='h00000ac4;  wr_data_rom[21169]='h00000000;
    rd_cycle[21170] = 1'b1;  wr_cycle[21170] = 1'b0;  addr_rom[21170]='h00000ac8;  wr_data_rom[21170]='h00000000;
    rd_cycle[21171] = 1'b1;  wr_cycle[21171] = 1'b0;  addr_rom[21171]='h00000acc;  wr_data_rom[21171]='h00000000;
    rd_cycle[21172] = 1'b1;  wr_cycle[21172] = 1'b0;  addr_rom[21172]='h00000ad0;  wr_data_rom[21172]='h00000000;
    rd_cycle[21173] = 1'b1;  wr_cycle[21173] = 1'b0;  addr_rom[21173]='h00000ad4;  wr_data_rom[21173]='h00000000;
    rd_cycle[21174] = 1'b1;  wr_cycle[21174] = 1'b0;  addr_rom[21174]='h00000ad8;  wr_data_rom[21174]='h00000000;
    rd_cycle[21175] = 1'b1;  wr_cycle[21175] = 1'b0;  addr_rom[21175]='h00000adc;  wr_data_rom[21175]='h00000000;
    rd_cycle[21176] = 1'b1;  wr_cycle[21176] = 1'b0;  addr_rom[21176]='h00000ae0;  wr_data_rom[21176]='h00000000;
    rd_cycle[21177] = 1'b1;  wr_cycle[21177] = 1'b0;  addr_rom[21177]='h00000ae4;  wr_data_rom[21177]='h00000000;
    rd_cycle[21178] = 1'b1;  wr_cycle[21178] = 1'b0;  addr_rom[21178]='h00000ae8;  wr_data_rom[21178]='h00000000;
    rd_cycle[21179] = 1'b1;  wr_cycle[21179] = 1'b0;  addr_rom[21179]='h00000aec;  wr_data_rom[21179]='h00000000;
    rd_cycle[21180] = 1'b1;  wr_cycle[21180] = 1'b0;  addr_rom[21180]='h00000af0;  wr_data_rom[21180]='h00000000;
    rd_cycle[21181] = 1'b1;  wr_cycle[21181] = 1'b0;  addr_rom[21181]='h00000af4;  wr_data_rom[21181]='h00000000;
    rd_cycle[21182] = 1'b1;  wr_cycle[21182] = 1'b0;  addr_rom[21182]='h00000af8;  wr_data_rom[21182]='h00000000;
    rd_cycle[21183] = 1'b1;  wr_cycle[21183] = 1'b0;  addr_rom[21183]='h00000afc;  wr_data_rom[21183]='h00000000;
    rd_cycle[21184] = 1'b1;  wr_cycle[21184] = 1'b0;  addr_rom[21184]='h00000b00;  wr_data_rom[21184]='h00000000;
    rd_cycle[21185] = 1'b1;  wr_cycle[21185] = 1'b0;  addr_rom[21185]='h00000b04;  wr_data_rom[21185]='h00000000;
    rd_cycle[21186] = 1'b1;  wr_cycle[21186] = 1'b0;  addr_rom[21186]='h00000b08;  wr_data_rom[21186]='h00000000;
    rd_cycle[21187] = 1'b1;  wr_cycle[21187] = 1'b0;  addr_rom[21187]='h00000b0c;  wr_data_rom[21187]='h00000000;
    rd_cycle[21188] = 1'b1;  wr_cycle[21188] = 1'b0;  addr_rom[21188]='h00000b10;  wr_data_rom[21188]='h00000000;
    rd_cycle[21189] = 1'b1;  wr_cycle[21189] = 1'b0;  addr_rom[21189]='h00000b14;  wr_data_rom[21189]='h00000000;
    rd_cycle[21190] = 1'b1;  wr_cycle[21190] = 1'b0;  addr_rom[21190]='h00000b18;  wr_data_rom[21190]='h00000000;
    rd_cycle[21191] = 1'b1;  wr_cycle[21191] = 1'b0;  addr_rom[21191]='h00000b1c;  wr_data_rom[21191]='h00000000;
    rd_cycle[21192] = 1'b1;  wr_cycle[21192] = 1'b0;  addr_rom[21192]='h00000b20;  wr_data_rom[21192]='h00000000;
    rd_cycle[21193] = 1'b1;  wr_cycle[21193] = 1'b0;  addr_rom[21193]='h00000b24;  wr_data_rom[21193]='h00000000;
    rd_cycle[21194] = 1'b1;  wr_cycle[21194] = 1'b0;  addr_rom[21194]='h00000b28;  wr_data_rom[21194]='h00000000;
    rd_cycle[21195] = 1'b1;  wr_cycle[21195] = 1'b0;  addr_rom[21195]='h00000b2c;  wr_data_rom[21195]='h00000000;
    rd_cycle[21196] = 1'b1;  wr_cycle[21196] = 1'b0;  addr_rom[21196]='h00000b30;  wr_data_rom[21196]='h00000000;
    rd_cycle[21197] = 1'b1;  wr_cycle[21197] = 1'b0;  addr_rom[21197]='h00000b34;  wr_data_rom[21197]='h00000000;
    rd_cycle[21198] = 1'b1;  wr_cycle[21198] = 1'b0;  addr_rom[21198]='h00000b38;  wr_data_rom[21198]='h00000000;
    rd_cycle[21199] = 1'b1;  wr_cycle[21199] = 1'b0;  addr_rom[21199]='h00000b3c;  wr_data_rom[21199]='h00000000;
    rd_cycle[21200] = 1'b1;  wr_cycle[21200] = 1'b0;  addr_rom[21200]='h00000b40;  wr_data_rom[21200]='h00000000;
    rd_cycle[21201] = 1'b1;  wr_cycle[21201] = 1'b0;  addr_rom[21201]='h00000b44;  wr_data_rom[21201]='h00000000;
    rd_cycle[21202] = 1'b1;  wr_cycle[21202] = 1'b0;  addr_rom[21202]='h00000b48;  wr_data_rom[21202]='h00000000;
    rd_cycle[21203] = 1'b1;  wr_cycle[21203] = 1'b0;  addr_rom[21203]='h00000b4c;  wr_data_rom[21203]='h00000000;
    rd_cycle[21204] = 1'b1;  wr_cycle[21204] = 1'b0;  addr_rom[21204]='h00000b50;  wr_data_rom[21204]='h00000000;
    rd_cycle[21205] = 1'b1;  wr_cycle[21205] = 1'b0;  addr_rom[21205]='h00000b54;  wr_data_rom[21205]='h00000000;
    rd_cycle[21206] = 1'b1;  wr_cycle[21206] = 1'b0;  addr_rom[21206]='h00000b58;  wr_data_rom[21206]='h00000000;
    rd_cycle[21207] = 1'b1;  wr_cycle[21207] = 1'b0;  addr_rom[21207]='h00000b5c;  wr_data_rom[21207]='h00000000;
    rd_cycle[21208] = 1'b1;  wr_cycle[21208] = 1'b0;  addr_rom[21208]='h00000b60;  wr_data_rom[21208]='h00000000;
    rd_cycle[21209] = 1'b1;  wr_cycle[21209] = 1'b0;  addr_rom[21209]='h00000b64;  wr_data_rom[21209]='h00000000;
    rd_cycle[21210] = 1'b1;  wr_cycle[21210] = 1'b0;  addr_rom[21210]='h00000b68;  wr_data_rom[21210]='h00000000;
    rd_cycle[21211] = 1'b1;  wr_cycle[21211] = 1'b0;  addr_rom[21211]='h00000b6c;  wr_data_rom[21211]='h00000000;
    rd_cycle[21212] = 1'b1;  wr_cycle[21212] = 1'b0;  addr_rom[21212]='h00000b70;  wr_data_rom[21212]='h00000000;
    rd_cycle[21213] = 1'b1;  wr_cycle[21213] = 1'b0;  addr_rom[21213]='h00000b74;  wr_data_rom[21213]='h00000000;
    rd_cycle[21214] = 1'b1;  wr_cycle[21214] = 1'b0;  addr_rom[21214]='h00000b78;  wr_data_rom[21214]='h00000000;
    rd_cycle[21215] = 1'b1;  wr_cycle[21215] = 1'b0;  addr_rom[21215]='h00000b7c;  wr_data_rom[21215]='h00000000;
    rd_cycle[21216] = 1'b1;  wr_cycle[21216] = 1'b0;  addr_rom[21216]='h00000b80;  wr_data_rom[21216]='h00000000;
    rd_cycle[21217] = 1'b1;  wr_cycle[21217] = 1'b0;  addr_rom[21217]='h00000b84;  wr_data_rom[21217]='h00000000;
    rd_cycle[21218] = 1'b1;  wr_cycle[21218] = 1'b0;  addr_rom[21218]='h00000b88;  wr_data_rom[21218]='h00000000;
    rd_cycle[21219] = 1'b1;  wr_cycle[21219] = 1'b0;  addr_rom[21219]='h00000b8c;  wr_data_rom[21219]='h00000000;
    rd_cycle[21220] = 1'b1;  wr_cycle[21220] = 1'b0;  addr_rom[21220]='h00000b90;  wr_data_rom[21220]='h00000000;
    rd_cycle[21221] = 1'b1;  wr_cycle[21221] = 1'b0;  addr_rom[21221]='h00000b94;  wr_data_rom[21221]='h00000000;
    rd_cycle[21222] = 1'b1;  wr_cycle[21222] = 1'b0;  addr_rom[21222]='h00000b98;  wr_data_rom[21222]='h00000000;
    rd_cycle[21223] = 1'b1;  wr_cycle[21223] = 1'b0;  addr_rom[21223]='h00000b9c;  wr_data_rom[21223]='h00000000;
    rd_cycle[21224] = 1'b1;  wr_cycle[21224] = 1'b0;  addr_rom[21224]='h00000ba0;  wr_data_rom[21224]='h00000000;
    rd_cycle[21225] = 1'b1;  wr_cycle[21225] = 1'b0;  addr_rom[21225]='h00000ba4;  wr_data_rom[21225]='h00000000;
    rd_cycle[21226] = 1'b1;  wr_cycle[21226] = 1'b0;  addr_rom[21226]='h00000ba8;  wr_data_rom[21226]='h00000000;
    rd_cycle[21227] = 1'b1;  wr_cycle[21227] = 1'b0;  addr_rom[21227]='h00000bac;  wr_data_rom[21227]='h00000000;
    rd_cycle[21228] = 1'b1;  wr_cycle[21228] = 1'b0;  addr_rom[21228]='h00000bb0;  wr_data_rom[21228]='h00000000;
    rd_cycle[21229] = 1'b1;  wr_cycle[21229] = 1'b0;  addr_rom[21229]='h00000bb4;  wr_data_rom[21229]='h00000000;
    rd_cycle[21230] = 1'b1;  wr_cycle[21230] = 1'b0;  addr_rom[21230]='h00000bb8;  wr_data_rom[21230]='h00000000;
    rd_cycle[21231] = 1'b1;  wr_cycle[21231] = 1'b0;  addr_rom[21231]='h00000bbc;  wr_data_rom[21231]='h00000000;
    rd_cycle[21232] = 1'b1;  wr_cycle[21232] = 1'b0;  addr_rom[21232]='h00000bc0;  wr_data_rom[21232]='h00000000;
    rd_cycle[21233] = 1'b1;  wr_cycle[21233] = 1'b0;  addr_rom[21233]='h00000bc4;  wr_data_rom[21233]='h00000000;
    rd_cycle[21234] = 1'b1;  wr_cycle[21234] = 1'b0;  addr_rom[21234]='h00000bc8;  wr_data_rom[21234]='h00000000;
    rd_cycle[21235] = 1'b1;  wr_cycle[21235] = 1'b0;  addr_rom[21235]='h00000bcc;  wr_data_rom[21235]='h00000000;
    rd_cycle[21236] = 1'b1;  wr_cycle[21236] = 1'b0;  addr_rom[21236]='h00000bd0;  wr_data_rom[21236]='h00000000;
    rd_cycle[21237] = 1'b1;  wr_cycle[21237] = 1'b0;  addr_rom[21237]='h00000bd4;  wr_data_rom[21237]='h00000000;
    rd_cycle[21238] = 1'b1;  wr_cycle[21238] = 1'b0;  addr_rom[21238]='h00000bd8;  wr_data_rom[21238]='h00000000;
    rd_cycle[21239] = 1'b1;  wr_cycle[21239] = 1'b0;  addr_rom[21239]='h00000bdc;  wr_data_rom[21239]='h00000000;
    rd_cycle[21240] = 1'b1;  wr_cycle[21240] = 1'b0;  addr_rom[21240]='h00000be0;  wr_data_rom[21240]='h00000000;
    rd_cycle[21241] = 1'b1;  wr_cycle[21241] = 1'b0;  addr_rom[21241]='h00000be4;  wr_data_rom[21241]='h00000000;
    rd_cycle[21242] = 1'b1;  wr_cycle[21242] = 1'b0;  addr_rom[21242]='h00000be8;  wr_data_rom[21242]='h00000000;
    rd_cycle[21243] = 1'b1;  wr_cycle[21243] = 1'b0;  addr_rom[21243]='h00000bec;  wr_data_rom[21243]='h00000000;
    rd_cycle[21244] = 1'b1;  wr_cycle[21244] = 1'b0;  addr_rom[21244]='h00000bf0;  wr_data_rom[21244]='h00000000;
    rd_cycle[21245] = 1'b1;  wr_cycle[21245] = 1'b0;  addr_rom[21245]='h00000bf4;  wr_data_rom[21245]='h00000000;
    rd_cycle[21246] = 1'b1;  wr_cycle[21246] = 1'b0;  addr_rom[21246]='h00000bf8;  wr_data_rom[21246]='h00000000;
    rd_cycle[21247] = 1'b1;  wr_cycle[21247] = 1'b0;  addr_rom[21247]='h00000bfc;  wr_data_rom[21247]='h00000000;
    rd_cycle[21248] = 1'b1;  wr_cycle[21248] = 1'b0;  addr_rom[21248]='h00000c00;  wr_data_rom[21248]='h00000000;
    rd_cycle[21249] = 1'b1;  wr_cycle[21249] = 1'b0;  addr_rom[21249]='h00000c04;  wr_data_rom[21249]='h00000000;
    rd_cycle[21250] = 1'b1;  wr_cycle[21250] = 1'b0;  addr_rom[21250]='h00000c08;  wr_data_rom[21250]='h00000000;
    rd_cycle[21251] = 1'b1;  wr_cycle[21251] = 1'b0;  addr_rom[21251]='h00000c0c;  wr_data_rom[21251]='h00000000;
    rd_cycle[21252] = 1'b1;  wr_cycle[21252] = 1'b0;  addr_rom[21252]='h00000c10;  wr_data_rom[21252]='h00000000;
    rd_cycle[21253] = 1'b1;  wr_cycle[21253] = 1'b0;  addr_rom[21253]='h00000c14;  wr_data_rom[21253]='h00000000;
    rd_cycle[21254] = 1'b1;  wr_cycle[21254] = 1'b0;  addr_rom[21254]='h00000c18;  wr_data_rom[21254]='h00000000;
    rd_cycle[21255] = 1'b1;  wr_cycle[21255] = 1'b0;  addr_rom[21255]='h00000c1c;  wr_data_rom[21255]='h00000000;
    rd_cycle[21256] = 1'b1;  wr_cycle[21256] = 1'b0;  addr_rom[21256]='h00000c20;  wr_data_rom[21256]='h00000000;
    rd_cycle[21257] = 1'b1;  wr_cycle[21257] = 1'b0;  addr_rom[21257]='h00000c24;  wr_data_rom[21257]='h00000000;
    rd_cycle[21258] = 1'b1;  wr_cycle[21258] = 1'b0;  addr_rom[21258]='h00000c28;  wr_data_rom[21258]='h00000000;
    rd_cycle[21259] = 1'b1;  wr_cycle[21259] = 1'b0;  addr_rom[21259]='h00000c2c;  wr_data_rom[21259]='h00000000;
    rd_cycle[21260] = 1'b1;  wr_cycle[21260] = 1'b0;  addr_rom[21260]='h00000c30;  wr_data_rom[21260]='h00000000;
    rd_cycle[21261] = 1'b1;  wr_cycle[21261] = 1'b0;  addr_rom[21261]='h00000c34;  wr_data_rom[21261]='h00000000;
    rd_cycle[21262] = 1'b1;  wr_cycle[21262] = 1'b0;  addr_rom[21262]='h00000c38;  wr_data_rom[21262]='h00000000;
    rd_cycle[21263] = 1'b1;  wr_cycle[21263] = 1'b0;  addr_rom[21263]='h00000c3c;  wr_data_rom[21263]='h00000000;
    rd_cycle[21264] = 1'b1;  wr_cycle[21264] = 1'b0;  addr_rom[21264]='h00000c40;  wr_data_rom[21264]='h00000000;
    rd_cycle[21265] = 1'b1;  wr_cycle[21265] = 1'b0;  addr_rom[21265]='h00000c44;  wr_data_rom[21265]='h00000000;
    rd_cycle[21266] = 1'b1;  wr_cycle[21266] = 1'b0;  addr_rom[21266]='h00000c48;  wr_data_rom[21266]='h00000000;
    rd_cycle[21267] = 1'b1;  wr_cycle[21267] = 1'b0;  addr_rom[21267]='h00000c4c;  wr_data_rom[21267]='h00000000;
    rd_cycle[21268] = 1'b1;  wr_cycle[21268] = 1'b0;  addr_rom[21268]='h00000c50;  wr_data_rom[21268]='h00000000;
    rd_cycle[21269] = 1'b1;  wr_cycle[21269] = 1'b0;  addr_rom[21269]='h00000c54;  wr_data_rom[21269]='h00000000;
    rd_cycle[21270] = 1'b1;  wr_cycle[21270] = 1'b0;  addr_rom[21270]='h00000c58;  wr_data_rom[21270]='h00000000;
    rd_cycle[21271] = 1'b1;  wr_cycle[21271] = 1'b0;  addr_rom[21271]='h00000c5c;  wr_data_rom[21271]='h00000000;
    rd_cycle[21272] = 1'b1;  wr_cycle[21272] = 1'b0;  addr_rom[21272]='h00000c60;  wr_data_rom[21272]='h00000000;
    rd_cycle[21273] = 1'b1;  wr_cycle[21273] = 1'b0;  addr_rom[21273]='h00000c64;  wr_data_rom[21273]='h00000000;
    rd_cycle[21274] = 1'b1;  wr_cycle[21274] = 1'b0;  addr_rom[21274]='h00000c68;  wr_data_rom[21274]='h00000000;
    rd_cycle[21275] = 1'b1;  wr_cycle[21275] = 1'b0;  addr_rom[21275]='h00000c6c;  wr_data_rom[21275]='h00000000;
    rd_cycle[21276] = 1'b1;  wr_cycle[21276] = 1'b0;  addr_rom[21276]='h00000c70;  wr_data_rom[21276]='h00000000;
    rd_cycle[21277] = 1'b1;  wr_cycle[21277] = 1'b0;  addr_rom[21277]='h00000c74;  wr_data_rom[21277]='h00000000;
    rd_cycle[21278] = 1'b1;  wr_cycle[21278] = 1'b0;  addr_rom[21278]='h00000c78;  wr_data_rom[21278]='h00000000;
    rd_cycle[21279] = 1'b1;  wr_cycle[21279] = 1'b0;  addr_rom[21279]='h00000c7c;  wr_data_rom[21279]='h00000000;
    rd_cycle[21280] = 1'b1;  wr_cycle[21280] = 1'b0;  addr_rom[21280]='h00000c80;  wr_data_rom[21280]='h00000000;
    rd_cycle[21281] = 1'b1;  wr_cycle[21281] = 1'b0;  addr_rom[21281]='h00000c84;  wr_data_rom[21281]='h00000000;
    rd_cycle[21282] = 1'b1;  wr_cycle[21282] = 1'b0;  addr_rom[21282]='h00000c88;  wr_data_rom[21282]='h00000000;
    rd_cycle[21283] = 1'b1;  wr_cycle[21283] = 1'b0;  addr_rom[21283]='h00000c8c;  wr_data_rom[21283]='h00000000;
    rd_cycle[21284] = 1'b1;  wr_cycle[21284] = 1'b0;  addr_rom[21284]='h00000c90;  wr_data_rom[21284]='h00000000;
    rd_cycle[21285] = 1'b1;  wr_cycle[21285] = 1'b0;  addr_rom[21285]='h00000c94;  wr_data_rom[21285]='h00000000;
    rd_cycle[21286] = 1'b1;  wr_cycle[21286] = 1'b0;  addr_rom[21286]='h00000c98;  wr_data_rom[21286]='h00000000;
    rd_cycle[21287] = 1'b1;  wr_cycle[21287] = 1'b0;  addr_rom[21287]='h00000c9c;  wr_data_rom[21287]='h00000000;
    rd_cycle[21288] = 1'b1;  wr_cycle[21288] = 1'b0;  addr_rom[21288]='h00000ca0;  wr_data_rom[21288]='h00000000;
    rd_cycle[21289] = 1'b1;  wr_cycle[21289] = 1'b0;  addr_rom[21289]='h00000ca4;  wr_data_rom[21289]='h00000000;
    rd_cycle[21290] = 1'b1;  wr_cycle[21290] = 1'b0;  addr_rom[21290]='h00000ca8;  wr_data_rom[21290]='h00000000;
    rd_cycle[21291] = 1'b1;  wr_cycle[21291] = 1'b0;  addr_rom[21291]='h00000cac;  wr_data_rom[21291]='h00000000;
    rd_cycle[21292] = 1'b1;  wr_cycle[21292] = 1'b0;  addr_rom[21292]='h00000cb0;  wr_data_rom[21292]='h00000000;
    rd_cycle[21293] = 1'b1;  wr_cycle[21293] = 1'b0;  addr_rom[21293]='h00000cb4;  wr_data_rom[21293]='h00000000;
    rd_cycle[21294] = 1'b1;  wr_cycle[21294] = 1'b0;  addr_rom[21294]='h00000cb8;  wr_data_rom[21294]='h00000000;
    rd_cycle[21295] = 1'b1;  wr_cycle[21295] = 1'b0;  addr_rom[21295]='h00000cbc;  wr_data_rom[21295]='h00000000;
    rd_cycle[21296] = 1'b1;  wr_cycle[21296] = 1'b0;  addr_rom[21296]='h00000cc0;  wr_data_rom[21296]='h00000000;
    rd_cycle[21297] = 1'b1;  wr_cycle[21297] = 1'b0;  addr_rom[21297]='h00000cc4;  wr_data_rom[21297]='h00000000;
    rd_cycle[21298] = 1'b1;  wr_cycle[21298] = 1'b0;  addr_rom[21298]='h00000cc8;  wr_data_rom[21298]='h00000000;
    rd_cycle[21299] = 1'b1;  wr_cycle[21299] = 1'b0;  addr_rom[21299]='h00000ccc;  wr_data_rom[21299]='h00000000;
    rd_cycle[21300] = 1'b1;  wr_cycle[21300] = 1'b0;  addr_rom[21300]='h00000cd0;  wr_data_rom[21300]='h00000000;
    rd_cycle[21301] = 1'b1;  wr_cycle[21301] = 1'b0;  addr_rom[21301]='h00000cd4;  wr_data_rom[21301]='h00000000;
    rd_cycle[21302] = 1'b1;  wr_cycle[21302] = 1'b0;  addr_rom[21302]='h00000cd8;  wr_data_rom[21302]='h00000000;
    rd_cycle[21303] = 1'b1;  wr_cycle[21303] = 1'b0;  addr_rom[21303]='h00000cdc;  wr_data_rom[21303]='h00000000;
    rd_cycle[21304] = 1'b1;  wr_cycle[21304] = 1'b0;  addr_rom[21304]='h00000ce0;  wr_data_rom[21304]='h00000000;
    rd_cycle[21305] = 1'b1;  wr_cycle[21305] = 1'b0;  addr_rom[21305]='h00000ce4;  wr_data_rom[21305]='h00000000;
    rd_cycle[21306] = 1'b1;  wr_cycle[21306] = 1'b0;  addr_rom[21306]='h00000ce8;  wr_data_rom[21306]='h00000000;
    rd_cycle[21307] = 1'b1;  wr_cycle[21307] = 1'b0;  addr_rom[21307]='h00000cec;  wr_data_rom[21307]='h00000000;
    rd_cycle[21308] = 1'b1;  wr_cycle[21308] = 1'b0;  addr_rom[21308]='h00000cf0;  wr_data_rom[21308]='h00000000;
    rd_cycle[21309] = 1'b1;  wr_cycle[21309] = 1'b0;  addr_rom[21309]='h00000cf4;  wr_data_rom[21309]='h00000000;
    rd_cycle[21310] = 1'b1;  wr_cycle[21310] = 1'b0;  addr_rom[21310]='h00000cf8;  wr_data_rom[21310]='h00000000;
    rd_cycle[21311] = 1'b1;  wr_cycle[21311] = 1'b0;  addr_rom[21311]='h00000cfc;  wr_data_rom[21311]='h00000000;
    rd_cycle[21312] = 1'b1;  wr_cycle[21312] = 1'b0;  addr_rom[21312]='h00000d00;  wr_data_rom[21312]='h00000000;
    rd_cycle[21313] = 1'b1;  wr_cycle[21313] = 1'b0;  addr_rom[21313]='h00000d04;  wr_data_rom[21313]='h00000000;
    rd_cycle[21314] = 1'b1;  wr_cycle[21314] = 1'b0;  addr_rom[21314]='h00000d08;  wr_data_rom[21314]='h00000000;
    rd_cycle[21315] = 1'b1;  wr_cycle[21315] = 1'b0;  addr_rom[21315]='h00000d0c;  wr_data_rom[21315]='h00000000;
    rd_cycle[21316] = 1'b1;  wr_cycle[21316] = 1'b0;  addr_rom[21316]='h00000d10;  wr_data_rom[21316]='h00000000;
    rd_cycle[21317] = 1'b1;  wr_cycle[21317] = 1'b0;  addr_rom[21317]='h00000d14;  wr_data_rom[21317]='h00000000;
    rd_cycle[21318] = 1'b1;  wr_cycle[21318] = 1'b0;  addr_rom[21318]='h00000d18;  wr_data_rom[21318]='h00000000;
    rd_cycle[21319] = 1'b1;  wr_cycle[21319] = 1'b0;  addr_rom[21319]='h00000d1c;  wr_data_rom[21319]='h00000000;
    rd_cycle[21320] = 1'b1;  wr_cycle[21320] = 1'b0;  addr_rom[21320]='h00000d20;  wr_data_rom[21320]='h00000000;
    rd_cycle[21321] = 1'b1;  wr_cycle[21321] = 1'b0;  addr_rom[21321]='h00000d24;  wr_data_rom[21321]='h00000000;
    rd_cycle[21322] = 1'b1;  wr_cycle[21322] = 1'b0;  addr_rom[21322]='h00000d28;  wr_data_rom[21322]='h00000000;
    rd_cycle[21323] = 1'b1;  wr_cycle[21323] = 1'b0;  addr_rom[21323]='h00000d2c;  wr_data_rom[21323]='h00000000;
    rd_cycle[21324] = 1'b1;  wr_cycle[21324] = 1'b0;  addr_rom[21324]='h00000d30;  wr_data_rom[21324]='h00000000;
    rd_cycle[21325] = 1'b1;  wr_cycle[21325] = 1'b0;  addr_rom[21325]='h00000d34;  wr_data_rom[21325]='h00000000;
    rd_cycle[21326] = 1'b1;  wr_cycle[21326] = 1'b0;  addr_rom[21326]='h00000d38;  wr_data_rom[21326]='h00000000;
    rd_cycle[21327] = 1'b1;  wr_cycle[21327] = 1'b0;  addr_rom[21327]='h00000d3c;  wr_data_rom[21327]='h00000000;
    rd_cycle[21328] = 1'b1;  wr_cycle[21328] = 1'b0;  addr_rom[21328]='h00000d40;  wr_data_rom[21328]='h00000000;
    rd_cycle[21329] = 1'b1;  wr_cycle[21329] = 1'b0;  addr_rom[21329]='h00000d44;  wr_data_rom[21329]='h00000000;
    rd_cycle[21330] = 1'b1;  wr_cycle[21330] = 1'b0;  addr_rom[21330]='h00000d48;  wr_data_rom[21330]='h00000000;
    rd_cycle[21331] = 1'b1;  wr_cycle[21331] = 1'b0;  addr_rom[21331]='h00000d4c;  wr_data_rom[21331]='h00000000;
    rd_cycle[21332] = 1'b1;  wr_cycle[21332] = 1'b0;  addr_rom[21332]='h00000d50;  wr_data_rom[21332]='h00000000;
    rd_cycle[21333] = 1'b1;  wr_cycle[21333] = 1'b0;  addr_rom[21333]='h00000d54;  wr_data_rom[21333]='h00000000;
    rd_cycle[21334] = 1'b1;  wr_cycle[21334] = 1'b0;  addr_rom[21334]='h00000d58;  wr_data_rom[21334]='h00000000;
    rd_cycle[21335] = 1'b1;  wr_cycle[21335] = 1'b0;  addr_rom[21335]='h00000d5c;  wr_data_rom[21335]='h00000000;
    rd_cycle[21336] = 1'b1;  wr_cycle[21336] = 1'b0;  addr_rom[21336]='h00000d60;  wr_data_rom[21336]='h00000000;
    rd_cycle[21337] = 1'b1;  wr_cycle[21337] = 1'b0;  addr_rom[21337]='h00000d64;  wr_data_rom[21337]='h00000000;
    rd_cycle[21338] = 1'b1;  wr_cycle[21338] = 1'b0;  addr_rom[21338]='h00000d68;  wr_data_rom[21338]='h00000000;
    rd_cycle[21339] = 1'b1;  wr_cycle[21339] = 1'b0;  addr_rom[21339]='h00000d6c;  wr_data_rom[21339]='h00000000;
    rd_cycle[21340] = 1'b1;  wr_cycle[21340] = 1'b0;  addr_rom[21340]='h00000d70;  wr_data_rom[21340]='h00000000;
    rd_cycle[21341] = 1'b1;  wr_cycle[21341] = 1'b0;  addr_rom[21341]='h00000d74;  wr_data_rom[21341]='h00000000;
    rd_cycle[21342] = 1'b1;  wr_cycle[21342] = 1'b0;  addr_rom[21342]='h00000d78;  wr_data_rom[21342]='h00000000;
    rd_cycle[21343] = 1'b1;  wr_cycle[21343] = 1'b0;  addr_rom[21343]='h00000d7c;  wr_data_rom[21343]='h00000000;
    rd_cycle[21344] = 1'b1;  wr_cycle[21344] = 1'b0;  addr_rom[21344]='h00000d80;  wr_data_rom[21344]='h00000000;
    rd_cycle[21345] = 1'b1;  wr_cycle[21345] = 1'b0;  addr_rom[21345]='h00000d84;  wr_data_rom[21345]='h00000000;
    rd_cycle[21346] = 1'b1;  wr_cycle[21346] = 1'b0;  addr_rom[21346]='h00000d88;  wr_data_rom[21346]='h00000000;
    rd_cycle[21347] = 1'b1;  wr_cycle[21347] = 1'b0;  addr_rom[21347]='h00000d8c;  wr_data_rom[21347]='h00000000;
    rd_cycle[21348] = 1'b1;  wr_cycle[21348] = 1'b0;  addr_rom[21348]='h00000d90;  wr_data_rom[21348]='h00000000;
    rd_cycle[21349] = 1'b1;  wr_cycle[21349] = 1'b0;  addr_rom[21349]='h00000d94;  wr_data_rom[21349]='h00000000;
    rd_cycle[21350] = 1'b1;  wr_cycle[21350] = 1'b0;  addr_rom[21350]='h00000d98;  wr_data_rom[21350]='h00000000;
    rd_cycle[21351] = 1'b1;  wr_cycle[21351] = 1'b0;  addr_rom[21351]='h00000d9c;  wr_data_rom[21351]='h00000000;
    rd_cycle[21352] = 1'b1;  wr_cycle[21352] = 1'b0;  addr_rom[21352]='h00000da0;  wr_data_rom[21352]='h00000000;
    rd_cycle[21353] = 1'b1;  wr_cycle[21353] = 1'b0;  addr_rom[21353]='h00000da4;  wr_data_rom[21353]='h00000000;
    rd_cycle[21354] = 1'b1;  wr_cycle[21354] = 1'b0;  addr_rom[21354]='h00000da8;  wr_data_rom[21354]='h00000000;
    rd_cycle[21355] = 1'b1;  wr_cycle[21355] = 1'b0;  addr_rom[21355]='h00000dac;  wr_data_rom[21355]='h00000000;
    rd_cycle[21356] = 1'b1;  wr_cycle[21356] = 1'b0;  addr_rom[21356]='h00000db0;  wr_data_rom[21356]='h00000000;
    rd_cycle[21357] = 1'b1;  wr_cycle[21357] = 1'b0;  addr_rom[21357]='h00000db4;  wr_data_rom[21357]='h00000000;
    rd_cycle[21358] = 1'b1;  wr_cycle[21358] = 1'b0;  addr_rom[21358]='h00000db8;  wr_data_rom[21358]='h00000000;
    rd_cycle[21359] = 1'b1;  wr_cycle[21359] = 1'b0;  addr_rom[21359]='h00000dbc;  wr_data_rom[21359]='h00000000;
    rd_cycle[21360] = 1'b1;  wr_cycle[21360] = 1'b0;  addr_rom[21360]='h00000dc0;  wr_data_rom[21360]='h00000000;
    rd_cycle[21361] = 1'b1;  wr_cycle[21361] = 1'b0;  addr_rom[21361]='h00000dc4;  wr_data_rom[21361]='h00000000;
    rd_cycle[21362] = 1'b1;  wr_cycle[21362] = 1'b0;  addr_rom[21362]='h00000dc8;  wr_data_rom[21362]='h00000000;
    rd_cycle[21363] = 1'b1;  wr_cycle[21363] = 1'b0;  addr_rom[21363]='h00000dcc;  wr_data_rom[21363]='h00000000;
    rd_cycle[21364] = 1'b1;  wr_cycle[21364] = 1'b0;  addr_rom[21364]='h00000dd0;  wr_data_rom[21364]='h00000000;
    rd_cycle[21365] = 1'b1;  wr_cycle[21365] = 1'b0;  addr_rom[21365]='h00000dd4;  wr_data_rom[21365]='h00000000;
    rd_cycle[21366] = 1'b1;  wr_cycle[21366] = 1'b0;  addr_rom[21366]='h00000dd8;  wr_data_rom[21366]='h00000000;
    rd_cycle[21367] = 1'b1;  wr_cycle[21367] = 1'b0;  addr_rom[21367]='h00000ddc;  wr_data_rom[21367]='h00000000;
    rd_cycle[21368] = 1'b1;  wr_cycle[21368] = 1'b0;  addr_rom[21368]='h00000de0;  wr_data_rom[21368]='h00000000;
    rd_cycle[21369] = 1'b1;  wr_cycle[21369] = 1'b0;  addr_rom[21369]='h00000de4;  wr_data_rom[21369]='h00000000;
    rd_cycle[21370] = 1'b1;  wr_cycle[21370] = 1'b0;  addr_rom[21370]='h00000de8;  wr_data_rom[21370]='h00000000;
    rd_cycle[21371] = 1'b1;  wr_cycle[21371] = 1'b0;  addr_rom[21371]='h00000dec;  wr_data_rom[21371]='h00000000;
    rd_cycle[21372] = 1'b1;  wr_cycle[21372] = 1'b0;  addr_rom[21372]='h00000df0;  wr_data_rom[21372]='h00000000;
    rd_cycle[21373] = 1'b1;  wr_cycle[21373] = 1'b0;  addr_rom[21373]='h00000df4;  wr_data_rom[21373]='h00000000;
    rd_cycle[21374] = 1'b1;  wr_cycle[21374] = 1'b0;  addr_rom[21374]='h00000df8;  wr_data_rom[21374]='h00000000;
    rd_cycle[21375] = 1'b1;  wr_cycle[21375] = 1'b0;  addr_rom[21375]='h00000dfc;  wr_data_rom[21375]='h00000000;
    rd_cycle[21376] = 1'b1;  wr_cycle[21376] = 1'b0;  addr_rom[21376]='h00000e00;  wr_data_rom[21376]='h00000000;
    rd_cycle[21377] = 1'b1;  wr_cycle[21377] = 1'b0;  addr_rom[21377]='h00000e04;  wr_data_rom[21377]='h00000000;
    rd_cycle[21378] = 1'b1;  wr_cycle[21378] = 1'b0;  addr_rom[21378]='h00000e08;  wr_data_rom[21378]='h00000000;
    rd_cycle[21379] = 1'b1;  wr_cycle[21379] = 1'b0;  addr_rom[21379]='h00000e0c;  wr_data_rom[21379]='h00000000;
    rd_cycle[21380] = 1'b1;  wr_cycle[21380] = 1'b0;  addr_rom[21380]='h00000e10;  wr_data_rom[21380]='h00000000;
    rd_cycle[21381] = 1'b1;  wr_cycle[21381] = 1'b0;  addr_rom[21381]='h00000e14;  wr_data_rom[21381]='h00000000;
    rd_cycle[21382] = 1'b1;  wr_cycle[21382] = 1'b0;  addr_rom[21382]='h00000e18;  wr_data_rom[21382]='h00000000;
    rd_cycle[21383] = 1'b1;  wr_cycle[21383] = 1'b0;  addr_rom[21383]='h00000e1c;  wr_data_rom[21383]='h00000000;
    rd_cycle[21384] = 1'b1;  wr_cycle[21384] = 1'b0;  addr_rom[21384]='h00000e20;  wr_data_rom[21384]='h00000000;
    rd_cycle[21385] = 1'b1;  wr_cycle[21385] = 1'b0;  addr_rom[21385]='h00000e24;  wr_data_rom[21385]='h00000000;
    rd_cycle[21386] = 1'b1;  wr_cycle[21386] = 1'b0;  addr_rom[21386]='h00000e28;  wr_data_rom[21386]='h00000000;
    rd_cycle[21387] = 1'b1;  wr_cycle[21387] = 1'b0;  addr_rom[21387]='h00000e2c;  wr_data_rom[21387]='h00000000;
    rd_cycle[21388] = 1'b1;  wr_cycle[21388] = 1'b0;  addr_rom[21388]='h00000e30;  wr_data_rom[21388]='h00000000;
    rd_cycle[21389] = 1'b1;  wr_cycle[21389] = 1'b0;  addr_rom[21389]='h00000e34;  wr_data_rom[21389]='h00000000;
    rd_cycle[21390] = 1'b1;  wr_cycle[21390] = 1'b0;  addr_rom[21390]='h00000e38;  wr_data_rom[21390]='h00000000;
    rd_cycle[21391] = 1'b1;  wr_cycle[21391] = 1'b0;  addr_rom[21391]='h00000e3c;  wr_data_rom[21391]='h00000000;
    rd_cycle[21392] = 1'b1;  wr_cycle[21392] = 1'b0;  addr_rom[21392]='h00000e40;  wr_data_rom[21392]='h00000000;
    rd_cycle[21393] = 1'b1;  wr_cycle[21393] = 1'b0;  addr_rom[21393]='h00000e44;  wr_data_rom[21393]='h00000000;
    rd_cycle[21394] = 1'b1;  wr_cycle[21394] = 1'b0;  addr_rom[21394]='h00000e48;  wr_data_rom[21394]='h00000000;
    rd_cycle[21395] = 1'b1;  wr_cycle[21395] = 1'b0;  addr_rom[21395]='h00000e4c;  wr_data_rom[21395]='h00000000;
    rd_cycle[21396] = 1'b1;  wr_cycle[21396] = 1'b0;  addr_rom[21396]='h00000e50;  wr_data_rom[21396]='h00000000;
    rd_cycle[21397] = 1'b1;  wr_cycle[21397] = 1'b0;  addr_rom[21397]='h00000e54;  wr_data_rom[21397]='h00000000;
    rd_cycle[21398] = 1'b1;  wr_cycle[21398] = 1'b0;  addr_rom[21398]='h00000e58;  wr_data_rom[21398]='h00000000;
    rd_cycle[21399] = 1'b1;  wr_cycle[21399] = 1'b0;  addr_rom[21399]='h00000e5c;  wr_data_rom[21399]='h00000000;
    rd_cycle[21400] = 1'b1;  wr_cycle[21400] = 1'b0;  addr_rom[21400]='h00000e60;  wr_data_rom[21400]='h00000000;
    rd_cycle[21401] = 1'b1;  wr_cycle[21401] = 1'b0;  addr_rom[21401]='h00000e64;  wr_data_rom[21401]='h00000000;
    rd_cycle[21402] = 1'b1;  wr_cycle[21402] = 1'b0;  addr_rom[21402]='h00000e68;  wr_data_rom[21402]='h00000000;
    rd_cycle[21403] = 1'b1;  wr_cycle[21403] = 1'b0;  addr_rom[21403]='h00000e6c;  wr_data_rom[21403]='h00000000;
    rd_cycle[21404] = 1'b1;  wr_cycle[21404] = 1'b0;  addr_rom[21404]='h00000e70;  wr_data_rom[21404]='h00000000;
    rd_cycle[21405] = 1'b1;  wr_cycle[21405] = 1'b0;  addr_rom[21405]='h00000e74;  wr_data_rom[21405]='h00000000;
    rd_cycle[21406] = 1'b1;  wr_cycle[21406] = 1'b0;  addr_rom[21406]='h00000e78;  wr_data_rom[21406]='h00000000;
    rd_cycle[21407] = 1'b1;  wr_cycle[21407] = 1'b0;  addr_rom[21407]='h00000e7c;  wr_data_rom[21407]='h00000000;
    rd_cycle[21408] = 1'b1;  wr_cycle[21408] = 1'b0;  addr_rom[21408]='h00000e80;  wr_data_rom[21408]='h00000000;
    rd_cycle[21409] = 1'b1;  wr_cycle[21409] = 1'b0;  addr_rom[21409]='h00000e84;  wr_data_rom[21409]='h00000000;
    rd_cycle[21410] = 1'b1;  wr_cycle[21410] = 1'b0;  addr_rom[21410]='h00000e88;  wr_data_rom[21410]='h00000000;
    rd_cycle[21411] = 1'b1;  wr_cycle[21411] = 1'b0;  addr_rom[21411]='h00000e8c;  wr_data_rom[21411]='h00000000;
    rd_cycle[21412] = 1'b1;  wr_cycle[21412] = 1'b0;  addr_rom[21412]='h00000e90;  wr_data_rom[21412]='h00000000;
    rd_cycle[21413] = 1'b1;  wr_cycle[21413] = 1'b0;  addr_rom[21413]='h00000e94;  wr_data_rom[21413]='h00000000;
    rd_cycle[21414] = 1'b1;  wr_cycle[21414] = 1'b0;  addr_rom[21414]='h00000e98;  wr_data_rom[21414]='h00000000;
    rd_cycle[21415] = 1'b1;  wr_cycle[21415] = 1'b0;  addr_rom[21415]='h00000e9c;  wr_data_rom[21415]='h00000000;
    rd_cycle[21416] = 1'b1;  wr_cycle[21416] = 1'b0;  addr_rom[21416]='h00000ea0;  wr_data_rom[21416]='h00000000;
    rd_cycle[21417] = 1'b1;  wr_cycle[21417] = 1'b0;  addr_rom[21417]='h00000ea4;  wr_data_rom[21417]='h00000000;
    rd_cycle[21418] = 1'b1;  wr_cycle[21418] = 1'b0;  addr_rom[21418]='h00000ea8;  wr_data_rom[21418]='h00000000;
    rd_cycle[21419] = 1'b1;  wr_cycle[21419] = 1'b0;  addr_rom[21419]='h00000eac;  wr_data_rom[21419]='h00000000;
    rd_cycle[21420] = 1'b1;  wr_cycle[21420] = 1'b0;  addr_rom[21420]='h00000eb0;  wr_data_rom[21420]='h00000000;
    rd_cycle[21421] = 1'b1;  wr_cycle[21421] = 1'b0;  addr_rom[21421]='h00000eb4;  wr_data_rom[21421]='h00000000;
    rd_cycle[21422] = 1'b1;  wr_cycle[21422] = 1'b0;  addr_rom[21422]='h00000eb8;  wr_data_rom[21422]='h00000000;
    rd_cycle[21423] = 1'b1;  wr_cycle[21423] = 1'b0;  addr_rom[21423]='h00000ebc;  wr_data_rom[21423]='h00000000;
    rd_cycle[21424] = 1'b1;  wr_cycle[21424] = 1'b0;  addr_rom[21424]='h00000ec0;  wr_data_rom[21424]='h00000000;
    rd_cycle[21425] = 1'b1;  wr_cycle[21425] = 1'b0;  addr_rom[21425]='h00000ec4;  wr_data_rom[21425]='h00000000;
    rd_cycle[21426] = 1'b1;  wr_cycle[21426] = 1'b0;  addr_rom[21426]='h00000ec8;  wr_data_rom[21426]='h00000000;
    rd_cycle[21427] = 1'b1;  wr_cycle[21427] = 1'b0;  addr_rom[21427]='h00000ecc;  wr_data_rom[21427]='h00000000;
    rd_cycle[21428] = 1'b1;  wr_cycle[21428] = 1'b0;  addr_rom[21428]='h00000ed0;  wr_data_rom[21428]='h00000000;
    rd_cycle[21429] = 1'b1;  wr_cycle[21429] = 1'b0;  addr_rom[21429]='h00000ed4;  wr_data_rom[21429]='h00000000;
    rd_cycle[21430] = 1'b1;  wr_cycle[21430] = 1'b0;  addr_rom[21430]='h00000ed8;  wr_data_rom[21430]='h00000000;
    rd_cycle[21431] = 1'b1;  wr_cycle[21431] = 1'b0;  addr_rom[21431]='h00000edc;  wr_data_rom[21431]='h00000000;
    rd_cycle[21432] = 1'b1;  wr_cycle[21432] = 1'b0;  addr_rom[21432]='h00000ee0;  wr_data_rom[21432]='h00000000;
    rd_cycle[21433] = 1'b1;  wr_cycle[21433] = 1'b0;  addr_rom[21433]='h00000ee4;  wr_data_rom[21433]='h00000000;
    rd_cycle[21434] = 1'b1;  wr_cycle[21434] = 1'b0;  addr_rom[21434]='h00000ee8;  wr_data_rom[21434]='h00000000;
    rd_cycle[21435] = 1'b1;  wr_cycle[21435] = 1'b0;  addr_rom[21435]='h00000eec;  wr_data_rom[21435]='h00000000;
    rd_cycle[21436] = 1'b1;  wr_cycle[21436] = 1'b0;  addr_rom[21436]='h00000ef0;  wr_data_rom[21436]='h00000000;
    rd_cycle[21437] = 1'b1;  wr_cycle[21437] = 1'b0;  addr_rom[21437]='h00000ef4;  wr_data_rom[21437]='h00000000;
    rd_cycle[21438] = 1'b1;  wr_cycle[21438] = 1'b0;  addr_rom[21438]='h00000ef8;  wr_data_rom[21438]='h00000000;
    rd_cycle[21439] = 1'b1;  wr_cycle[21439] = 1'b0;  addr_rom[21439]='h00000efc;  wr_data_rom[21439]='h00000000;
    rd_cycle[21440] = 1'b1;  wr_cycle[21440] = 1'b0;  addr_rom[21440]='h00000f00;  wr_data_rom[21440]='h00000000;
    rd_cycle[21441] = 1'b1;  wr_cycle[21441] = 1'b0;  addr_rom[21441]='h00000f04;  wr_data_rom[21441]='h00000000;
    rd_cycle[21442] = 1'b1;  wr_cycle[21442] = 1'b0;  addr_rom[21442]='h00000f08;  wr_data_rom[21442]='h00000000;
    rd_cycle[21443] = 1'b1;  wr_cycle[21443] = 1'b0;  addr_rom[21443]='h00000f0c;  wr_data_rom[21443]='h00000000;
    rd_cycle[21444] = 1'b1;  wr_cycle[21444] = 1'b0;  addr_rom[21444]='h00000f10;  wr_data_rom[21444]='h00000000;
    rd_cycle[21445] = 1'b1;  wr_cycle[21445] = 1'b0;  addr_rom[21445]='h00000f14;  wr_data_rom[21445]='h00000000;
    rd_cycle[21446] = 1'b1;  wr_cycle[21446] = 1'b0;  addr_rom[21446]='h00000f18;  wr_data_rom[21446]='h00000000;
    rd_cycle[21447] = 1'b1;  wr_cycle[21447] = 1'b0;  addr_rom[21447]='h00000f1c;  wr_data_rom[21447]='h00000000;
    rd_cycle[21448] = 1'b1;  wr_cycle[21448] = 1'b0;  addr_rom[21448]='h00000f20;  wr_data_rom[21448]='h00000000;
    rd_cycle[21449] = 1'b1;  wr_cycle[21449] = 1'b0;  addr_rom[21449]='h00000f24;  wr_data_rom[21449]='h00000000;
    rd_cycle[21450] = 1'b1;  wr_cycle[21450] = 1'b0;  addr_rom[21450]='h00000f28;  wr_data_rom[21450]='h00000000;
    rd_cycle[21451] = 1'b1;  wr_cycle[21451] = 1'b0;  addr_rom[21451]='h00000f2c;  wr_data_rom[21451]='h00000000;
    rd_cycle[21452] = 1'b1;  wr_cycle[21452] = 1'b0;  addr_rom[21452]='h00000f30;  wr_data_rom[21452]='h00000000;
    rd_cycle[21453] = 1'b1;  wr_cycle[21453] = 1'b0;  addr_rom[21453]='h00000f34;  wr_data_rom[21453]='h00000000;
    rd_cycle[21454] = 1'b1;  wr_cycle[21454] = 1'b0;  addr_rom[21454]='h00000f38;  wr_data_rom[21454]='h00000000;
    rd_cycle[21455] = 1'b1;  wr_cycle[21455] = 1'b0;  addr_rom[21455]='h00000f3c;  wr_data_rom[21455]='h00000000;
    rd_cycle[21456] = 1'b1;  wr_cycle[21456] = 1'b0;  addr_rom[21456]='h00000f40;  wr_data_rom[21456]='h00000000;
    rd_cycle[21457] = 1'b1;  wr_cycle[21457] = 1'b0;  addr_rom[21457]='h00000f44;  wr_data_rom[21457]='h00000000;
    rd_cycle[21458] = 1'b1;  wr_cycle[21458] = 1'b0;  addr_rom[21458]='h00000f48;  wr_data_rom[21458]='h00000000;
    rd_cycle[21459] = 1'b1;  wr_cycle[21459] = 1'b0;  addr_rom[21459]='h00000f4c;  wr_data_rom[21459]='h00000000;
    rd_cycle[21460] = 1'b1;  wr_cycle[21460] = 1'b0;  addr_rom[21460]='h00000f50;  wr_data_rom[21460]='h00000000;
    rd_cycle[21461] = 1'b1;  wr_cycle[21461] = 1'b0;  addr_rom[21461]='h00000f54;  wr_data_rom[21461]='h00000000;
    rd_cycle[21462] = 1'b1;  wr_cycle[21462] = 1'b0;  addr_rom[21462]='h00000f58;  wr_data_rom[21462]='h00000000;
    rd_cycle[21463] = 1'b1;  wr_cycle[21463] = 1'b0;  addr_rom[21463]='h00000f5c;  wr_data_rom[21463]='h00000000;
    rd_cycle[21464] = 1'b1;  wr_cycle[21464] = 1'b0;  addr_rom[21464]='h00000f60;  wr_data_rom[21464]='h00000000;
    rd_cycle[21465] = 1'b1;  wr_cycle[21465] = 1'b0;  addr_rom[21465]='h00000f64;  wr_data_rom[21465]='h00000000;
    rd_cycle[21466] = 1'b1;  wr_cycle[21466] = 1'b0;  addr_rom[21466]='h00000f68;  wr_data_rom[21466]='h00000000;
    rd_cycle[21467] = 1'b1;  wr_cycle[21467] = 1'b0;  addr_rom[21467]='h00000f6c;  wr_data_rom[21467]='h00000000;
    rd_cycle[21468] = 1'b1;  wr_cycle[21468] = 1'b0;  addr_rom[21468]='h00000f70;  wr_data_rom[21468]='h00000000;
    rd_cycle[21469] = 1'b1;  wr_cycle[21469] = 1'b0;  addr_rom[21469]='h00000f74;  wr_data_rom[21469]='h00000000;
    rd_cycle[21470] = 1'b1;  wr_cycle[21470] = 1'b0;  addr_rom[21470]='h00000f78;  wr_data_rom[21470]='h00000000;
    rd_cycle[21471] = 1'b1;  wr_cycle[21471] = 1'b0;  addr_rom[21471]='h00000f7c;  wr_data_rom[21471]='h00000000;
    rd_cycle[21472] = 1'b1;  wr_cycle[21472] = 1'b0;  addr_rom[21472]='h00000f80;  wr_data_rom[21472]='h00000000;
    rd_cycle[21473] = 1'b1;  wr_cycle[21473] = 1'b0;  addr_rom[21473]='h00000f84;  wr_data_rom[21473]='h00000000;
    rd_cycle[21474] = 1'b1;  wr_cycle[21474] = 1'b0;  addr_rom[21474]='h00000f88;  wr_data_rom[21474]='h00000000;
    rd_cycle[21475] = 1'b1;  wr_cycle[21475] = 1'b0;  addr_rom[21475]='h00000f8c;  wr_data_rom[21475]='h00000000;
    rd_cycle[21476] = 1'b1;  wr_cycle[21476] = 1'b0;  addr_rom[21476]='h00000f90;  wr_data_rom[21476]='h00000000;
    rd_cycle[21477] = 1'b1;  wr_cycle[21477] = 1'b0;  addr_rom[21477]='h00000f94;  wr_data_rom[21477]='h00000000;
    rd_cycle[21478] = 1'b1;  wr_cycle[21478] = 1'b0;  addr_rom[21478]='h00000f98;  wr_data_rom[21478]='h00000000;
    rd_cycle[21479] = 1'b1;  wr_cycle[21479] = 1'b0;  addr_rom[21479]='h00000f9c;  wr_data_rom[21479]='h00000000;
    rd_cycle[21480] = 1'b1;  wr_cycle[21480] = 1'b0;  addr_rom[21480]='h00000fa0;  wr_data_rom[21480]='h00000000;
    rd_cycle[21481] = 1'b1;  wr_cycle[21481] = 1'b0;  addr_rom[21481]='h00000fa4;  wr_data_rom[21481]='h00000000;
    rd_cycle[21482] = 1'b1;  wr_cycle[21482] = 1'b0;  addr_rom[21482]='h00000fa8;  wr_data_rom[21482]='h00000000;
    rd_cycle[21483] = 1'b1;  wr_cycle[21483] = 1'b0;  addr_rom[21483]='h00000fac;  wr_data_rom[21483]='h00000000;
    rd_cycle[21484] = 1'b1;  wr_cycle[21484] = 1'b0;  addr_rom[21484]='h00000fb0;  wr_data_rom[21484]='h00000000;
    rd_cycle[21485] = 1'b1;  wr_cycle[21485] = 1'b0;  addr_rom[21485]='h00000fb4;  wr_data_rom[21485]='h00000000;
    rd_cycle[21486] = 1'b1;  wr_cycle[21486] = 1'b0;  addr_rom[21486]='h00000fb8;  wr_data_rom[21486]='h00000000;
    rd_cycle[21487] = 1'b1;  wr_cycle[21487] = 1'b0;  addr_rom[21487]='h00000fbc;  wr_data_rom[21487]='h00000000;
    rd_cycle[21488] = 1'b1;  wr_cycle[21488] = 1'b0;  addr_rom[21488]='h00000fc0;  wr_data_rom[21488]='h00000000;
    rd_cycle[21489] = 1'b1;  wr_cycle[21489] = 1'b0;  addr_rom[21489]='h00000fc4;  wr_data_rom[21489]='h00000000;
    rd_cycle[21490] = 1'b1;  wr_cycle[21490] = 1'b0;  addr_rom[21490]='h00000fc8;  wr_data_rom[21490]='h00000000;
    rd_cycle[21491] = 1'b1;  wr_cycle[21491] = 1'b0;  addr_rom[21491]='h00000fcc;  wr_data_rom[21491]='h00000000;
    rd_cycle[21492] = 1'b1;  wr_cycle[21492] = 1'b0;  addr_rom[21492]='h00000fd0;  wr_data_rom[21492]='h00000000;
    rd_cycle[21493] = 1'b1;  wr_cycle[21493] = 1'b0;  addr_rom[21493]='h00000fd4;  wr_data_rom[21493]='h00000000;
    rd_cycle[21494] = 1'b1;  wr_cycle[21494] = 1'b0;  addr_rom[21494]='h00000fd8;  wr_data_rom[21494]='h00000000;
    rd_cycle[21495] = 1'b1;  wr_cycle[21495] = 1'b0;  addr_rom[21495]='h00000fdc;  wr_data_rom[21495]='h00000000;
    rd_cycle[21496] = 1'b1;  wr_cycle[21496] = 1'b0;  addr_rom[21496]='h00000fe0;  wr_data_rom[21496]='h00000000;
    rd_cycle[21497] = 1'b1;  wr_cycle[21497] = 1'b0;  addr_rom[21497]='h00000fe4;  wr_data_rom[21497]='h00000000;
    rd_cycle[21498] = 1'b1;  wr_cycle[21498] = 1'b0;  addr_rom[21498]='h00000fe8;  wr_data_rom[21498]='h00000000;
    rd_cycle[21499] = 1'b1;  wr_cycle[21499] = 1'b0;  addr_rom[21499]='h00000fec;  wr_data_rom[21499]='h00000000;
    rd_cycle[21500] = 1'b1;  wr_cycle[21500] = 1'b0;  addr_rom[21500]='h00000ff0;  wr_data_rom[21500]='h00000000;
    rd_cycle[21501] = 1'b1;  wr_cycle[21501] = 1'b0;  addr_rom[21501]='h00000ff4;  wr_data_rom[21501]='h00000000;
    rd_cycle[21502] = 1'b1;  wr_cycle[21502] = 1'b0;  addr_rom[21502]='h00000ff8;  wr_data_rom[21502]='h00000000;
    rd_cycle[21503] = 1'b1;  wr_cycle[21503] = 1'b0;  addr_rom[21503]='h00000ffc;  wr_data_rom[21503]='h00000000;
    rd_cycle[21504] = 1'b1;  wr_cycle[21504] = 1'b0;  addr_rom[21504]='h00001000;  wr_data_rom[21504]='h00000000;
    rd_cycle[21505] = 1'b1;  wr_cycle[21505] = 1'b0;  addr_rom[21505]='h00001004;  wr_data_rom[21505]='h00000000;
    rd_cycle[21506] = 1'b1;  wr_cycle[21506] = 1'b0;  addr_rom[21506]='h00001008;  wr_data_rom[21506]='h00000000;
    rd_cycle[21507] = 1'b1;  wr_cycle[21507] = 1'b0;  addr_rom[21507]='h0000100c;  wr_data_rom[21507]='h00000000;
    rd_cycle[21508] = 1'b1;  wr_cycle[21508] = 1'b0;  addr_rom[21508]='h00001010;  wr_data_rom[21508]='h00000000;
    rd_cycle[21509] = 1'b1;  wr_cycle[21509] = 1'b0;  addr_rom[21509]='h00001014;  wr_data_rom[21509]='h00000000;
    rd_cycle[21510] = 1'b1;  wr_cycle[21510] = 1'b0;  addr_rom[21510]='h00001018;  wr_data_rom[21510]='h00000000;
    rd_cycle[21511] = 1'b1;  wr_cycle[21511] = 1'b0;  addr_rom[21511]='h0000101c;  wr_data_rom[21511]='h00000000;
    rd_cycle[21512] = 1'b1;  wr_cycle[21512] = 1'b0;  addr_rom[21512]='h00001020;  wr_data_rom[21512]='h00000000;
    rd_cycle[21513] = 1'b1;  wr_cycle[21513] = 1'b0;  addr_rom[21513]='h00001024;  wr_data_rom[21513]='h00000000;
    rd_cycle[21514] = 1'b1;  wr_cycle[21514] = 1'b0;  addr_rom[21514]='h00001028;  wr_data_rom[21514]='h00000000;
    rd_cycle[21515] = 1'b1;  wr_cycle[21515] = 1'b0;  addr_rom[21515]='h0000102c;  wr_data_rom[21515]='h00000000;
    rd_cycle[21516] = 1'b1;  wr_cycle[21516] = 1'b0;  addr_rom[21516]='h00001030;  wr_data_rom[21516]='h00000000;
    rd_cycle[21517] = 1'b1;  wr_cycle[21517] = 1'b0;  addr_rom[21517]='h00001034;  wr_data_rom[21517]='h00000000;
    rd_cycle[21518] = 1'b1;  wr_cycle[21518] = 1'b0;  addr_rom[21518]='h00001038;  wr_data_rom[21518]='h00000000;
    rd_cycle[21519] = 1'b1;  wr_cycle[21519] = 1'b0;  addr_rom[21519]='h0000103c;  wr_data_rom[21519]='h00000000;
    rd_cycle[21520] = 1'b1;  wr_cycle[21520] = 1'b0;  addr_rom[21520]='h00001040;  wr_data_rom[21520]='h00000000;
    rd_cycle[21521] = 1'b1;  wr_cycle[21521] = 1'b0;  addr_rom[21521]='h00001044;  wr_data_rom[21521]='h00000000;
    rd_cycle[21522] = 1'b1;  wr_cycle[21522] = 1'b0;  addr_rom[21522]='h00001048;  wr_data_rom[21522]='h00000000;
    rd_cycle[21523] = 1'b1;  wr_cycle[21523] = 1'b0;  addr_rom[21523]='h0000104c;  wr_data_rom[21523]='h00000000;
    rd_cycle[21524] = 1'b1;  wr_cycle[21524] = 1'b0;  addr_rom[21524]='h00001050;  wr_data_rom[21524]='h00000000;
    rd_cycle[21525] = 1'b1;  wr_cycle[21525] = 1'b0;  addr_rom[21525]='h00001054;  wr_data_rom[21525]='h00000000;
    rd_cycle[21526] = 1'b1;  wr_cycle[21526] = 1'b0;  addr_rom[21526]='h00001058;  wr_data_rom[21526]='h00000000;
    rd_cycle[21527] = 1'b1;  wr_cycle[21527] = 1'b0;  addr_rom[21527]='h0000105c;  wr_data_rom[21527]='h00000000;
    rd_cycle[21528] = 1'b1;  wr_cycle[21528] = 1'b0;  addr_rom[21528]='h00001060;  wr_data_rom[21528]='h00000000;
    rd_cycle[21529] = 1'b1;  wr_cycle[21529] = 1'b0;  addr_rom[21529]='h00001064;  wr_data_rom[21529]='h00000000;
    rd_cycle[21530] = 1'b1;  wr_cycle[21530] = 1'b0;  addr_rom[21530]='h00001068;  wr_data_rom[21530]='h00000000;
    rd_cycle[21531] = 1'b1;  wr_cycle[21531] = 1'b0;  addr_rom[21531]='h0000106c;  wr_data_rom[21531]='h00000000;
    rd_cycle[21532] = 1'b1;  wr_cycle[21532] = 1'b0;  addr_rom[21532]='h00001070;  wr_data_rom[21532]='h00000000;
    rd_cycle[21533] = 1'b1;  wr_cycle[21533] = 1'b0;  addr_rom[21533]='h00001074;  wr_data_rom[21533]='h00000000;
    rd_cycle[21534] = 1'b1;  wr_cycle[21534] = 1'b0;  addr_rom[21534]='h00001078;  wr_data_rom[21534]='h00000000;
    rd_cycle[21535] = 1'b1;  wr_cycle[21535] = 1'b0;  addr_rom[21535]='h0000107c;  wr_data_rom[21535]='h00000000;
    rd_cycle[21536] = 1'b1;  wr_cycle[21536] = 1'b0;  addr_rom[21536]='h00001080;  wr_data_rom[21536]='h00000000;
    rd_cycle[21537] = 1'b1;  wr_cycle[21537] = 1'b0;  addr_rom[21537]='h00001084;  wr_data_rom[21537]='h00000000;
    rd_cycle[21538] = 1'b1;  wr_cycle[21538] = 1'b0;  addr_rom[21538]='h00001088;  wr_data_rom[21538]='h00000000;
    rd_cycle[21539] = 1'b1;  wr_cycle[21539] = 1'b0;  addr_rom[21539]='h0000108c;  wr_data_rom[21539]='h00000000;
    rd_cycle[21540] = 1'b1;  wr_cycle[21540] = 1'b0;  addr_rom[21540]='h00001090;  wr_data_rom[21540]='h00000000;
    rd_cycle[21541] = 1'b1;  wr_cycle[21541] = 1'b0;  addr_rom[21541]='h00001094;  wr_data_rom[21541]='h00000000;
    rd_cycle[21542] = 1'b1;  wr_cycle[21542] = 1'b0;  addr_rom[21542]='h00001098;  wr_data_rom[21542]='h00000000;
    rd_cycle[21543] = 1'b1;  wr_cycle[21543] = 1'b0;  addr_rom[21543]='h0000109c;  wr_data_rom[21543]='h00000000;
    rd_cycle[21544] = 1'b1;  wr_cycle[21544] = 1'b0;  addr_rom[21544]='h000010a0;  wr_data_rom[21544]='h00000000;
    rd_cycle[21545] = 1'b1;  wr_cycle[21545] = 1'b0;  addr_rom[21545]='h000010a4;  wr_data_rom[21545]='h00000000;
    rd_cycle[21546] = 1'b1;  wr_cycle[21546] = 1'b0;  addr_rom[21546]='h000010a8;  wr_data_rom[21546]='h00000000;
    rd_cycle[21547] = 1'b1;  wr_cycle[21547] = 1'b0;  addr_rom[21547]='h000010ac;  wr_data_rom[21547]='h00000000;
    rd_cycle[21548] = 1'b1;  wr_cycle[21548] = 1'b0;  addr_rom[21548]='h000010b0;  wr_data_rom[21548]='h00000000;
    rd_cycle[21549] = 1'b1;  wr_cycle[21549] = 1'b0;  addr_rom[21549]='h000010b4;  wr_data_rom[21549]='h00000000;
    rd_cycle[21550] = 1'b1;  wr_cycle[21550] = 1'b0;  addr_rom[21550]='h000010b8;  wr_data_rom[21550]='h00000000;
    rd_cycle[21551] = 1'b1;  wr_cycle[21551] = 1'b0;  addr_rom[21551]='h000010bc;  wr_data_rom[21551]='h00000000;
    rd_cycle[21552] = 1'b1;  wr_cycle[21552] = 1'b0;  addr_rom[21552]='h000010c0;  wr_data_rom[21552]='h00000000;
    rd_cycle[21553] = 1'b1;  wr_cycle[21553] = 1'b0;  addr_rom[21553]='h000010c4;  wr_data_rom[21553]='h00000000;
    rd_cycle[21554] = 1'b1;  wr_cycle[21554] = 1'b0;  addr_rom[21554]='h000010c8;  wr_data_rom[21554]='h00000000;
    rd_cycle[21555] = 1'b1;  wr_cycle[21555] = 1'b0;  addr_rom[21555]='h000010cc;  wr_data_rom[21555]='h00000000;
    rd_cycle[21556] = 1'b1;  wr_cycle[21556] = 1'b0;  addr_rom[21556]='h000010d0;  wr_data_rom[21556]='h00000000;
    rd_cycle[21557] = 1'b1;  wr_cycle[21557] = 1'b0;  addr_rom[21557]='h000010d4;  wr_data_rom[21557]='h00000000;
    rd_cycle[21558] = 1'b1;  wr_cycle[21558] = 1'b0;  addr_rom[21558]='h000010d8;  wr_data_rom[21558]='h00000000;
    rd_cycle[21559] = 1'b1;  wr_cycle[21559] = 1'b0;  addr_rom[21559]='h000010dc;  wr_data_rom[21559]='h00000000;
    rd_cycle[21560] = 1'b1;  wr_cycle[21560] = 1'b0;  addr_rom[21560]='h000010e0;  wr_data_rom[21560]='h00000000;
    rd_cycle[21561] = 1'b1;  wr_cycle[21561] = 1'b0;  addr_rom[21561]='h000010e4;  wr_data_rom[21561]='h00000000;
    rd_cycle[21562] = 1'b1;  wr_cycle[21562] = 1'b0;  addr_rom[21562]='h000010e8;  wr_data_rom[21562]='h00000000;
    rd_cycle[21563] = 1'b1;  wr_cycle[21563] = 1'b0;  addr_rom[21563]='h000010ec;  wr_data_rom[21563]='h00000000;
    rd_cycle[21564] = 1'b1;  wr_cycle[21564] = 1'b0;  addr_rom[21564]='h000010f0;  wr_data_rom[21564]='h00000000;
    rd_cycle[21565] = 1'b1;  wr_cycle[21565] = 1'b0;  addr_rom[21565]='h000010f4;  wr_data_rom[21565]='h00000000;
    rd_cycle[21566] = 1'b1;  wr_cycle[21566] = 1'b0;  addr_rom[21566]='h000010f8;  wr_data_rom[21566]='h00000000;
    rd_cycle[21567] = 1'b1;  wr_cycle[21567] = 1'b0;  addr_rom[21567]='h000010fc;  wr_data_rom[21567]='h00000000;
    rd_cycle[21568] = 1'b1;  wr_cycle[21568] = 1'b0;  addr_rom[21568]='h00001100;  wr_data_rom[21568]='h00000000;
    rd_cycle[21569] = 1'b1;  wr_cycle[21569] = 1'b0;  addr_rom[21569]='h00001104;  wr_data_rom[21569]='h00000000;
    rd_cycle[21570] = 1'b1;  wr_cycle[21570] = 1'b0;  addr_rom[21570]='h00001108;  wr_data_rom[21570]='h00000000;
    rd_cycle[21571] = 1'b1;  wr_cycle[21571] = 1'b0;  addr_rom[21571]='h0000110c;  wr_data_rom[21571]='h00000000;
    rd_cycle[21572] = 1'b1;  wr_cycle[21572] = 1'b0;  addr_rom[21572]='h00001110;  wr_data_rom[21572]='h00000000;
    rd_cycle[21573] = 1'b1;  wr_cycle[21573] = 1'b0;  addr_rom[21573]='h00001114;  wr_data_rom[21573]='h00000000;
    rd_cycle[21574] = 1'b1;  wr_cycle[21574] = 1'b0;  addr_rom[21574]='h00001118;  wr_data_rom[21574]='h00000000;
    rd_cycle[21575] = 1'b1;  wr_cycle[21575] = 1'b0;  addr_rom[21575]='h0000111c;  wr_data_rom[21575]='h00000000;
    rd_cycle[21576] = 1'b1;  wr_cycle[21576] = 1'b0;  addr_rom[21576]='h00001120;  wr_data_rom[21576]='h00000000;
    rd_cycle[21577] = 1'b1;  wr_cycle[21577] = 1'b0;  addr_rom[21577]='h00001124;  wr_data_rom[21577]='h00000000;
    rd_cycle[21578] = 1'b1;  wr_cycle[21578] = 1'b0;  addr_rom[21578]='h00001128;  wr_data_rom[21578]='h00000000;
    rd_cycle[21579] = 1'b1;  wr_cycle[21579] = 1'b0;  addr_rom[21579]='h0000112c;  wr_data_rom[21579]='h00000000;
    rd_cycle[21580] = 1'b1;  wr_cycle[21580] = 1'b0;  addr_rom[21580]='h00001130;  wr_data_rom[21580]='h00000000;
    rd_cycle[21581] = 1'b1;  wr_cycle[21581] = 1'b0;  addr_rom[21581]='h00001134;  wr_data_rom[21581]='h00000000;
    rd_cycle[21582] = 1'b1;  wr_cycle[21582] = 1'b0;  addr_rom[21582]='h00001138;  wr_data_rom[21582]='h00000000;
    rd_cycle[21583] = 1'b1;  wr_cycle[21583] = 1'b0;  addr_rom[21583]='h0000113c;  wr_data_rom[21583]='h00000000;
    rd_cycle[21584] = 1'b1;  wr_cycle[21584] = 1'b0;  addr_rom[21584]='h00001140;  wr_data_rom[21584]='h00000000;
    rd_cycle[21585] = 1'b1;  wr_cycle[21585] = 1'b0;  addr_rom[21585]='h00001144;  wr_data_rom[21585]='h00000000;
    rd_cycle[21586] = 1'b1;  wr_cycle[21586] = 1'b0;  addr_rom[21586]='h00001148;  wr_data_rom[21586]='h00000000;
    rd_cycle[21587] = 1'b1;  wr_cycle[21587] = 1'b0;  addr_rom[21587]='h0000114c;  wr_data_rom[21587]='h00000000;
    rd_cycle[21588] = 1'b1;  wr_cycle[21588] = 1'b0;  addr_rom[21588]='h00001150;  wr_data_rom[21588]='h00000000;
    rd_cycle[21589] = 1'b1;  wr_cycle[21589] = 1'b0;  addr_rom[21589]='h00001154;  wr_data_rom[21589]='h00000000;
    rd_cycle[21590] = 1'b1;  wr_cycle[21590] = 1'b0;  addr_rom[21590]='h00001158;  wr_data_rom[21590]='h00000000;
    rd_cycle[21591] = 1'b1;  wr_cycle[21591] = 1'b0;  addr_rom[21591]='h0000115c;  wr_data_rom[21591]='h00000000;
    rd_cycle[21592] = 1'b1;  wr_cycle[21592] = 1'b0;  addr_rom[21592]='h00001160;  wr_data_rom[21592]='h00000000;
    rd_cycle[21593] = 1'b1;  wr_cycle[21593] = 1'b0;  addr_rom[21593]='h00001164;  wr_data_rom[21593]='h00000000;
    rd_cycle[21594] = 1'b1;  wr_cycle[21594] = 1'b0;  addr_rom[21594]='h00001168;  wr_data_rom[21594]='h00000000;
    rd_cycle[21595] = 1'b1;  wr_cycle[21595] = 1'b0;  addr_rom[21595]='h0000116c;  wr_data_rom[21595]='h00000000;
    rd_cycle[21596] = 1'b1;  wr_cycle[21596] = 1'b0;  addr_rom[21596]='h00001170;  wr_data_rom[21596]='h00000000;
    rd_cycle[21597] = 1'b1;  wr_cycle[21597] = 1'b0;  addr_rom[21597]='h00001174;  wr_data_rom[21597]='h00000000;
    rd_cycle[21598] = 1'b1;  wr_cycle[21598] = 1'b0;  addr_rom[21598]='h00001178;  wr_data_rom[21598]='h00000000;
    rd_cycle[21599] = 1'b1;  wr_cycle[21599] = 1'b0;  addr_rom[21599]='h0000117c;  wr_data_rom[21599]='h00000000;
    rd_cycle[21600] = 1'b1;  wr_cycle[21600] = 1'b0;  addr_rom[21600]='h00001180;  wr_data_rom[21600]='h00000000;
    rd_cycle[21601] = 1'b1;  wr_cycle[21601] = 1'b0;  addr_rom[21601]='h00001184;  wr_data_rom[21601]='h00000000;
    rd_cycle[21602] = 1'b1;  wr_cycle[21602] = 1'b0;  addr_rom[21602]='h00001188;  wr_data_rom[21602]='h00000000;
    rd_cycle[21603] = 1'b1;  wr_cycle[21603] = 1'b0;  addr_rom[21603]='h0000118c;  wr_data_rom[21603]='h00000000;
    rd_cycle[21604] = 1'b1;  wr_cycle[21604] = 1'b0;  addr_rom[21604]='h00001190;  wr_data_rom[21604]='h00000000;
    rd_cycle[21605] = 1'b1;  wr_cycle[21605] = 1'b0;  addr_rom[21605]='h00001194;  wr_data_rom[21605]='h00000000;
    rd_cycle[21606] = 1'b1;  wr_cycle[21606] = 1'b0;  addr_rom[21606]='h00001198;  wr_data_rom[21606]='h00000000;
    rd_cycle[21607] = 1'b1;  wr_cycle[21607] = 1'b0;  addr_rom[21607]='h0000119c;  wr_data_rom[21607]='h00000000;
    rd_cycle[21608] = 1'b1;  wr_cycle[21608] = 1'b0;  addr_rom[21608]='h000011a0;  wr_data_rom[21608]='h00000000;
    rd_cycle[21609] = 1'b1;  wr_cycle[21609] = 1'b0;  addr_rom[21609]='h000011a4;  wr_data_rom[21609]='h00000000;
    rd_cycle[21610] = 1'b1;  wr_cycle[21610] = 1'b0;  addr_rom[21610]='h000011a8;  wr_data_rom[21610]='h00000000;
    rd_cycle[21611] = 1'b1;  wr_cycle[21611] = 1'b0;  addr_rom[21611]='h000011ac;  wr_data_rom[21611]='h00000000;
    rd_cycle[21612] = 1'b1;  wr_cycle[21612] = 1'b0;  addr_rom[21612]='h000011b0;  wr_data_rom[21612]='h00000000;
    rd_cycle[21613] = 1'b1;  wr_cycle[21613] = 1'b0;  addr_rom[21613]='h000011b4;  wr_data_rom[21613]='h00000000;
    rd_cycle[21614] = 1'b1;  wr_cycle[21614] = 1'b0;  addr_rom[21614]='h000011b8;  wr_data_rom[21614]='h00000000;
    rd_cycle[21615] = 1'b1;  wr_cycle[21615] = 1'b0;  addr_rom[21615]='h000011bc;  wr_data_rom[21615]='h00000000;
    rd_cycle[21616] = 1'b1;  wr_cycle[21616] = 1'b0;  addr_rom[21616]='h000011c0;  wr_data_rom[21616]='h00000000;
    rd_cycle[21617] = 1'b1;  wr_cycle[21617] = 1'b0;  addr_rom[21617]='h000011c4;  wr_data_rom[21617]='h00000000;
    rd_cycle[21618] = 1'b1;  wr_cycle[21618] = 1'b0;  addr_rom[21618]='h000011c8;  wr_data_rom[21618]='h00000000;
    rd_cycle[21619] = 1'b1;  wr_cycle[21619] = 1'b0;  addr_rom[21619]='h000011cc;  wr_data_rom[21619]='h00000000;
    rd_cycle[21620] = 1'b1;  wr_cycle[21620] = 1'b0;  addr_rom[21620]='h000011d0;  wr_data_rom[21620]='h00000000;
    rd_cycle[21621] = 1'b1;  wr_cycle[21621] = 1'b0;  addr_rom[21621]='h000011d4;  wr_data_rom[21621]='h00000000;
    rd_cycle[21622] = 1'b1;  wr_cycle[21622] = 1'b0;  addr_rom[21622]='h000011d8;  wr_data_rom[21622]='h00000000;
    rd_cycle[21623] = 1'b1;  wr_cycle[21623] = 1'b0;  addr_rom[21623]='h000011dc;  wr_data_rom[21623]='h00000000;
    rd_cycle[21624] = 1'b1;  wr_cycle[21624] = 1'b0;  addr_rom[21624]='h000011e0;  wr_data_rom[21624]='h00000000;
    rd_cycle[21625] = 1'b1;  wr_cycle[21625] = 1'b0;  addr_rom[21625]='h000011e4;  wr_data_rom[21625]='h00000000;
    rd_cycle[21626] = 1'b1;  wr_cycle[21626] = 1'b0;  addr_rom[21626]='h000011e8;  wr_data_rom[21626]='h00000000;
    rd_cycle[21627] = 1'b1;  wr_cycle[21627] = 1'b0;  addr_rom[21627]='h000011ec;  wr_data_rom[21627]='h00000000;
    rd_cycle[21628] = 1'b1;  wr_cycle[21628] = 1'b0;  addr_rom[21628]='h000011f0;  wr_data_rom[21628]='h00000000;
    rd_cycle[21629] = 1'b1;  wr_cycle[21629] = 1'b0;  addr_rom[21629]='h000011f4;  wr_data_rom[21629]='h00000000;
    rd_cycle[21630] = 1'b1;  wr_cycle[21630] = 1'b0;  addr_rom[21630]='h000011f8;  wr_data_rom[21630]='h00000000;
    rd_cycle[21631] = 1'b1;  wr_cycle[21631] = 1'b0;  addr_rom[21631]='h000011fc;  wr_data_rom[21631]='h00000000;
    rd_cycle[21632] = 1'b1;  wr_cycle[21632] = 1'b0;  addr_rom[21632]='h00001200;  wr_data_rom[21632]='h00000000;
    rd_cycle[21633] = 1'b1;  wr_cycle[21633] = 1'b0;  addr_rom[21633]='h00001204;  wr_data_rom[21633]='h00000000;
    rd_cycle[21634] = 1'b1;  wr_cycle[21634] = 1'b0;  addr_rom[21634]='h00001208;  wr_data_rom[21634]='h00000000;
    rd_cycle[21635] = 1'b1;  wr_cycle[21635] = 1'b0;  addr_rom[21635]='h0000120c;  wr_data_rom[21635]='h00000000;
    rd_cycle[21636] = 1'b1;  wr_cycle[21636] = 1'b0;  addr_rom[21636]='h00001210;  wr_data_rom[21636]='h00000000;
    rd_cycle[21637] = 1'b1;  wr_cycle[21637] = 1'b0;  addr_rom[21637]='h00001214;  wr_data_rom[21637]='h00000000;
    rd_cycle[21638] = 1'b1;  wr_cycle[21638] = 1'b0;  addr_rom[21638]='h00001218;  wr_data_rom[21638]='h00000000;
    rd_cycle[21639] = 1'b1;  wr_cycle[21639] = 1'b0;  addr_rom[21639]='h0000121c;  wr_data_rom[21639]='h00000000;
    rd_cycle[21640] = 1'b1;  wr_cycle[21640] = 1'b0;  addr_rom[21640]='h00001220;  wr_data_rom[21640]='h00000000;
    rd_cycle[21641] = 1'b1;  wr_cycle[21641] = 1'b0;  addr_rom[21641]='h00001224;  wr_data_rom[21641]='h00000000;
    rd_cycle[21642] = 1'b1;  wr_cycle[21642] = 1'b0;  addr_rom[21642]='h00001228;  wr_data_rom[21642]='h00000000;
    rd_cycle[21643] = 1'b1;  wr_cycle[21643] = 1'b0;  addr_rom[21643]='h0000122c;  wr_data_rom[21643]='h00000000;
    rd_cycle[21644] = 1'b1;  wr_cycle[21644] = 1'b0;  addr_rom[21644]='h00001230;  wr_data_rom[21644]='h00000000;
    rd_cycle[21645] = 1'b1;  wr_cycle[21645] = 1'b0;  addr_rom[21645]='h00001234;  wr_data_rom[21645]='h00000000;
    rd_cycle[21646] = 1'b1;  wr_cycle[21646] = 1'b0;  addr_rom[21646]='h00001238;  wr_data_rom[21646]='h00000000;
    rd_cycle[21647] = 1'b1;  wr_cycle[21647] = 1'b0;  addr_rom[21647]='h0000123c;  wr_data_rom[21647]='h00000000;
    rd_cycle[21648] = 1'b1;  wr_cycle[21648] = 1'b0;  addr_rom[21648]='h00001240;  wr_data_rom[21648]='h00000000;
    rd_cycle[21649] = 1'b1;  wr_cycle[21649] = 1'b0;  addr_rom[21649]='h00001244;  wr_data_rom[21649]='h00000000;
    rd_cycle[21650] = 1'b1;  wr_cycle[21650] = 1'b0;  addr_rom[21650]='h00001248;  wr_data_rom[21650]='h00000000;
    rd_cycle[21651] = 1'b1;  wr_cycle[21651] = 1'b0;  addr_rom[21651]='h0000124c;  wr_data_rom[21651]='h00000000;
    rd_cycle[21652] = 1'b1;  wr_cycle[21652] = 1'b0;  addr_rom[21652]='h00001250;  wr_data_rom[21652]='h00000000;
    rd_cycle[21653] = 1'b1;  wr_cycle[21653] = 1'b0;  addr_rom[21653]='h00001254;  wr_data_rom[21653]='h00000000;
    rd_cycle[21654] = 1'b1;  wr_cycle[21654] = 1'b0;  addr_rom[21654]='h00001258;  wr_data_rom[21654]='h00000000;
    rd_cycle[21655] = 1'b1;  wr_cycle[21655] = 1'b0;  addr_rom[21655]='h0000125c;  wr_data_rom[21655]='h00000000;
    rd_cycle[21656] = 1'b1;  wr_cycle[21656] = 1'b0;  addr_rom[21656]='h00001260;  wr_data_rom[21656]='h00000000;
    rd_cycle[21657] = 1'b1;  wr_cycle[21657] = 1'b0;  addr_rom[21657]='h00001264;  wr_data_rom[21657]='h00000000;
    rd_cycle[21658] = 1'b1;  wr_cycle[21658] = 1'b0;  addr_rom[21658]='h00001268;  wr_data_rom[21658]='h00000000;
    rd_cycle[21659] = 1'b1;  wr_cycle[21659] = 1'b0;  addr_rom[21659]='h0000126c;  wr_data_rom[21659]='h00000000;
    rd_cycle[21660] = 1'b1;  wr_cycle[21660] = 1'b0;  addr_rom[21660]='h00001270;  wr_data_rom[21660]='h00000000;
    rd_cycle[21661] = 1'b1;  wr_cycle[21661] = 1'b0;  addr_rom[21661]='h00001274;  wr_data_rom[21661]='h00000000;
    rd_cycle[21662] = 1'b1;  wr_cycle[21662] = 1'b0;  addr_rom[21662]='h00001278;  wr_data_rom[21662]='h00000000;
    rd_cycle[21663] = 1'b1;  wr_cycle[21663] = 1'b0;  addr_rom[21663]='h0000127c;  wr_data_rom[21663]='h00000000;
    rd_cycle[21664] = 1'b1;  wr_cycle[21664] = 1'b0;  addr_rom[21664]='h00001280;  wr_data_rom[21664]='h00000000;
    rd_cycle[21665] = 1'b1;  wr_cycle[21665] = 1'b0;  addr_rom[21665]='h00001284;  wr_data_rom[21665]='h00000000;
    rd_cycle[21666] = 1'b1;  wr_cycle[21666] = 1'b0;  addr_rom[21666]='h00001288;  wr_data_rom[21666]='h00000000;
    rd_cycle[21667] = 1'b1;  wr_cycle[21667] = 1'b0;  addr_rom[21667]='h0000128c;  wr_data_rom[21667]='h00000000;
    rd_cycle[21668] = 1'b1;  wr_cycle[21668] = 1'b0;  addr_rom[21668]='h00001290;  wr_data_rom[21668]='h00000000;
    rd_cycle[21669] = 1'b1;  wr_cycle[21669] = 1'b0;  addr_rom[21669]='h00001294;  wr_data_rom[21669]='h00000000;
    rd_cycle[21670] = 1'b1;  wr_cycle[21670] = 1'b0;  addr_rom[21670]='h00001298;  wr_data_rom[21670]='h00000000;
    rd_cycle[21671] = 1'b1;  wr_cycle[21671] = 1'b0;  addr_rom[21671]='h0000129c;  wr_data_rom[21671]='h00000000;
    rd_cycle[21672] = 1'b1;  wr_cycle[21672] = 1'b0;  addr_rom[21672]='h000012a0;  wr_data_rom[21672]='h00000000;
    rd_cycle[21673] = 1'b1;  wr_cycle[21673] = 1'b0;  addr_rom[21673]='h000012a4;  wr_data_rom[21673]='h00000000;
    rd_cycle[21674] = 1'b1;  wr_cycle[21674] = 1'b0;  addr_rom[21674]='h000012a8;  wr_data_rom[21674]='h00000000;
    rd_cycle[21675] = 1'b1;  wr_cycle[21675] = 1'b0;  addr_rom[21675]='h000012ac;  wr_data_rom[21675]='h00000000;
    rd_cycle[21676] = 1'b1;  wr_cycle[21676] = 1'b0;  addr_rom[21676]='h000012b0;  wr_data_rom[21676]='h00000000;
    rd_cycle[21677] = 1'b1;  wr_cycle[21677] = 1'b0;  addr_rom[21677]='h000012b4;  wr_data_rom[21677]='h00000000;
    rd_cycle[21678] = 1'b1;  wr_cycle[21678] = 1'b0;  addr_rom[21678]='h000012b8;  wr_data_rom[21678]='h00000000;
    rd_cycle[21679] = 1'b1;  wr_cycle[21679] = 1'b0;  addr_rom[21679]='h000012bc;  wr_data_rom[21679]='h00000000;
    rd_cycle[21680] = 1'b1;  wr_cycle[21680] = 1'b0;  addr_rom[21680]='h000012c0;  wr_data_rom[21680]='h00000000;
    rd_cycle[21681] = 1'b1;  wr_cycle[21681] = 1'b0;  addr_rom[21681]='h000012c4;  wr_data_rom[21681]='h00000000;
    rd_cycle[21682] = 1'b1;  wr_cycle[21682] = 1'b0;  addr_rom[21682]='h000012c8;  wr_data_rom[21682]='h00000000;
    rd_cycle[21683] = 1'b1;  wr_cycle[21683] = 1'b0;  addr_rom[21683]='h000012cc;  wr_data_rom[21683]='h00000000;
    rd_cycle[21684] = 1'b1;  wr_cycle[21684] = 1'b0;  addr_rom[21684]='h000012d0;  wr_data_rom[21684]='h00000000;
    rd_cycle[21685] = 1'b1;  wr_cycle[21685] = 1'b0;  addr_rom[21685]='h000012d4;  wr_data_rom[21685]='h00000000;
    rd_cycle[21686] = 1'b1;  wr_cycle[21686] = 1'b0;  addr_rom[21686]='h000012d8;  wr_data_rom[21686]='h00000000;
    rd_cycle[21687] = 1'b1;  wr_cycle[21687] = 1'b0;  addr_rom[21687]='h000012dc;  wr_data_rom[21687]='h00000000;
    rd_cycle[21688] = 1'b1;  wr_cycle[21688] = 1'b0;  addr_rom[21688]='h000012e0;  wr_data_rom[21688]='h00000000;
    rd_cycle[21689] = 1'b1;  wr_cycle[21689] = 1'b0;  addr_rom[21689]='h000012e4;  wr_data_rom[21689]='h00000000;
    rd_cycle[21690] = 1'b1;  wr_cycle[21690] = 1'b0;  addr_rom[21690]='h000012e8;  wr_data_rom[21690]='h00000000;
    rd_cycle[21691] = 1'b1;  wr_cycle[21691] = 1'b0;  addr_rom[21691]='h000012ec;  wr_data_rom[21691]='h00000000;
    rd_cycle[21692] = 1'b1;  wr_cycle[21692] = 1'b0;  addr_rom[21692]='h000012f0;  wr_data_rom[21692]='h00000000;
    rd_cycle[21693] = 1'b1;  wr_cycle[21693] = 1'b0;  addr_rom[21693]='h000012f4;  wr_data_rom[21693]='h00000000;
    rd_cycle[21694] = 1'b1;  wr_cycle[21694] = 1'b0;  addr_rom[21694]='h000012f8;  wr_data_rom[21694]='h00000000;
    rd_cycle[21695] = 1'b1;  wr_cycle[21695] = 1'b0;  addr_rom[21695]='h000012fc;  wr_data_rom[21695]='h00000000;
    rd_cycle[21696] = 1'b1;  wr_cycle[21696] = 1'b0;  addr_rom[21696]='h00001300;  wr_data_rom[21696]='h00000000;
    rd_cycle[21697] = 1'b1;  wr_cycle[21697] = 1'b0;  addr_rom[21697]='h00001304;  wr_data_rom[21697]='h00000000;
    rd_cycle[21698] = 1'b1;  wr_cycle[21698] = 1'b0;  addr_rom[21698]='h00001308;  wr_data_rom[21698]='h00000000;
    rd_cycle[21699] = 1'b1;  wr_cycle[21699] = 1'b0;  addr_rom[21699]='h0000130c;  wr_data_rom[21699]='h00000000;
    rd_cycle[21700] = 1'b1;  wr_cycle[21700] = 1'b0;  addr_rom[21700]='h00001310;  wr_data_rom[21700]='h00000000;
    rd_cycle[21701] = 1'b1;  wr_cycle[21701] = 1'b0;  addr_rom[21701]='h00001314;  wr_data_rom[21701]='h00000000;
    rd_cycle[21702] = 1'b1;  wr_cycle[21702] = 1'b0;  addr_rom[21702]='h00001318;  wr_data_rom[21702]='h00000000;
    rd_cycle[21703] = 1'b1;  wr_cycle[21703] = 1'b0;  addr_rom[21703]='h0000131c;  wr_data_rom[21703]='h00000000;
    rd_cycle[21704] = 1'b1;  wr_cycle[21704] = 1'b0;  addr_rom[21704]='h00001320;  wr_data_rom[21704]='h00000000;
    rd_cycle[21705] = 1'b1;  wr_cycle[21705] = 1'b0;  addr_rom[21705]='h00001324;  wr_data_rom[21705]='h00000000;
    rd_cycle[21706] = 1'b1;  wr_cycle[21706] = 1'b0;  addr_rom[21706]='h00001328;  wr_data_rom[21706]='h00000000;
    rd_cycle[21707] = 1'b1;  wr_cycle[21707] = 1'b0;  addr_rom[21707]='h0000132c;  wr_data_rom[21707]='h00000000;
    rd_cycle[21708] = 1'b1;  wr_cycle[21708] = 1'b0;  addr_rom[21708]='h00001330;  wr_data_rom[21708]='h00000000;
    rd_cycle[21709] = 1'b1;  wr_cycle[21709] = 1'b0;  addr_rom[21709]='h00001334;  wr_data_rom[21709]='h00000000;
    rd_cycle[21710] = 1'b1;  wr_cycle[21710] = 1'b0;  addr_rom[21710]='h00001338;  wr_data_rom[21710]='h00000000;
    rd_cycle[21711] = 1'b1;  wr_cycle[21711] = 1'b0;  addr_rom[21711]='h0000133c;  wr_data_rom[21711]='h00000000;
    rd_cycle[21712] = 1'b1;  wr_cycle[21712] = 1'b0;  addr_rom[21712]='h00001340;  wr_data_rom[21712]='h00000000;
    rd_cycle[21713] = 1'b1;  wr_cycle[21713] = 1'b0;  addr_rom[21713]='h00001344;  wr_data_rom[21713]='h00000000;
    rd_cycle[21714] = 1'b1;  wr_cycle[21714] = 1'b0;  addr_rom[21714]='h00001348;  wr_data_rom[21714]='h00000000;
    rd_cycle[21715] = 1'b1;  wr_cycle[21715] = 1'b0;  addr_rom[21715]='h0000134c;  wr_data_rom[21715]='h00000000;
    rd_cycle[21716] = 1'b1;  wr_cycle[21716] = 1'b0;  addr_rom[21716]='h00001350;  wr_data_rom[21716]='h00000000;
    rd_cycle[21717] = 1'b1;  wr_cycle[21717] = 1'b0;  addr_rom[21717]='h00001354;  wr_data_rom[21717]='h00000000;
    rd_cycle[21718] = 1'b1;  wr_cycle[21718] = 1'b0;  addr_rom[21718]='h00001358;  wr_data_rom[21718]='h00000000;
    rd_cycle[21719] = 1'b1;  wr_cycle[21719] = 1'b0;  addr_rom[21719]='h0000135c;  wr_data_rom[21719]='h00000000;
    rd_cycle[21720] = 1'b1;  wr_cycle[21720] = 1'b0;  addr_rom[21720]='h00001360;  wr_data_rom[21720]='h00000000;
    rd_cycle[21721] = 1'b1;  wr_cycle[21721] = 1'b0;  addr_rom[21721]='h00001364;  wr_data_rom[21721]='h00000000;
    rd_cycle[21722] = 1'b1;  wr_cycle[21722] = 1'b0;  addr_rom[21722]='h00001368;  wr_data_rom[21722]='h00000000;
    rd_cycle[21723] = 1'b1;  wr_cycle[21723] = 1'b0;  addr_rom[21723]='h0000136c;  wr_data_rom[21723]='h00000000;
    rd_cycle[21724] = 1'b1;  wr_cycle[21724] = 1'b0;  addr_rom[21724]='h00001370;  wr_data_rom[21724]='h00000000;
    rd_cycle[21725] = 1'b1;  wr_cycle[21725] = 1'b0;  addr_rom[21725]='h00001374;  wr_data_rom[21725]='h00000000;
    rd_cycle[21726] = 1'b1;  wr_cycle[21726] = 1'b0;  addr_rom[21726]='h00001378;  wr_data_rom[21726]='h00000000;
    rd_cycle[21727] = 1'b1;  wr_cycle[21727] = 1'b0;  addr_rom[21727]='h0000137c;  wr_data_rom[21727]='h00000000;
    rd_cycle[21728] = 1'b1;  wr_cycle[21728] = 1'b0;  addr_rom[21728]='h00001380;  wr_data_rom[21728]='h00000000;
    rd_cycle[21729] = 1'b1;  wr_cycle[21729] = 1'b0;  addr_rom[21729]='h00001384;  wr_data_rom[21729]='h00000000;
    rd_cycle[21730] = 1'b1;  wr_cycle[21730] = 1'b0;  addr_rom[21730]='h00001388;  wr_data_rom[21730]='h00000000;
    rd_cycle[21731] = 1'b1;  wr_cycle[21731] = 1'b0;  addr_rom[21731]='h0000138c;  wr_data_rom[21731]='h00000000;
    rd_cycle[21732] = 1'b1;  wr_cycle[21732] = 1'b0;  addr_rom[21732]='h00001390;  wr_data_rom[21732]='h00000000;
    rd_cycle[21733] = 1'b1;  wr_cycle[21733] = 1'b0;  addr_rom[21733]='h00001394;  wr_data_rom[21733]='h00000000;
    rd_cycle[21734] = 1'b1;  wr_cycle[21734] = 1'b0;  addr_rom[21734]='h00001398;  wr_data_rom[21734]='h00000000;
    rd_cycle[21735] = 1'b1;  wr_cycle[21735] = 1'b0;  addr_rom[21735]='h0000139c;  wr_data_rom[21735]='h00000000;
    rd_cycle[21736] = 1'b1;  wr_cycle[21736] = 1'b0;  addr_rom[21736]='h000013a0;  wr_data_rom[21736]='h00000000;
    rd_cycle[21737] = 1'b1;  wr_cycle[21737] = 1'b0;  addr_rom[21737]='h000013a4;  wr_data_rom[21737]='h00000000;
    rd_cycle[21738] = 1'b1;  wr_cycle[21738] = 1'b0;  addr_rom[21738]='h000013a8;  wr_data_rom[21738]='h00000000;
    rd_cycle[21739] = 1'b1;  wr_cycle[21739] = 1'b0;  addr_rom[21739]='h000013ac;  wr_data_rom[21739]='h00000000;
    rd_cycle[21740] = 1'b1;  wr_cycle[21740] = 1'b0;  addr_rom[21740]='h000013b0;  wr_data_rom[21740]='h00000000;
    rd_cycle[21741] = 1'b1;  wr_cycle[21741] = 1'b0;  addr_rom[21741]='h000013b4;  wr_data_rom[21741]='h00000000;
    rd_cycle[21742] = 1'b1;  wr_cycle[21742] = 1'b0;  addr_rom[21742]='h000013b8;  wr_data_rom[21742]='h00000000;
    rd_cycle[21743] = 1'b1;  wr_cycle[21743] = 1'b0;  addr_rom[21743]='h000013bc;  wr_data_rom[21743]='h00000000;
    rd_cycle[21744] = 1'b1;  wr_cycle[21744] = 1'b0;  addr_rom[21744]='h000013c0;  wr_data_rom[21744]='h00000000;
    rd_cycle[21745] = 1'b1;  wr_cycle[21745] = 1'b0;  addr_rom[21745]='h000013c4;  wr_data_rom[21745]='h00000000;
    rd_cycle[21746] = 1'b1;  wr_cycle[21746] = 1'b0;  addr_rom[21746]='h000013c8;  wr_data_rom[21746]='h00000000;
    rd_cycle[21747] = 1'b1;  wr_cycle[21747] = 1'b0;  addr_rom[21747]='h000013cc;  wr_data_rom[21747]='h00000000;
    rd_cycle[21748] = 1'b1;  wr_cycle[21748] = 1'b0;  addr_rom[21748]='h000013d0;  wr_data_rom[21748]='h00000000;
    rd_cycle[21749] = 1'b1;  wr_cycle[21749] = 1'b0;  addr_rom[21749]='h000013d4;  wr_data_rom[21749]='h00000000;
    rd_cycle[21750] = 1'b1;  wr_cycle[21750] = 1'b0;  addr_rom[21750]='h000013d8;  wr_data_rom[21750]='h00000000;
    rd_cycle[21751] = 1'b1;  wr_cycle[21751] = 1'b0;  addr_rom[21751]='h000013dc;  wr_data_rom[21751]='h00000000;
    rd_cycle[21752] = 1'b1;  wr_cycle[21752] = 1'b0;  addr_rom[21752]='h000013e0;  wr_data_rom[21752]='h00000000;
    rd_cycle[21753] = 1'b1;  wr_cycle[21753] = 1'b0;  addr_rom[21753]='h000013e4;  wr_data_rom[21753]='h00000000;
    rd_cycle[21754] = 1'b1;  wr_cycle[21754] = 1'b0;  addr_rom[21754]='h000013e8;  wr_data_rom[21754]='h00000000;
    rd_cycle[21755] = 1'b1;  wr_cycle[21755] = 1'b0;  addr_rom[21755]='h000013ec;  wr_data_rom[21755]='h00000000;
    rd_cycle[21756] = 1'b1;  wr_cycle[21756] = 1'b0;  addr_rom[21756]='h000013f0;  wr_data_rom[21756]='h00000000;
    rd_cycle[21757] = 1'b1;  wr_cycle[21757] = 1'b0;  addr_rom[21757]='h000013f4;  wr_data_rom[21757]='h00000000;
    rd_cycle[21758] = 1'b1;  wr_cycle[21758] = 1'b0;  addr_rom[21758]='h000013f8;  wr_data_rom[21758]='h00000000;
    rd_cycle[21759] = 1'b1;  wr_cycle[21759] = 1'b0;  addr_rom[21759]='h000013fc;  wr_data_rom[21759]='h00000000;
    rd_cycle[21760] = 1'b1;  wr_cycle[21760] = 1'b0;  addr_rom[21760]='h00001400;  wr_data_rom[21760]='h00000000;
    rd_cycle[21761] = 1'b1;  wr_cycle[21761] = 1'b0;  addr_rom[21761]='h00001404;  wr_data_rom[21761]='h00000000;
    rd_cycle[21762] = 1'b1;  wr_cycle[21762] = 1'b0;  addr_rom[21762]='h00001408;  wr_data_rom[21762]='h00000000;
    rd_cycle[21763] = 1'b1;  wr_cycle[21763] = 1'b0;  addr_rom[21763]='h0000140c;  wr_data_rom[21763]='h00000000;
    rd_cycle[21764] = 1'b1;  wr_cycle[21764] = 1'b0;  addr_rom[21764]='h00001410;  wr_data_rom[21764]='h00000000;
    rd_cycle[21765] = 1'b1;  wr_cycle[21765] = 1'b0;  addr_rom[21765]='h00001414;  wr_data_rom[21765]='h00000000;
    rd_cycle[21766] = 1'b1;  wr_cycle[21766] = 1'b0;  addr_rom[21766]='h00001418;  wr_data_rom[21766]='h00000000;
    rd_cycle[21767] = 1'b1;  wr_cycle[21767] = 1'b0;  addr_rom[21767]='h0000141c;  wr_data_rom[21767]='h00000000;
    rd_cycle[21768] = 1'b1;  wr_cycle[21768] = 1'b0;  addr_rom[21768]='h00001420;  wr_data_rom[21768]='h00000000;
    rd_cycle[21769] = 1'b1;  wr_cycle[21769] = 1'b0;  addr_rom[21769]='h00001424;  wr_data_rom[21769]='h00000000;
    rd_cycle[21770] = 1'b1;  wr_cycle[21770] = 1'b0;  addr_rom[21770]='h00001428;  wr_data_rom[21770]='h00000000;
    rd_cycle[21771] = 1'b1;  wr_cycle[21771] = 1'b0;  addr_rom[21771]='h0000142c;  wr_data_rom[21771]='h00000000;
    rd_cycle[21772] = 1'b1;  wr_cycle[21772] = 1'b0;  addr_rom[21772]='h00001430;  wr_data_rom[21772]='h00000000;
    rd_cycle[21773] = 1'b1;  wr_cycle[21773] = 1'b0;  addr_rom[21773]='h00001434;  wr_data_rom[21773]='h00000000;
    rd_cycle[21774] = 1'b1;  wr_cycle[21774] = 1'b0;  addr_rom[21774]='h00001438;  wr_data_rom[21774]='h00000000;
    rd_cycle[21775] = 1'b1;  wr_cycle[21775] = 1'b0;  addr_rom[21775]='h0000143c;  wr_data_rom[21775]='h00000000;
    rd_cycle[21776] = 1'b1;  wr_cycle[21776] = 1'b0;  addr_rom[21776]='h00001440;  wr_data_rom[21776]='h00000000;
    rd_cycle[21777] = 1'b1;  wr_cycle[21777] = 1'b0;  addr_rom[21777]='h00001444;  wr_data_rom[21777]='h00000000;
    rd_cycle[21778] = 1'b1;  wr_cycle[21778] = 1'b0;  addr_rom[21778]='h00001448;  wr_data_rom[21778]='h00000000;
    rd_cycle[21779] = 1'b1;  wr_cycle[21779] = 1'b0;  addr_rom[21779]='h0000144c;  wr_data_rom[21779]='h00000000;
    rd_cycle[21780] = 1'b1;  wr_cycle[21780] = 1'b0;  addr_rom[21780]='h00001450;  wr_data_rom[21780]='h00000000;
    rd_cycle[21781] = 1'b1;  wr_cycle[21781] = 1'b0;  addr_rom[21781]='h00001454;  wr_data_rom[21781]='h00000000;
    rd_cycle[21782] = 1'b1;  wr_cycle[21782] = 1'b0;  addr_rom[21782]='h00001458;  wr_data_rom[21782]='h00000000;
    rd_cycle[21783] = 1'b1;  wr_cycle[21783] = 1'b0;  addr_rom[21783]='h0000145c;  wr_data_rom[21783]='h00000000;
    rd_cycle[21784] = 1'b1;  wr_cycle[21784] = 1'b0;  addr_rom[21784]='h00001460;  wr_data_rom[21784]='h00000000;
    rd_cycle[21785] = 1'b1;  wr_cycle[21785] = 1'b0;  addr_rom[21785]='h00001464;  wr_data_rom[21785]='h00000000;
    rd_cycle[21786] = 1'b1;  wr_cycle[21786] = 1'b0;  addr_rom[21786]='h00001468;  wr_data_rom[21786]='h00000000;
    rd_cycle[21787] = 1'b1;  wr_cycle[21787] = 1'b0;  addr_rom[21787]='h0000146c;  wr_data_rom[21787]='h00000000;
    rd_cycle[21788] = 1'b1;  wr_cycle[21788] = 1'b0;  addr_rom[21788]='h00001470;  wr_data_rom[21788]='h00000000;
    rd_cycle[21789] = 1'b1;  wr_cycle[21789] = 1'b0;  addr_rom[21789]='h00001474;  wr_data_rom[21789]='h00000000;
    rd_cycle[21790] = 1'b1;  wr_cycle[21790] = 1'b0;  addr_rom[21790]='h00001478;  wr_data_rom[21790]='h00000000;
    rd_cycle[21791] = 1'b1;  wr_cycle[21791] = 1'b0;  addr_rom[21791]='h0000147c;  wr_data_rom[21791]='h00000000;
    rd_cycle[21792] = 1'b1;  wr_cycle[21792] = 1'b0;  addr_rom[21792]='h00001480;  wr_data_rom[21792]='h00000000;
    rd_cycle[21793] = 1'b1;  wr_cycle[21793] = 1'b0;  addr_rom[21793]='h00001484;  wr_data_rom[21793]='h00000000;
    rd_cycle[21794] = 1'b1;  wr_cycle[21794] = 1'b0;  addr_rom[21794]='h00001488;  wr_data_rom[21794]='h00000000;
    rd_cycle[21795] = 1'b1;  wr_cycle[21795] = 1'b0;  addr_rom[21795]='h0000148c;  wr_data_rom[21795]='h00000000;
    rd_cycle[21796] = 1'b1;  wr_cycle[21796] = 1'b0;  addr_rom[21796]='h00001490;  wr_data_rom[21796]='h00000000;
    rd_cycle[21797] = 1'b1;  wr_cycle[21797] = 1'b0;  addr_rom[21797]='h00001494;  wr_data_rom[21797]='h00000000;
    rd_cycle[21798] = 1'b1;  wr_cycle[21798] = 1'b0;  addr_rom[21798]='h00001498;  wr_data_rom[21798]='h00000000;
    rd_cycle[21799] = 1'b1;  wr_cycle[21799] = 1'b0;  addr_rom[21799]='h0000149c;  wr_data_rom[21799]='h00000000;
    rd_cycle[21800] = 1'b1;  wr_cycle[21800] = 1'b0;  addr_rom[21800]='h000014a0;  wr_data_rom[21800]='h00000000;
    rd_cycle[21801] = 1'b1;  wr_cycle[21801] = 1'b0;  addr_rom[21801]='h000014a4;  wr_data_rom[21801]='h00000000;
    rd_cycle[21802] = 1'b1;  wr_cycle[21802] = 1'b0;  addr_rom[21802]='h000014a8;  wr_data_rom[21802]='h00000000;
    rd_cycle[21803] = 1'b1;  wr_cycle[21803] = 1'b0;  addr_rom[21803]='h000014ac;  wr_data_rom[21803]='h00000000;
    rd_cycle[21804] = 1'b1;  wr_cycle[21804] = 1'b0;  addr_rom[21804]='h000014b0;  wr_data_rom[21804]='h00000000;
    rd_cycle[21805] = 1'b1;  wr_cycle[21805] = 1'b0;  addr_rom[21805]='h000014b4;  wr_data_rom[21805]='h00000000;
    rd_cycle[21806] = 1'b1;  wr_cycle[21806] = 1'b0;  addr_rom[21806]='h000014b8;  wr_data_rom[21806]='h00000000;
    rd_cycle[21807] = 1'b1;  wr_cycle[21807] = 1'b0;  addr_rom[21807]='h000014bc;  wr_data_rom[21807]='h00000000;
    rd_cycle[21808] = 1'b1;  wr_cycle[21808] = 1'b0;  addr_rom[21808]='h000014c0;  wr_data_rom[21808]='h00000000;
    rd_cycle[21809] = 1'b1;  wr_cycle[21809] = 1'b0;  addr_rom[21809]='h000014c4;  wr_data_rom[21809]='h00000000;
    rd_cycle[21810] = 1'b1;  wr_cycle[21810] = 1'b0;  addr_rom[21810]='h000014c8;  wr_data_rom[21810]='h00000000;
    rd_cycle[21811] = 1'b1;  wr_cycle[21811] = 1'b0;  addr_rom[21811]='h000014cc;  wr_data_rom[21811]='h00000000;
    rd_cycle[21812] = 1'b1;  wr_cycle[21812] = 1'b0;  addr_rom[21812]='h000014d0;  wr_data_rom[21812]='h00000000;
    rd_cycle[21813] = 1'b1;  wr_cycle[21813] = 1'b0;  addr_rom[21813]='h000014d4;  wr_data_rom[21813]='h00000000;
    rd_cycle[21814] = 1'b1;  wr_cycle[21814] = 1'b0;  addr_rom[21814]='h000014d8;  wr_data_rom[21814]='h00000000;
    rd_cycle[21815] = 1'b1;  wr_cycle[21815] = 1'b0;  addr_rom[21815]='h000014dc;  wr_data_rom[21815]='h00000000;
    rd_cycle[21816] = 1'b1;  wr_cycle[21816] = 1'b0;  addr_rom[21816]='h000014e0;  wr_data_rom[21816]='h00000000;
    rd_cycle[21817] = 1'b1;  wr_cycle[21817] = 1'b0;  addr_rom[21817]='h000014e4;  wr_data_rom[21817]='h00000000;
    rd_cycle[21818] = 1'b1;  wr_cycle[21818] = 1'b0;  addr_rom[21818]='h000014e8;  wr_data_rom[21818]='h00000000;
    rd_cycle[21819] = 1'b1;  wr_cycle[21819] = 1'b0;  addr_rom[21819]='h000014ec;  wr_data_rom[21819]='h00000000;
    rd_cycle[21820] = 1'b1;  wr_cycle[21820] = 1'b0;  addr_rom[21820]='h000014f0;  wr_data_rom[21820]='h00000000;
    rd_cycle[21821] = 1'b1;  wr_cycle[21821] = 1'b0;  addr_rom[21821]='h000014f4;  wr_data_rom[21821]='h00000000;
    rd_cycle[21822] = 1'b1;  wr_cycle[21822] = 1'b0;  addr_rom[21822]='h000014f8;  wr_data_rom[21822]='h00000000;
    rd_cycle[21823] = 1'b1;  wr_cycle[21823] = 1'b0;  addr_rom[21823]='h000014fc;  wr_data_rom[21823]='h00000000;
    rd_cycle[21824] = 1'b1;  wr_cycle[21824] = 1'b0;  addr_rom[21824]='h00001500;  wr_data_rom[21824]='h00000000;
    rd_cycle[21825] = 1'b1;  wr_cycle[21825] = 1'b0;  addr_rom[21825]='h00001504;  wr_data_rom[21825]='h00000000;
    rd_cycle[21826] = 1'b1;  wr_cycle[21826] = 1'b0;  addr_rom[21826]='h00001508;  wr_data_rom[21826]='h00000000;
    rd_cycle[21827] = 1'b1;  wr_cycle[21827] = 1'b0;  addr_rom[21827]='h0000150c;  wr_data_rom[21827]='h00000000;
    rd_cycle[21828] = 1'b1;  wr_cycle[21828] = 1'b0;  addr_rom[21828]='h00001510;  wr_data_rom[21828]='h00000000;
    rd_cycle[21829] = 1'b1;  wr_cycle[21829] = 1'b0;  addr_rom[21829]='h00001514;  wr_data_rom[21829]='h00000000;
    rd_cycle[21830] = 1'b1;  wr_cycle[21830] = 1'b0;  addr_rom[21830]='h00001518;  wr_data_rom[21830]='h00000000;
    rd_cycle[21831] = 1'b1;  wr_cycle[21831] = 1'b0;  addr_rom[21831]='h0000151c;  wr_data_rom[21831]='h00000000;
    rd_cycle[21832] = 1'b1;  wr_cycle[21832] = 1'b0;  addr_rom[21832]='h00001520;  wr_data_rom[21832]='h00000000;
    rd_cycle[21833] = 1'b1;  wr_cycle[21833] = 1'b0;  addr_rom[21833]='h00001524;  wr_data_rom[21833]='h00000000;
    rd_cycle[21834] = 1'b1;  wr_cycle[21834] = 1'b0;  addr_rom[21834]='h00001528;  wr_data_rom[21834]='h00000000;
    rd_cycle[21835] = 1'b1;  wr_cycle[21835] = 1'b0;  addr_rom[21835]='h0000152c;  wr_data_rom[21835]='h00000000;
    rd_cycle[21836] = 1'b1;  wr_cycle[21836] = 1'b0;  addr_rom[21836]='h00001530;  wr_data_rom[21836]='h00000000;
    rd_cycle[21837] = 1'b1;  wr_cycle[21837] = 1'b0;  addr_rom[21837]='h00001534;  wr_data_rom[21837]='h00000000;
    rd_cycle[21838] = 1'b1;  wr_cycle[21838] = 1'b0;  addr_rom[21838]='h00001538;  wr_data_rom[21838]='h00000000;
    rd_cycle[21839] = 1'b1;  wr_cycle[21839] = 1'b0;  addr_rom[21839]='h0000153c;  wr_data_rom[21839]='h00000000;
    rd_cycle[21840] = 1'b1;  wr_cycle[21840] = 1'b0;  addr_rom[21840]='h00001540;  wr_data_rom[21840]='h00000000;
    rd_cycle[21841] = 1'b1;  wr_cycle[21841] = 1'b0;  addr_rom[21841]='h00001544;  wr_data_rom[21841]='h00000000;
    rd_cycle[21842] = 1'b1;  wr_cycle[21842] = 1'b0;  addr_rom[21842]='h00001548;  wr_data_rom[21842]='h00000000;
    rd_cycle[21843] = 1'b1;  wr_cycle[21843] = 1'b0;  addr_rom[21843]='h0000154c;  wr_data_rom[21843]='h00000000;
    rd_cycle[21844] = 1'b1;  wr_cycle[21844] = 1'b0;  addr_rom[21844]='h00001550;  wr_data_rom[21844]='h00000000;
    rd_cycle[21845] = 1'b1;  wr_cycle[21845] = 1'b0;  addr_rom[21845]='h00001554;  wr_data_rom[21845]='h00000000;
    rd_cycle[21846] = 1'b1;  wr_cycle[21846] = 1'b0;  addr_rom[21846]='h00001558;  wr_data_rom[21846]='h00000000;
    rd_cycle[21847] = 1'b1;  wr_cycle[21847] = 1'b0;  addr_rom[21847]='h0000155c;  wr_data_rom[21847]='h00000000;
    rd_cycle[21848] = 1'b1;  wr_cycle[21848] = 1'b0;  addr_rom[21848]='h00001560;  wr_data_rom[21848]='h00000000;
    rd_cycle[21849] = 1'b1;  wr_cycle[21849] = 1'b0;  addr_rom[21849]='h00001564;  wr_data_rom[21849]='h00000000;
    rd_cycle[21850] = 1'b1;  wr_cycle[21850] = 1'b0;  addr_rom[21850]='h00001568;  wr_data_rom[21850]='h00000000;
    rd_cycle[21851] = 1'b1;  wr_cycle[21851] = 1'b0;  addr_rom[21851]='h0000156c;  wr_data_rom[21851]='h00000000;
    rd_cycle[21852] = 1'b1;  wr_cycle[21852] = 1'b0;  addr_rom[21852]='h00001570;  wr_data_rom[21852]='h00000000;
    rd_cycle[21853] = 1'b1;  wr_cycle[21853] = 1'b0;  addr_rom[21853]='h00001574;  wr_data_rom[21853]='h00000000;
    rd_cycle[21854] = 1'b1;  wr_cycle[21854] = 1'b0;  addr_rom[21854]='h00001578;  wr_data_rom[21854]='h00000000;
    rd_cycle[21855] = 1'b1;  wr_cycle[21855] = 1'b0;  addr_rom[21855]='h0000157c;  wr_data_rom[21855]='h00000000;
    rd_cycle[21856] = 1'b1;  wr_cycle[21856] = 1'b0;  addr_rom[21856]='h00001580;  wr_data_rom[21856]='h00000000;
    rd_cycle[21857] = 1'b1;  wr_cycle[21857] = 1'b0;  addr_rom[21857]='h00001584;  wr_data_rom[21857]='h00000000;
    rd_cycle[21858] = 1'b1;  wr_cycle[21858] = 1'b0;  addr_rom[21858]='h00001588;  wr_data_rom[21858]='h00000000;
    rd_cycle[21859] = 1'b1;  wr_cycle[21859] = 1'b0;  addr_rom[21859]='h0000158c;  wr_data_rom[21859]='h00000000;
    rd_cycle[21860] = 1'b1;  wr_cycle[21860] = 1'b0;  addr_rom[21860]='h00001590;  wr_data_rom[21860]='h00000000;
    rd_cycle[21861] = 1'b1;  wr_cycle[21861] = 1'b0;  addr_rom[21861]='h00001594;  wr_data_rom[21861]='h00000000;
    rd_cycle[21862] = 1'b1;  wr_cycle[21862] = 1'b0;  addr_rom[21862]='h00001598;  wr_data_rom[21862]='h00000000;
    rd_cycle[21863] = 1'b1;  wr_cycle[21863] = 1'b0;  addr_rom[21863]='h0000159c;  wr_data_rom[21863]='h00000000;
    rd_cycle[21864] = 1'b1;  wr_cycle[21864] = 1'b0;  addr_rom[21864]='h000015a0;  wr_data_rom[21864]='h00000000;
    rd_cycle[21865] = 1'b1;  wr_cycle[21865] = 1'b0;  addr_rom[21865]='h000015a4;  wr_data_rom[21865]='h00000000;
    rd_cycle[21866] = 1'b1;  wr_cycle[21866] = 1'b0;  addr_rom[21866]='h000015a8;  wr_data_rom[21866]='h00000000;
    rd_cycle[21867] = 1'b1;  wr_cycle[21867] = 1'b0;  addr_rom[21867]='h000015ac;  wr_data_rom[21867]='h00000000;
    rd_cycle[21868] = 1'b1;  wr_cycle[21868] = 1'b0;  addr_rom[21868]='h000015b0;  wr_data_rom[21868]='h00000000;
    rd_cycle[21869] = 1'b1;  wr_cycle[21869] = 1'b0;  addr_rom[21869]='h000015b4;  wr_data_rom[21869]='h00000000;
    rd_cycle[21870] = 1'b1;  wr_cycle[21870] = 1'b0;  addr_rom[21870]='h000015b8;  wr_data_rom[21870]='h00000000;
    rd_cycle[21871] = 1'b1;  wr_cycle[21871] = 1'b0;  addr_rom[21871]='h000015bc;  wr_data_rom[21871]='h00000000;
    rd_cycle[21872] = 1'b1;  wr_cycle[21872] = 1'b0;  addr_rom[21872]='h000015c0;  wr_data_rom[21872]='h00000000;
    rd_cycle[21873] = 1'b1;  wr_cycle[21873] = 1'b0;  addr_rom[21873]='h000015c4;  wr_data_rom[21873]='h00000000;
    rd_cycle[21874] = 1'b1;  wr_cycle[21874] = 1'b0;  addr_rom[21874]='h000015c8;  wr_data_rom[21874]='h00000000;
    rd_cycle[21875] = 1'b1;  wr_cycle[21875] = 1'b0;  addr_rom[21875]='h000015cc;  wr_data_rom[21875]='h00000000;
    rd_cycle[21876] = 1'b1;  wr_cycle[21876] = 1'b0;  addr_rom[21876]='h000015d0;  wr_data_rom[21876]='h00000000;
    rd_cycle[21877] = 1'b1;  wr_cycle[21877] = 1'b0;  addr_rom[21877]='h000015d4;  wr_data_rom[21877]='h00000000;
    rd_cycle[21878] = 1'b1;  wr_cycle[21878] = 1'b0;  addr_rom[21878]='h000015d8;  wr_data_rom[21878]='h00000000;
    rd_cycle[21879] = 1'b1;  wr_cycle[21879] = 1'b0;  addr_rom[21879]='h000015dc;  wr_data_rom[21879]='h00000000;
    rd_cycle[21880] = 1'b1;  wr_cycle[21880] = 1'b0;  addr_rom[21880]='h000015e0;  wr_data_rom[21880]='h00000000;
    rd_cycle[21881] = 1'b1;  wr_cycle[21881] = 1'b0;  addr_rom[21881]='h000015e4;  wr_data_rom[21881]='h00000000;
    rd_cycle[21882] = 1'b1;  wr_cycle[21882] = 1'b0;  addr_rom[21882]='h000015e8;  wr_data_rom[21882]='h00000000;
    rd_cycle[21883] = 1'b1;  wr_cycle[21883] = 1'b0;  addr_rom[21883]='h000015ec;  wr_data_rom[21883]='h00000000;
    rd_cycle[21884] = 1'b1;  wr_cycle[21884] = 1'b0;  addr_rom[21884]='h000015f0;  wr_data_rom[21884]='h00000000;
    rd_cycle[21885] = 1'b1;  wr_cycle[21885] = 1'b0;  addr_rom[21885]='h000015f4;  wr_data_rom[21885]='h00000000;
    rd_cycle[21886] = 1'b1;  wr_cycle[21886] = 1'b0;  addr_rom[21886]='h000015f8;  wr_data_rom[21886]='h00000000;
    rd_cycle[21887] = 1'b1;  wr_cycle[21887] = 1'b0;  addr_rom[21887]='h000015fc;  wr_data_rom[21887]='h00000000;
    rd_cycle[21888] = 1'b1;  wr_cycle[21888] = 1'b0;  addr_rom[21888]='h00001600;  wr_data_rom[21888]='h00000000;
    rd_cycle[21889] = 1'b1;  wr_cycle[21889] = 1'b0;  addr_rom[21889]='h00001604;  wr_data_rom[21889]='h00000000;
    rd_cycle[21890] = 1'b1;  wr_cycle[21890] = 1'b0;  addr_rom[21890]='h00001608;  wr_data_rom[21890]='h00000000;
    rd_cycle[21891] = 1'b1;  wr_cycle[21891] = 1'b0;  addr_rom[21891]='h0000160c;  wr_data_rom[21891]='h00000000;
    rd_cycle[21892] = 1'b1;  wr_cycle[21892] = 1'b0;  addr_rom[21892]='h00001610;  wr_data_rom[21892]='h00000000;
    rd_cycle[21893] = 1'b1;  wr_cycle[21893] = 1'b0;  addr_rom[21893]='h00001614;  wr_data_rom[21893]='h00000000;
    rd_cycle[21894] = 1'b1;  wr_cycle[21894] = 1'b0;  addr_rom[21894]='h00001618;  wr_data_rom[21894]='h00000000;
    rd_cycle[21895] = 1'b1;  wr_cycle[21895] = 1'b0;  addr_rom[21895]='h0000161c;  wr_data_rom[21895]='h00000000;
    rd_cycle[21896] = 1'b1;  wr_cycle[21896] = 1'b0;  addr_rom[21896]='h00001620;  wr_data_rom[21896]='h00000000;
    rd_cycle[21897] = 1'b1;  wr_cycle[21897] = 1'b0;  addr_rom[21897]='h00001624;  wr_data_rom[21897]='h00000000;
    rd_cycle[21898] = 1'b1;  wr_cycle[21898] = 1'b0;  addr_rom[21898]='h00001628;  wr_data_rom[21898]='h00000000;
    rd_cycle[21899] = 1'b1;  wr_cycle[21899] = 1'b0;  addr_rom[21899]='h0000162c;  wr_data_rom[21899]='h00000000;
    rd_cycle[21900] = 1'b1;  wr_cycle[21900] = 1'b0;  addr_rom[21900]='h00001630;  wr_data_rom[21900]='h00000000;
    rd_cycle[21901] = 1'b1;  wr_cycle[21901] = 1'b0;  addr_rom[21901]='h00001634;  wr_data_rom[21901]='h00000000;
    rd_cycle[21902] = 1'b1;  wr_cycle[21902] = 1'b0;  addr_rom[21902]='h00001638;  wr_data_rom[21902]='h00000000;
    rd_cycle[21903] = 1'b1;  wr_cycle[21903] = 1'b0;  addr_rom[21903]='h0000163c;  wr_data_rom[21903]='h00000000;
    rd_cycle[21904] = 1'b1;  wr_cycle[21904] = 1'b0;  addr_rom[21904]='h00001640;  wr_data_rom[21904]='h00000000;
    rd_cycle[21905] = 1'b1;  wr_cycle[21905] = 1'b0;  addr_rom[21905]='h00001644;  wr_data_rom[21905]='h00000000;
    rd_cycle[21906] = 1'b1;  wr_cycle[21906] = 1'b0;  addr_rom[21906]='h00001648;  wr_data_rom[21906]='h00000000;
    rd_cycle[21907] = 1'b1;  wr_cycle[21907] = 1'b0;  addr_rom[21907]='h0000164c;  wr_data_rom[21907]='h00000000;
    rd_cycle[21908] = 1'b1;  wr_cycle[21908] = 1'b0;  addr_rom[21908]='h00001650;  wr_data_rom[21908]='h00000000;
    rd_cycle[21909] = 1'b1;  wr_cycle[21909] = 1'b0;  addr_rom[21909]='h00001654;  wr_data_rom[21909]='h00000000;
    rd_cycle[21910] = 1'b1;  wr_cycle[21910] = 1'b0;  addr_rom[21910]='h00001658;  wr_data_rom[21910]='h00000000;
    rd_cycle[21911] = 1'b1;  wr_cycle[21911] = 1'b0;  addr_rom[21911]='h0000165c;  wr_data_rom[21911]='h00000000;
    rd_cycle[21912] = 1'b1;  wr_cycle[21912] = 1'b0;  addr_rom[21912]='h00001660;  wr_data_rom[21912]='h00000000;
    rd_cycle[21913] = 1'b1;  wr_cycle[21913] = 1'b0;  addr_rom[21913]='h00001664;  wr_data_rom[21913]='h00000000;
    rd_cycle[21914] = 1'b1;  wr_cycle[21914] = 1'b0;  addr_rom[21914]='h00001668;  wr_data_rom[21914]='h00000000;
    rd_cycle[21915] = 1'b1;  wr_cycle[21915] = 1'b0;  addr_rom[21915]='h0000166c;  wr_data_rom[21915]='h00000000;
    rd_cycle[21916] = 1'b1;  wr_cycle[21916] = 1'b0;  addr_rom[21916]='h00001670;  wr_data_rom[21916]='h00000000;
    rd_cycle[21917] = 1'b1;  wr_cycle[21917] = 1'b0;  addr_rom[21917]='h00001674;  wr_data_rom[21917]='h00000000;
    rd_cycle[21918] = 1'b1;  wr_cycle[21918] = 1'b0;  addr_rom[21918]='h00001678;  wr_data_rom[21918]='h00000000;
    rd_cycle[21919] = 1'b1;  wr_cycle[21919] = 1'b0;  addr_rom[21919]='h0000167c;  wr_data_rom[21919]='h00000000;
    rd_cycle[21920] = 1'b1;  wr_cycle[21920] = 1'b0;  addr_rom[21920]='h00001680;  wr_data_rom[21920]='h00000000;
    rd_cycle[21921] = 1'b1;  wr_cycle[21921] = 1'b0;  addr_rom[21921]='h00001684;  wr_data_rom[21921]='h00000000;
    rd_cycle[21922] = 1'b1;  wr_cycle[21922] = 1'b0;  addr_rom[21922]='h00001688;  wr_data_rom[21922]='h00000000;
    rd_cycle[21923] = 1'b1;  wr_cycle[21923] = 1'b0;  addr_rom[21923]='h0000168c;  wr_data_rom[21923]='h00000000;
    rd_cycle[21924] = 1'b1;  wr_cycle[21924] = 1'b0;  addr_rom[21924]='h00001690;  wr_data_rom[21924]='h00000000;
    rd_cycle[21925] = 1'b1;  wr_cycle[21925] = 1'b0;  addr_rom[21925]='h00001694;  wr_data_rom[21925]='h00000000;
    rd_cycle[21926] = 1'b1;  wr_cycle[21926] = 1'b0;  addr_rom[21926]='h00001698;  wr_data_rom[21926]='h00000000;
    rd_cycle[21927] = 1'b1;  wr_cycle[21927] = 1'b0;  addr_rom[21927]='h0000169c;  wr_data_rom[21927]='h00000000;
    rd_cycle[21928] = 1'b1;  wr_cycle[21928] = 1'b0;  addr_rom[21928]='h000016a0;  wr_data_rom[21928]='h00000000;
    rd_cycle[21929] = 1'b1;  wr_cycle[21929] = 1'b0;  addr_rom[21929]='h000016a4;  wr_data_rom[21929]='h00000000;
    rd_cycle[21930] = 1'b1;  wr_cycle[21930] = 1'b0;  addr_rom[21930]='h000016a8;  wr_data_rom[21930]='h00000000;
    rd_cycle[21931] = 1'b1;  wr_cycle[21931] = 1'b0;  addr_rom[21931]='h000016ac;  wr_data_rom[21931]='h00000000;
    rd_cycle[21932] = 1'b1;  wr_cycle[21932] = 1'b0;  addr_rom[21932]='h000016b0;  wr_data_rom[21932]='h00000000;
    rd_cycle[21933] = 1'b1;  wr_cycle[21933] = 1'b0;  addr_rom[21933]='h000016b4;  wr_data_rom[21933]='h00000000;
    rd_cycle[21934] = 1'b1;  wr_cycle[21934] = 1'b0;  addr_rom[21934]='h000016b8;  wr_data_rom[21934]='h00000000;
    rd_cycle[21935] = 1'b1;  wr_cycle[21935] = 1'b0;  addr_rom[21935]='h000016bc;  wr_data_rom[21935]='h00000000;
    rd_cycle[21936] = 1'b1;  wr_cycle[21936] = 1'b0;  addr_rom[21936]='h000016c0;  wr_data_rom[21936]='h00000000;
    rd_cycle[21937] = 1'b1;  wr_cycle[21937] = 1'b0;  addr_rom[21937]='h000016c4;  wr_data_rom[21937]='h00000000;
    rd_cycle[21938] = 1'b1;  wr_cycle[21938] = 1'b0;  addr_rom[21938]='h000016c8;  wr_data_rom[21938]='h00000000;
    rd_cycle[21939] = 1'b1;  wr_cycle[21939] = 1'b0;  addr_rom[21939]='h000016cc;  wr_data_rom[21939]='h00000000;
    rd_cycle[21940] = 1'b1;  wr_cycle[21940] = 1'b0;  addr_rom[21940]='h000016d0;  wr_data_rom[21940]='h00000000;
    rd_cycle[21941] = 1'b1;  wr_cycle[21941] = 1'b0;  addr_rom[21941]='h000016d4;  wr_data_rom[21941]='h00000000;
    rd_cycle[21942] = 1'b1;  wr_cycle[21942] = 1'b0;  addr_rom[21942]='h000016d8;  wr_data_rom[21942]='h00000000;
    rd_cycle[21943] = 1'b1;  wr_cycle[21943] = 1'b0;  addr_rom[21943]='h000016dc;  wr_data_rom[21943]='h00000000;
    rd_cycle[21944] = 1'b1;  wr_cycle[21944] = 1'b0;  addr_rom[21944]='h000016e0;  wr_data_rom[21944]='h00000000;
    rd_cycle[21945] = 1'b1;  wr_cycle[21945] = 1'b0;  addr_rom[21945]='h000016e4;  wr_data_rom[21945]='h00000000;
    rd_cycle[21946] = 1'b1;  wr_cycle[21946] = 1'b0;  addr_rom[21946]='h000016e8;  wr_data_rom[21946]='h00000000;
    rd_cycle[21947] = 1'b1;  wr_cycle[21947] = 1'b0;  addr_rom[21947]='h000016ec;  wr_data_rom[21947]='h00000000;
    rd_cycle[21948] = 1'b1;  wr_cycle[21948] = 1'b0;  addr_rom[21948]='h000016f0;  wr_data_rom[21948]='h00000000;
    rd_cycle[21949] = 1'b1;  wr_cycle[21949] = 1'b0;  addr_rom[21949]='h000016f4;  wr_data_rom[21949]='h00000000;
    rd_cycle[21950] = 1'b1;  wr_cycle[21950] = 1'b0;  addr_rom[21950]='h000016f8;  wr_data_rom[21950]='h00000000;
    rd_cycle[21951] = 1'b1;  wr_cycle[21951] = 1'b0;  addr_rom[21951]='h000016fc;  wr_data_rom[21951]='h00000000;
    rd_cycle[21952] = 1'b1;  wr_cycle[21952] = 1'b0;  addr_rom[21952]='h00001700;  wr_data_rom[21952]='h00000000;
    rd_cycle[21953] = 1'b1;  wr_cycle[21953] = 1'b0;  addr_rom[21953]='h00001704;  wr_data_rom[21953]='h00000000;
    rd_cycle[21954] = 1'b1;  wr_cycle[21954] = 1'b0;  addr_rom[21954]='h00001708;  wr_data_rom[21954]='h00000000;
    rd_cycle[21955] = 1'b1;  wr_cycle[21955] = 1'b0;  addr_rom[21955]='h0000170c;  wr_data_rom[21955]='h00000000;
    rd_cycle[21956] = 1'b1;  wr_cycle[21956] = 1'b0;  addr_rom[21956]='h00001710;  wr_data_rom[21956]='h00000000;
    rd_cycle[21957] = 1'b1;  wr_cycle[21957] = 1'b0;  addr_rom[21957]='h00001714;  wr_data_rom[21957]='h00000000;
    rd_cycle[21958] = 1'b1;  wr_cycle[21958] = 1'b0;  addr_rom[21958]='h00001718;  wr_data_rom[21958]='h00000000;
    rd_cycle[21959] = 1'b1;  wr_cycle[21959] = 1'b0;  addr_rom[21959]='h0000171c;  wr_data_rom[21959]='h00000000;
    rd_cycle[21960] = 1'b1;  wr_cycle[21960] = 1'b0;  addr_rom[21960]='h00001720;  wr_data_rom[21960]='h00000000;
    rd_cycle[21961] = 1'b1;  wr_cycle[21961] = 1'b0;  addr_rom[21961]='h00001724;  wr_data_rom[21961]='h00000000;
    rd_cycle[21962] = 1'b1;  wr_cycle[21962] = 1'b0;  addr_rom[21962]='h00001728;  wr_data_rom[21962]='h00000000;
    rd_cycle[21963] = 1'b1;  wr_cycle[21963] = 1'b0;  addr_rom[21963]='h0000172c;  wr_data_rom[21963]='h00000000;
    rd_cycle[21964] = 1'b1;  wr_cycle[21964] = 1'b0;  addr_rom[21964]='h00001730;  wr_data_rom[21964]='h00000000;
    rd_cycle[21965] = 1'b1;  wr_cycle[21965] = 1'b0;  addr_rom[21965]='h00001734;  wr_data_rom[21965]='h00000000;
    rd_cycle[21966] = 1'b1;  wr_cycle[21966] = 1'b0;  addr_rom[21966]='h00001738;  wr_data_rom[21966]='h00000000;
    rd_cycle[21967] = 1'b1;  wr_cycle[21967] = 1'b0;  addr_rom[21967]='h0000173c;  wr_data_rom[21967]='h00000000;
    rd_cycle[21968] = 1'b1;  wr_cycle[21968] = 1'b0;  addr_rom[21968]='h00001740;  wr_data_rom[21968]='h00000000;
    rd_cycle[21969] = 1'b1;  wr_cycle[21969] = 1'b0;  addr_rom[21969]='h00001744;  wr_data_rom[21969]='h00000000;
    rd_cycle[21970] = 1'b1;  wr_cycle[21970] = 1'b0;  addr_rom[21970]='h00001748;  wr_data_rom[21970]='h00000000;
    rd_cycle[21971] = 1'b1;  wr_cycle[21971] = 1'b0;  addr_rom[21971]='h0000174c;  wr_data_rom[21971]='h00000000;
    rd_cycle[21972] = 1'b1;  wr_cycle[21972] = 1'b0;  addr_rom[21972]='h00001750;  wr_data_rom[21972]='h00000000;
    rd_cycle[21973] = 1'b1;  wr_cycle[21973] = 1'b0;  addr_rom[21973]='h00001754;  wr_data_rom[21973]='h00000000;
    rd_cycle[21974] = 1'b1;  wr_cycle[21974] = 1'b0;  addr_rom[21974]='h00001758;  wr_data_rom[21974]='h00000000;
    rd_cycle[21975] = 1'b1;  wr_cycle[21975] = 1'b0;  addr_rom[21975]='h0000175c;  wr_data_rom[21975]='h00000000;
    rd_cycle[21976] = 1'b1;  wr_cycle[21976] = 1'b0;  addr_rom[21976]='h00001760;  wr_data_rom[21976]='h00000000;
    rd_cycle[21977] = 1'b1;  wr_cycle[21977] = 1'b0;  addr_rom[21977]='h00001764;  wr_data_rom[21977]='h00000000;
    rd_cycle[21978] = 1'b1;  wr_cycle[21978] = 1'b0;  addr_rom[21978]='h00001768;  wr_data_rom[21978]='h00000000;
    rd_cycle[21979] = 1'b1;  wr_cycle[21979] = 1'b0;  addr_rom[21979]='h0000176c;  wr_data_rom[21979]='h00000000;
    rd_cycle[21980] = 1'b1;  wr_cycle[21980] = 1'b0;  addr_rom[21980]='h00001770;  wr_data_rom[21980]='h00000000;
    rd_cycle[21981] = 1'b1;  wr_cycle[21981] = 1'b0;  addr_rom[21981]='h00001774;  wr_data_rom[21981]='h00000000;
    rd_cycle[21982] = 1'b1;  wr_cycle[21982] = 1'b0;  addr_rom[21982]='h00001778;  wr_data_rom[21982]='h00000000;
    rd_cycle[21983] = 1'b1;  wr_cycle[21983] = 1'b0;  addr_rom[21983]='h0000177c;  wr_data_rom[21983]='h00000000;
    rd_cycle[21984] = 1'b1;  wr_cycle[21984] = 1'b0;  addr_rom[21984]='h00001780;  wr_data_rom[21984]='h00000000;
    rd_cycle[21985] = 1'b1;  wr_cycle[21985] = 1'b0;  addr_rom[21985]='h00001784;  wr_data_rom[21985]='h00000000;
    rd_cycle[21986] = 1'b1;  wr_cycle[21986] = 1'b0;  addr_rom[21986]='h00001788;  wr_data_rom[21986]='h00000000;
    rd_cycle[21987] = 1'b1;  wr_cycle[21987] = 1'b0;  addr_rom[21987]='h0000178c;  wr_data_rom[21987]='h00000000;
    rd_cycle[21988] = 1'b1;  wr_cycle[21988] = 1'b0;  addr_rom[21988]='h00001790;  wr_data_rom[21988]='h00000000;
    rd_cycle[21989] = 1'b1;  wr_cycle[21989] = 1'b0;  addr_rom[21989]='h00001794;  wr_data_rom[21989]='h00000000;
    rd_cycle[21990] = 1'b1;  wr_cycle[21990] = 1'b0;  addr_rom[21990]='h00001798;  wr_data_rom[21990]='h00000000;
    rd_cycle[21991] = 1'b1;  wr_cycle[21991] = 1'b0;  addr_rom[21991]='h0000179c;  wr_data_rom[21991]='h00000000;
    rd_cycle[21992] = 1'b1;  wr_cycle[21992] = 1'b0;  addr_rom[21992]='h000017a0;  wr_data_rom[21992]='h00000000;
    rd_cycle[21993] = 1'b1;  wr_cycle[21993] = 1'b0;  addr_rom[21993]='h000017a4;  wr_data_rom[21993]='h00000000;
    rd_cycle[21994] = 1'b1;  wr_cycle[21994] = 1'b0;  addr_rom[21994]='h000017a8;  wr_data_rom[21994]='h00000000;
    rd_cycle[21995] = 1'b1;  wr_cycle[21995] = 1'b0;  addr_rom[21995]='h000017ac;  wr_data_rom[21995]='h00000000;
    rd_cycle[21996] = 1'b1;  wr_cycle[21996] = 1'b0;  addr_rom[21996]='h000017b0;  wr_data_rom[21996]='h00000000;
    rd_cycle[21997] = 1'b1;  wr_cycle[21997] = 1'b0;  addr_rom[21997]='h000017b4;  wr_data_rom[21997]='h00000000;
    rd_cycle[21998] = 1'b1;  wr_cycle[21998] = 1'b0;  addr_rom[21998]='h000017b8;  wr_data_rom[21998]='h00000000;
    rd_cycle[21999] = 1'b1;  wr_cycle[21999] = 1'b0;  addr_rom[21999]='h000017bc;  wr_data_rom[21999]='h00000000;
    rd_cycle[22000] = 1'b1;  wr_cycle[22000] = 1'b0;  addr_rom[22000]='h000017c0;  wr_data_rom[22000]='h00000000;
    rd_cycle[22001] = 1'b1;  wr_cycle[22001] = 1'b0;  addr_rom[22001]='h000017c4;  wr_data_rom[22001]='h00000000;
    rd_cycle[22002] = 1'b1;  wr_cycle[22002] = 1'b0;  addr_rom[22002]='h000017c8;  wr_data_rom[22002]='h00000000;
    rd_cycle[22003] = 1'b1;  wr_cycle[22003] = 1'b0;  addr_rom[22003]='h000017cc;  wr_data_rom[22003]='h00000000;
    rd_cycle[22004] = 1'b1;  wr_cycle[22004] = 1'b0;  addr_rom[22004]='h000017d0;  wr_data_rom[22004]='h00000000;
    rd_cycle[22005] = 1'b1;  wr_cycle[22005] = 1'b0;  addr_rom[22005]='h000017d4;  wr_data_rom[22005]='h00000000;
    rd_cycle[22006] = 1'b1;  wr_cycle[22006] = 1'b0;  addr_rom[22006]='h000017d8;  wr_data_rom[22006]='h00000000;
    rd_cycle[22007] = 1'b1;  wr_cycle[22007] = 1'b0;  addr_rom[22007]='h000017dc;  wr_data_rom[22007]='h00000000;
    rd_cycle[22008] = 1'b1;  wr_cycle[22008] = 1'b0;  addr_rom[22008]='h000017e0;  wr_data_rom[22008]='h00000000;
    rd_cycle[22009] = 1'b1;  wr_cycle[22009] = 1'b0;  addr_rom[22009]='h000017e4;  wr_data_rom[22009]='h00000000;
    rd_cycle[22010] = 1'b1;  wr_cycle[22010] = 1'b0;  addr_rom[22010]='h000017e8;  wr_data_rom[22010]='h00000000;
    rd_cycle[22011] = 1'b1;  wr_cycle[22011] = 1'b0;  addr_rom[22011]='h000017ec;  wr_data_rom[22011]='h00000000;
    rd_cycle[22012] = 1'b1;  wr_cycle[22012] = 1'b0;  addr_rom[22012]='h000017f0;  wr_data_rom[22012]='h00000000;
    rd_cycle[22013] = 1'b1;  wr_cycle[22013] = 1'b0;  addr_rom[22013]='h000017f4;  wr_data_rom[22013]='h00000000;
    rd_cycle[22014] = 1'b1;  wr_cycle[22014] = 1'b0;  addr_rom[22014]='h000017f8;  wr_data_rom[22014]='h00000000;
    rd_cycle[22015] = 1'b1;  wr_cycle[22015] = 1'b0;  addr_rom[22015]='h000017fc;  wr_data_rom[22015]='h00000000;
    rd_cycle[22016] = 1'b1;  wr_cycle[22016] = 1'b0;  addr_rom[22016]='h00001800;  wr_data_rom[22016]='h00000000;
    rd_cycle[22017] = 1'b1;  wr_cycle[22017] = 1'b0;  addr_rom[22017]='h00001804;  wr_data_rom[22017]='h00000000;
    rd_cycle[22018] = 1'b1;  wr_cycle[22018] = 1'b0;  addr_rom[22018]='h00001808;  wr_data_rom[22018]='h00000000;
    rd_cycle[22019] = 1'b1;  wr_cycle[22019] = 1'b0;  addr_rom[22019]='h0000180c;  wr_data_rom[22019]='h00000000;
    rd_cycle[22020] = 1'b1;  wr_cycle[22020] = 1'b0;  addr_rom[22020]='h00001810;  wr_data_rom[22020]='h00000000;
    rd_cycle[22021] = 1'b1;  wr_cycle[22021] = 1'b0;  addr_rom[22021]='h00001814;  wr_data_rom[22021]='h00000000;
    rd_cycle[22022] = 1'b1;  wr_cycle[22022] = 1'b0;  addr_rom[22022]='h00001818;  wr_data_rom[22022]='h00000000;
    rd_cycle[22023] = 1'b1;  wr_cycle[22023] = 1'b0;  addr_rom[22023]='h0000181c;  wr_data_rom[22023]='h00000000;
    rd_cycle[22024] = 1'b1;  wr_cycle[22024] = 1'b0;  addr_rom[22024]='h00001820;  wr_data_rom[22024]='h00000000;
    rd_cycle[22025] = 1'b1;  wr_cycle[22025] = 1'b0;  addr_rom[22025]='h00001824;  wr_data_rom[22025]='h00000000;
    rd_cycle[22026] = 1'b1;  wr_cycle[22026] = 1'b0;  addr_rom[22026]='h00001828;  wr_data_rom[22026]='h00000000;
    rd_cycle[22027] = 1'b1;  wr_cycle[22027] = 1'b0;  addr_rom[22027]='h0000182c;  wr_data_rom[22027]='h00000000;
    rd_cycle[22028] = 1'b1;  wr_cycle[22028] = 1'b0;  addr_rom[22028]='h00001830;  wr_data_rom[22028]='h00000000;
    rd_cycle[22029] = 1'b1;  wr_cycle[22029] = 1'b0;  addr_rom[22029]='h00001834;  wr_data_rom[22029]='h00000000;
    rd_cycle[22030] = 1'b1;  wr_cycle[22030] = 1'b0;  addr_rom[22030]='h00001838;  wr_data_rom[22030]='h00000000;
    rd_cycle[22031] = 1'b1;  wr_cycle[22031] = 1'b0;  addr_rom[22031]='h0000183c;  wr_data_rom[22031]='h00000000;
    rd_cycle[22032] = 1'b1;  wr_cycle[22032] = 1'b0;  addr_rom[22032]='h00001840;  wr_data_rom[22032]='h00000000;
    rd_cycle[22033] = 1'b1;  wr_cycle[22033] = 1'b0;  addr_rom[22033]='h00001844;  wr_data_rom[22033]='h00000000;
    rd_cycle[22034] = 1'b1;  wr_cycle[22034] = 1'b0;  addr_rom[22034]='h00001848;  wr_data_rom[22034]='h00000000;
    rd_cycle[22035] = 1'b1;  wr_cycle[22035] = 1'b0;  addr_rom[22035]='h0000184c;  wr_data_rom[22035]='h00000000;
    rd_cycle[22036] = 1'b1;  wr_cycle[22036] = 1'b0;  addr_rom[22036]='h00001850;  wr_data_rom[22036]='h00000000;
    rd_cycle[22037] = 1'b1;  wr_cycle[22037] = 1'b0;  addr_rom[22037]='h00001854;  wr_data_rom[22037]='h00000000;
    rd_cycle[22038] = 1'b1;  wr_cycle[22038] = 1'b0;  addr_rom[22038]='h00001858;  wr_data_rom[22038]='h00000000;
    rd_cycle[22039] = 1'b1;  wr_cycle[22039] = 1'b0;  addr_rom[22039]='h0000185c;  wr_data_rom[22039]='h00000000;
    rd_cycle[22040] = 1'b1;  wr_cycle[22040] = 1'b0;  addr_rom[22040]='h00001860;  wr_data_rom[22040]='h00000000;
    rd_cycle[22041] = 1'b1;  wr_cycle[22041] = 1'b0;  addr_rom[22041]='h00001864;  wr_data_rom[22041]='h00000000;
    rd_cycle[22042] = 1'b1;  wr_cycle[22042] = 1'b0;  addr_rom[22042]='h00001868;  wr_data_rom[22042]='h00000000;
    rd_cycle[22043] = 1'b1;  wr_cycle[22043] = 1'b0;  addr_rom[22043]='h0000186c;  wr_data_rom[22043]='h00000000;
    rd_cycle[22044] = 1'b1;  wr_cycle[22044] = 1'b0;  addr_rom[22044]='h00001870;  wr_data_rom[22044]='h00000000;
    rd_cycle[22045] = 1'b1;  wr_cycle[22045] = 1'b0;  addr_rom[22045]='h00001874;  wr_data_rom[22045]='h00000000;
    rd_cycle[22046] = 1'b1;  wr_cycle[22046] = 1'b0;  addr_rom[22046]='h00001878;  wr_data_rom[22046]='h00000000;
    rd_cycle[22047] = 1'b1;  wr_cycle[22047] = 1'b0;  addr_rom[22047]='h0000187c;  wr_data_rom[22047]='h00000000;
    rd_cycle[22048] = 1'b1;  wr_cycle[22048] = 1'b0;  addr_rom[22048]='h00001880;  wr_data_rom[22048]='h00000000;
    rd_cycle[22049] = 1'b1;  wr_cycle[22049] = 1'b0;  addr_rom[22049]='h00001884;  wr_data_rom[22049]='h00000000;
    rd_cycle[22050] = 1'b1;  wr_cycle[22050] = 1'b0;  addr_rom[22050]='h00001888;  wr_data_rom[22050]='h00000000;
    rd_cycle[22051] = 1'b1;  wr_cycle[22051] = 1'b0;  addr_rom[22051]='h0000188c;  wr_data_rom[22051]='h00000000;
    rd_cycle[22052] = 1'b1;  wr_cycle[22052] = 1'b0;  addr_rom[22052]='h00001890;  wr_data_rom[22052]='h00000000;
    rd_cycle[22053] = 1'b1;  wr_cycle[22053] = 1'b0;  addr_rom[22053]='h00001894;  wr_data_rom[22053]='h00000000;
    rd_cycle[22054] = 1'b1;  wr_cycle[22054] = 1'b0;  addr_rom[22054]='h00001898;  wr_data_rom[22054]='h00000000;
    rd_cycle[22055] = 1'b1;  wr_cycle[22055] = 1'b0;  addr_rom[22055]='h0000189c;  wr_data_rom[22055]='h00000000;
    rd_cycle[22056] = 1'b1;  wr_cycle[22056] = 1'b0;  addr_rom[22056]='h000018a0;  wr_data_rom[22056]='h00000000;
    rd_cycle[22057] = 1'b1;  wr_cycle[22057] = 1'b0;  addr_rom[22057]='h000018a4;  wr_data_rom[22057]='h00000000;
    rd_cycle[22058] = 1'b1;  wr_cycle[22058] = 1'b0;  addr_rom[22058]='h000018a8;  wr_data_rom[22058]='h00000000;
    rd_cycle[22059] = 1'b1;  wr_cycle[22059] = 1'b0;  addr_rom[22059]='h000018ac;  wr_data_rom[22059]='h00000000;
    rd_cycle[22060] = 1'b1;  wr_cycle[22060] = 1'b0;  addr_rom[22060]='h000018b0;  wr_data_rom[22060]='h00000000;
    rd_cycle[22061] = 1'b1;  wr_cycle[22061] = 1'b0;  addr_rom[22061]='h000018b4;  wr_data_rom[22061]='h00000000;
    rd_cycle[22062] = 1'b1;  wr_cycle[22062] = 1'b0;  addr_rom[22062]='h000018b8;  wr_data_rom[22062]='h00000000;
    rd_cycle[22063] = 1'b1;  wr_cycle[22063] = 1'b0;  addr_rom[22063]='h000018bc;  wr_data_rom[22063]='h00000000;
    rd_cycle[22064] = 1'b1;  wr_cycle[22064] = 1'b0;  addr_rom[22064]='h000018c0;  wr_data_rom[22064]='h00000000;
    rd_cycle[22065] = 1'b1;  wr_cycle[22065] = 1'b0;  addr_rom[22065]='h000018c4;  wr_data_rom[22065]='h00000000;
    rd_cycle[22066] = 1'b1;  wr_cycle[22066] = 1'b0;  addr_rom[22066]='h000018c8;  wr_data_rom[22066]='h00000000;
    rd_cycle[22067] = 1'b1;  wr_cycle[22067] = 1'b0;  addr_rom[22067]='h000018cc;  wr_data_rom[22067]='h00000000;
    rd_cycle[22068] = 1'b1;  wr_cycle[22068] = 1'b0;  addr_rom[22068]='h000018d0;  wr_data_rom[22068]='h00000000;
    rd_cycle[22069] = 1'b1;  wr_cycle[22069] = 1'b0;  addr_rom[22069]='h000018d4;  wr_data_rom[22069]='h00000000;
    rd_cycle[22070] = 1'b1;  wr_cycle[22070] = 1'b0;  addr_rom[22070]='h000018d8;  wr_data_rom[22070]='h00000000;
    rd_cycle[22071] = 1'b1;  wr_cycle[22071] = 1'b0;  addr_rom[22071]='h000018dc;  wr_data_rom[22071]='h00000000;
    rd_cycle[22072] = 1'b1;  wr_cycle[22072] = 1'b0;  addr_rom[22072]='h000018e0;  wr_data_rom[22072]='h00000000;
    rd_cycle[22073] = 1'b1;  wr_cycle[22073] = 1'b0;  addr_rom[22073]='h000018e4;  wr_data_rom[22073]='h00000000;
    rd_cycle[22074] = 1'b1;  wr_cycle[22074] = 1'b0;  addr_rom[22074]='h000018e8;  wr_data_rom[22074]='h00000000;
    rd_cycle[22075] = 1'b1;  wr_cycle[22075] = 1'b0;  addr_rom[22075]='h000018ec;  wr_data_rom[22075]='h00000000;
    rd_cycle[22076] = 1'b1;  wr_cycle[22076] = 1'b0;  addr_rom[22076]='h000018f0;  wr_data_rom[22076]='h00000000;
    rd_cycle[22077] = 1'b1;  wr_cycle[22077] = 1'b0;  addr_rom[22077]='h000018f4;  wr_data_rom[22077]='h00000000;
    rd_cycle[22078] = 1'b1;  wr_cycle[22078] = 1'b0;  addr_rom[22078]='h000018f8;  wr_data_rom[22078]='h00000000;
    rd_cycle[22079] = 1'b1;  wr_cycle[22079] = 1'b0;  addr_rom[22079]='h000018fc;  wr_data_rom[22079]='h00000000;
    rd_cycle[22080] = 1'b1;  wr_cycle[22080] = 1'b0;  addr_rom[22080]='h00001900;  wr_data_rom[22080]='h00000000;
    rd_cycle[22081] = 1'b1;  wr_cycle[22081] = 1'b0;  addr_rom[22081]='h00001904;  wr_data_rom[22081]='h00000000;
    rd_cycle[22082] = 1'b1;  wr_cycle[22082] = 1'b0;  addr_rom[22082]='h00001908;  wr_data_rom[22082]='h00000000;
    rd_cycle[22083] = 1'b1;  wr_cycle[22083] = 1'b0;  addr_rom[22083]='h0000190c;  wr_data_rom[22083]='h00000000;
    rd_cycle[22084] = 1'b1;  wr_cycle[22084] = 1'b0;  addr_rom[22084]='h00001910;  wr_data_rom[22084]='h00000000;
    rd_cycle[22085] = 1'b1;  wr_cycle[22085] = 1'b0;  addr_rom[22085]='h00001914;  wr_data_rom[22085]='h00000000;
    rd_cycle[22086] = 1'b1;  wr_cycle[22086] = 1'b0;  addr_rom[22086]='h00001918;  wr_data_rom[22086]='h00000000;
    rd_cycle[22087] = 1'b1;  wr_cycle[22087] = 1'b0;  addr_rom[22087]='h0000191c;  wr_data_rom[22087]='h00000000;
    rd_cycle[22088] = 1'b1;  wr_cycle[22088] = 1'b0;  addr_rom[22088]='h00001920;  wr_data_rom[22088]='h00000000;
    rd_cycle[22089] = 1'b1;  wr_cycle[22089] = 1'b0;  addr_rom[22089]='h00001924;  wr_data_rom[22089]='h00000000;
    rd_cycle[22090] = 1'b1;  wr_cycle[22090] = 1'b0;  addr_rom[22090]='h00001928;  wr_data_rom[22090]='h00000000;
    rd_cycle[22091] = 1'b1;  wr_cycle[22091] = 1'b0;  addr_rom[22091]='h0000192c;  wr_data_rom[22091]='h00000000;
    rd_cycle[22092] = 1'b1;  wr_cycle[22092] = 1'b0;  addr_rom[22092]='h00001930;  wr_data_rom[22092]='h00000000;
    rd_cycle[22093] = 1'b1;  wr_cycle[22093] = 1'b0;  addr_rom[22093]='h00001934;  wr_data_rom[22093]='h00000000;
    rd_cycle[22094] = 1'b1;  wr_cycle[22094] = 1'b0;  addr_rom[22094]='h00001938;  wr_data_rom[22094]='h00000000;
    rd_cycle[22095] = 1'b1;  wr_cycle[22095] = 1'b0;  addr_rom[22095]='h0000193c;  wr_data_rom[22095]='h00000000;
    rd_cycle[22096] = 1'b1;  wr_cycle[22096] = 1'b0;  addr_rom[22096]='h00001940;  wr_data_rom[22096]='h00000000;
    rd_cycle[22097] = 1'b1;  wr_cycle[22097] = 1'b0;  addr_rom[22097]='h00001944;  wr_data_rom[22097]='h00000000;
    rd_cycle[22098] = 1'b1;  wr_cycle[22098] = 1'b0;  addr_rom[22098]='h00001948;  wr_data_rom[22098]='h00000000;
    rd_cycle[22099] = 1'b1;  wr_cycle[22099] = 1'b0;  addr_rom[22099]='h0000194c;  wr_data_rom[22099]='h00000000;
    rd_cycle[22100] = 1'b1;  wr_cycle[22100] = 1'b0;  addr_rom[22100]='h00001950;  wr_data_rom[22100]='h00000000;
    rd_cycle[22101] = 1'b1;  wr_cycle[22101] = 1'b0;  addr_rom[22101]='h00001954;  wr_data_rom[22101]='h00000000;
    rd_cycle[22102] = 1'b1;  wr_cycle[22102] = 1'b0;  addr_rom[22102]='h00001958;  wr_data_rom[22102]='h00000000;
    rd_cycle[22103] = 1'b1;  wr_cycle[22103] = 1'b0;  addr_rom[22103]='h0000195c;  wr_data_rom[22103]='h00000000;
    rd_cycle[22104] = 1'b1;  wr_cycle[22104] = 1'b0;  addr_rom[22104]='h00001960;  wr_data_rom[22104]='h00000000;
    rd_cycle[22105] = 1'b1;  wr_cycle[22105] = 1'b0;  addr_rom[22105]='h00001964;  wr_data_rom[22105]='h00000000;
    rd_cycle[22106] = 1'b1;  wr_cycle[22106] = 1'b0;  addr_rom[22106]='h00001968;  wr_data_rom[22106]='h00000000;
    rd_cycle[22107] = 1'b1;  wr_cycle[22107] = 1'b0;  addr_rom[22107]='h0000196c;  wr_data_rom[22107]='h00000000;
    rd_cycle[22108] = 1'b1;  wr_cycle[22108] = 1'b0;  addr_rom[22108]='h00001970;  wr_data_rom[22108]='h00000000;
    rd_cycle[22109] = 1'b1;  wr_cycle[22109] = 1'b0;  addr_rom[22109]='h00001974;  wr_data_rom[22109]='h00000000;
    rd_cycle[22110] = 1'b1;  wr_cycle[22110] = 1'b0;  addr_rom[22110]='h00001978;  wr_data_rom[22110]='h00000000;
    rd_cycle[22111] = 1'b1;  wr_cycle[22111] = 1'b0;  addr_rom[22111]='h0000197c;  wr_data_rom[22111]='h00000000;
    rd_cycle[22112] = 1'b1;  wr_cycle[22112] = 1'b0;  addr_rom[22112]='h00001980;  wr_data_rom[22112]='h00000000;
    rd_cycle[22113] = 1'b1;  wr_cycle[22113] = 1'b0;  addr_rom[22113]='h00001984;  wr_data_rom[22113]='h00000000;
    rd_cycle[22114] = 1'b1;  wr_cycle[22114] = 1'b0;  addr_rom[22114]='h00001988;  wr_data_rom[22114]='h00000000;
    rd_cycle[22115] = 1'b1;  wr_cycle[22115] = 1'b0;  addr_rom[22115]='h0000198c;  wr_data_rom[22115]='h00000000;
    rd_cycle[22116] = 1'b1;  wr_cycle[22116] = 1'b0;  addr_rom[22116]='h00001990;  wr_data_rom[22116]='h00000000;
    rd_cycle[22117] = 1'b1;  wr_cycle[22117] = 1'b0;  addr_rom[22117]='h00001994;  wr_data_rom[22117]='h00000000;
    rd_cycle[22118] = 1'b1;  wr_cycle[22118] = 1'b0;  addr_rom[22118]='h00001998;  wr_data_rom[22118]='h00000000;
    rd_cycle[22119] = 1'b1;  wr_cycle[22119] = 1'b0;  addr_rom[22119]='h0000199c;  wr_data_rom[22119]='h00000000;
    rd_cycle[22120] = 1'b1;  wr_cycle[22120] = 1'b0;  addr_rom[22120]='h000019a0;  wr_data_rom[22120]='h00000000;
    rd_cycle[22121] = 1'b1;  wr_cycle[22121] = 1'b0;  addr_rom[22121]='h000019a4;  wr_data_rom[22121]='h00000000;
    rd_cycle[22122] = 1'b1;  wr_cycle[22122] = 1'b0;  addr_rom[22122]='h000019a8;  wr_data_rom[22122]='h00000000;
    rd_cycle[22123] = 1'b1;  wr_cycle[22123] = 1'b0;  addr_rom[22123]='h000019ac;  wr_data_rom[22123]='h00000000;
    rd_cycle[22124] = 1'b1;  wr_cycle[22124] = 1'b0;  addr_rom[22124]='h000019b0;  wr_data_rom[22124]='h00000000;
    rd_cycle[22125] = 1'b1;  wr_cycle[22125] = 1'b0;  addr_rom[22125]='h000019b4;  wr_data_rom[22125]='h00000000;
    rd_cycle[22126] = 1'b1;  wr_cycle[22126] = 1'b0;  addr_rom[22126]='h000019b8;  wr_data_rom[22126]='h00000000;
    rd_cycle[22127] = 1'b1;  wr_cycle[22127] = 1'b0;  addr_rom[22127]='h000019bc;  wr_data_rom[22127]='h00000000;
    rd_cycle[22128] = 1'b1;  wr_cycle[22128] = 1'b0;  addr_rom[22128]='h000019c0;  wr_data_rom[22128]='h00000000;
    rd_cycle[22129] = 1'b1;  wr_cycle[22129] = 1'b0;  addr_rom[22129]='h000019c4;  wr_data_rom[22129]='h00000000;
    rd_cycle[22130] = 1'b1;  wr_cycle[22130] = 1'b0;  addr_rom[22130]='h000019c8;  wr_data_rom[22130]='h00000000;
    rd_cycle[22131] = 1'b1;  wr_cycle[22131] = 1'b0;  addr_rom[22131]='h000019cc;  wr_data_rom[22131]='h00000000;
    rd_cycle[22132] = 1'b1;  wr_cycle[22132] = 1'b0;  addr_rom[22132]='h000019d0;  wr_data_rom[22132]='h00000000;
    rd_cycle[22133] = 1'b1;  wr_cycle[22133] = 1'b0;  addr_rom[22133]='h000019d4;  wr_data_rom[22133]='h00000000;
    rd_cycle[22134] = 1'b1;  wr_cycle[22134] = 1'b0;  addr_rom[22134]='h000019d8;  wr_data_rom[22134]='h00000000;
    rd_cycle[22135] = 1'b1;  wr_cycle[22135] = 1'b0;  addr_rom[22135]='h000019dc;  wr_data_rom[22135]='h00000000;
    rd_cycle[22136] = 1'b1;  wr_cycle[22136] = 1'b0;  addr_rom[22136]='h000019e0;  wr_data_rom[22136]='h00000000;
    rd_cycle[22137] = 1'b1;  wr_cycle[22137] = 1'b0;  addr_rom[22137]='h000019e4;  wr_data_rom[22137]='h00000000;
    rd_cycle[22138] = 1'b1;  wr_cycle[22138] = 1'b0;  addr_rom[22138]='h000019e8;  wr_data_rom[22138]='h00000000;
    rd_cycle[22139] = 1'b1;  wr_cycle[22139] = 1'b0;  addr_rom[22139]='h000019ec;  wr_data_rom[22139]='h00000000;
    rd_cycle[22140] = 1'b1;  wr_cycle[22140] = 1'b0;  addr_rom[22140]='h000019f0;  wr_data_rom[22140]='h00000000;
    rd_cycle[22141] = 1'b1;  wr_cycle[22141] = 1'b0;  addr_rom[22141]='h000019f4;  wr_data_rom[22141]='h00000000;
    rd_cycle[22142] = 1'b1;  wr_cycle[22142] = 1'b0;  addr_rom[22142]='h000019f8;  wr_data_rom[22142]='h00000000;
    rd_cycle[22143] = 1'b1;  wr_cycle[22143] = 1'b0;  addr_rom[22143]='h000019fc;  wr_data_rom[22143]='h00000000;
    rd_cycle[22144] = 1'b1;  wr_cycle[22144] = 1'b0;  addr_rom[22144]='h00001a00;  wr_data_rom[22144]='h00000000;
    rd_cycle[22145] = 1'b1;  wr_cycle[22145] = 1'b0;  addr_rom[22145]='h00001a04;  wr_data_rom[22145]='h00000000;
    rd_cycle[22146] = 1'b1;  wr_cycle[22146] = 1'b0;  addr_rom[22146]='h00001a08;  wr_data_rom[22146]='h00000000;
    rd_cycle[22147] = 1'b1;  wr_cycle[22147] = 1'b0;  addr_rom[22147]='h00001a0c;  wr_data_rom[22147]='h00000000;
    rd_cycle[22148] = 1'b1;  wr_cycle[22148] = 1'b0;  addr_rom[22148]='h00001a10;  wr_data_rom[22148]='h00000000;
    rd_cycle[22149] = 1'b1;  wr_cycle[22149] = 1'b0;  addr_rom[22149]='h00001a14;  wr_data_rom[22149]='h00000000;
    rd_cycle[22150] = 1'b1;  wr_cycle[22150] = 1'b0;  addr_rom[22150]='h00001a18;  wr_data_rom[22150]='h00000000;
    rd_cycle[22151] = 1'b1;  wr_cycle[22151] = 1'b0;  addr_rom[22151]='h00001a1c;  wr_data_rom[22151]='h00000000;
    rd_cycle[22152] = 1'b1;  wr_cycle[22152] = 1'b0;  addr_rom[22152]='h00001a20;  wr_data_rom[22152]='h00000000;
    rd_cycle[22153] = 1'b1;  wr_cycle[22153] = 1'b0;  addr_rom[22153]='h00001a24;  wr_data_rom[22153]='h00000000;
    rd_cycle[22154] = 1'b1;  wr_cycle[22154] = 1'b0;  addr_rom[22154]='h00001a28;  wr_data_rom[22154]='h00000000;
    rd_cycle[22155] = 1'b1;  wr_cycle[22155] = 1'b0;  addr_rom[22155]='h00001a2c;  wr_data_rom[22155]='h00000000;
    rd_cycle[22156] = 1'b1;  wr_cycle[22156] = 1'b0;  addr_rom[22156]='h00001a30;  wr_data_rom[22156]='h00000000;
    rd_cycle[22157] = 1'b1;  wr_cycle[22157] = 1'b0;  addr_rom[22157]='h00001a34;  wr_data_rom[22157]='h00000000;
    rd_cycle[22158] = 1'b1;  wr_cycle[22158] = 1'b0;  addr_rom[22158]='h00001a38;  wr_data_rom[22158]='h00000000;
    rd_cycle[22159] = 1'b1;  wr_cycle[22159] = 1'b0;  addr_rom[22159]='h00001a3c;  wr_data_rom[22159]='h00000000;
    rd_cycle[22160] = 1'b1;  wr_cycle[22160] = 1'b0;  addr_rom[22160]='h00001a40;  wr_data_rom[22160]='h00000000;
    rd_cycle[22161] = 1'b1;  wr_cycle[22161] = 1'b0;  addr_rom[22161]='h00001a44;  wr_data_rom[22161]='h00000000;
    rd_cycle[22162] = 1'b1;  wr_cycle[22162] = 1'b0;  addr_rom[22162]='h00001a48;  wr_data_rom[22162]='h00000000;
    rd_cycle[22163] = 1'b1;  wr_cycle[22163] = 1'b0;  addr_rom[22163]='h00001a4c;  wr_data_rom[22163]='h00000000;
    rd_cycle[22164] = 1'b1;  wr_cycle[22164] = 1'b0;  addr_rom[22164]='h00001a50;  wr_data_rom[22164]='h00000000;
    rd_cycle[22165] = 1'b1;  wr_cycle[22165] = 1'b0;  addr_rom[22165]='h00001a54;  wr_data_rom[22165]='h00000000;
    rd_cycle[22166] = 1'b1;  wr_cycle[22166] = 1'b0;  addr_rom[22166]='h00001a58;  wr_data_rom[22166]='h00000000;
    rd_cycle[22167] = 1'b1;  wr_cycle[22167] = 1'b0;  addr_rom[22167]='h00001a5c;  wr_data_rom[22167]='h00000000;
    rd_cycle[22168] = 1'b1;  wr_cycle[22168] = 1'b0;  addr_rom[22168]='h00001a60;  wr_data_rom[22168]='h00000000;
    rd_cycle[22169] = 1'b1;  wr_cycle[22169] = 1'b0;  addr_rom[22169]='h00001a64;  wr_data_rom[22169]='h00000000;
    rd_cycle[22170] = 1'b1;  wr_cycle[22170] = 1'b0;  addr_rom[22170]='h00001a68;  wr_data_rom[22170]='h00000000;
    rd_cycle[22171] = 1'b1;  wr_cycle[22171] = 1'b0;  addr_rom[22171]='h00001a6c;  wr_data_rom[22171]='h00000000;
    rd_cycle[22172] = 1'b1;  wr_cycle[22172] = 1'b0;  addr_rom[22172]='h00001a70;  wr_data_rom[22172]='h00000000;
    rd_cycle[22173] = 1'b1;  wr_cycle[22173] = 1'b0;  addr_rom[22173]='h00001a74;  wr_data_rom[22173]='h00000000;
    rd_cycle[22174] = 1'b1;  wr_cycle[22174] = 1'b0;  addr_rom[22174]='h00001a78;  wr_data_rom[22174]='h00000000;
    rd_cycle[22175] = 1'b1;  wr_cycle[22175] = 1'b0;  addr_rom[22175]='h00001a7c;  wr_data_rom[22175]='h00000000;
    rd_cycle[22176] = 1'b1;  wr_cycle[22176] = 1'b0;  addr_rom[22176]='h00001a80;  wr_data_rom[22176]='h00000000;
    rd_cycle[22177] = 1'b1;  wr_cycle[22177] = 1'b0;  addr_rom[22177]='h00001a84;  wr_data_rom[22177]='h00000000;
    rd_cycle[22178] = 1'b1;  wr_cycle[22178] = 1'b0;  addr_rom[22178]='h00001a88;  wr_data_rom[22178]='h00000000;
    rd_cycle[22179] = 1'b1;  wr_cycle[22179] = 1'b0;  addr_rom[22179]='h00001a8c;  wr_data_rom[22179]='h00000000;
    rd_cycle[22180] = 1'b1;  wr_cycle[22180] = 1'b0;  addr_rom[22180]='h00001a90;  wr_data_rom[22180]='h00000000;
    rd_cycle[22181] = 1'b1;  wr_cycle[22181] = 1'b0;  addr_rom[22181]='h00001a94;  wr_data_rom[22181]='h00000000;
    rd_cycle[22182] = 1'b1;  wr_cycle[22182] = 1'b0;  addr_rom[22182]='h00001a98;  wr_data_rom[22182]='h00000000;
    rd_cycle[22183] = 1'b1;  wr_cycle[22183] = 1'b0;  addr_rom[22183]='h00001a9c;  wr_data_rom[22183]='h00000000;
    rd_cycle[22184] = 1'b1;  wr_cycle[22184] = 1'b0;  addr_rom[22184]='h00001aa0;  wr_data_rom[22184]='h00000000;
    rd_cycle[22185] = 1'b1;  wr_cycle[22185] = 1'b0;  addr_rom[22185]='h00001aa4;  wr_data_rom[22185]='h00000000;
    rd_cycle[22186] = 1'b1;  wr_cycle[22186] = 1'b0;  addr_rom[22186]='h00001aa8;  wr_data_rom[22186]='h00000000;
    rd_cycle[22187] = 1'b1;  wr_cycle[22187] = 1'b0;  addr_rom[22187]='h00001aac;  wr_data_rom[22187]='h00000000;
    rd_cycle[22188] = 1'b1;  wr_cycle[22188] = 1'b0;  addr_rom[22188]='h00001ab0;  wr_data_rom[22188]='h00000000;
    rd_cycle[22189] = 1'b1;  wr_cycle[22189] = 1'b0;  addr_rom[22189]='h00001ab4;  wr_data_rom[22189]='h00000000;
    rd_cycle[22190] = 1'b1;  wr_cycle[22190] = 1'b0;  addr_rom[22190]='h00001ab8;  wr_data_rom[22190]='h00000000;
    rd_cycle[22191] = 1'b1;  wr_cycle[22191] = 1'b0;  addr_rom[22191]='h00001abc;  wr_data_rom[22191]='h00000000;
    rd_cycle[22192] = 1'b1;  wr_cycle[22192] = 1'b0;  addr_rom[22192]='h00001ac0;  wr_data_rom[22192]='h00000000;
    rd_cycle[22193] = 1'b1;  wr_cycle[22193] = 1'b0;  addr_rom[22193]='h00001ac4;  wr_data_rom[22193]='h00000000;
    rd_cycle[22194] = 1'b1;  wr_cycle[22194] = 1'b0;  addr_rom[22194]='h00001ac8;  wr_data_rom[22194]='h00000000;
    rd_cycle[22195] = 1'b1;  wr_cycle[22195] = 1'b0;  addr_rom[22195]='h00001acc;  wr_data_rom[22195]='h00000000;
    rd_cycle[22196] = 1'b1;  wr_cycle[22196] = 1'b0;  addr_rom[22196]='h00001ad0;  wr_data_rom[22196]='h00000000;
    rd_cycle[22197] = 1'b1;  wr_cycle[22197] = 1'b0;  addr_rom[22197]='h00001ad4;  wr_data_rom[22197]='h00000000;
    rd_cycle[22198] = 1'b1;  wr_cycle[22198] = 1'b0;  addr_rom[22198]='h00001ad8;  wr_data_rom[22198]='h00000000;
    rd_cycle[22199] = 1'b1;  wr_cycle[22199] = 1'b0;  addr_rom[22199]='h00001adc;  wr_data_rom[22199]='h00000000;
    rd_cycle[22200] = 1'b1;  wr_cycle[22200] = 1'b0;  addr_rom[22200]='h00001ae0;  wr_data_rom[22200]='h00000000;
    rd_cycle[22201] = 1'b1;  wr_cycle[22201] = 1'b0;  addr_rom[22201]='h00001ae4;  wr_data_rom[22201]='h00000000;
    rd_cycle[22202] = 1'b1;  wr_cycle[22202] = 1'b0;  addr_rom[22202]='h00001ae8;  wr_data_rom[22202]='h00000000;
    rd_cycle[22203] = 1'b1;  wr_cycle[22203] = 1'b0;  addr_rom[22203]='h00001aec;  wr_data_rom[22203]='h00000000;
    rd_cycle[22204] = 1'b1;  wr_cycle[22204] = 1'b0;  addr_rom[22204]='h00001af0;  wr_data_rom[22204]='h00000000;
    rd_cycle[22205] = 1'b1;  wr_cycle[22205] = 1'b0;  addr_rom[22205]='h00001af4;  wr_data_rom[22205]='h00000000;
    rd_cycle[22206] = 1'b1;  wr_cycle[22206] = 1'b0;  addr_rom[22206]='h00001af8;  wr_data_rom[22206]='h00000000;
    rd_cycle[22207] = 1'b1;  wr_cycle[22207] = 1'b0;  addr_rom[22207]='h00001afc;  wr_data_rom[22207]='h00000000;
    rd_cycle[22208] = 1'b1;  wr_cycle[22208] = 1'b0;  addr_rom[22208]='h00001b00;  wr_data_rom[22208]='h00000000;
    rd_cycle[22209] = 1'b1;  wr_cycle[22209] = 1'b0;  addr_rom[22209]='h00001b04;  wr_data_rom[22209]='h00000000;
    rd_cycle[22210] = 1'b1;  wr_cycle[22210] = 1'b0;  addr_rom[22210]='h00001b08;  wr_data_rom[22210]='h00000000;
    rd_cycle[22211] = 1'b1;  wr_cycle[22211] = 1'b0;  addr_rom[22211]='h00001b0c;  wr_data_rom[22211]='h00000000;
    rd_cycle[22212] = 1'b1;  wr_cycle[22212] = 1'b0;  addr_rom[22212]='h00001b10;  wr_data_rom[22212]='h00000000;
    rd_cycle[22213] = 1'b1;  wr_cycle[22213] = 1'b0;  addr_rom[22213]='h00001b14;  wr_data_rom[22213]='h00000000;
    rd_cycle[22214] = 1'b1;  wr_cycle[22214] = 1'b0;  addr_rom[22214]='h00001b18;  wr_data_rom[22214]='h00000000;
    rd_cycle[22215] = 1'b1;  wr_cycle[22215] = 1'b0;  addr_rom[22215]='h00001b1c;  wr_data_rom[22215]='h00000000;
    rd_cycle[22216] = 1'b1;  wr_cycle[22216] = 1'b0;  addr_rom[22216]='h00001b20;  wr_data_rom[22216]='h00000000;
    rd_cycle[22217] = 1'b1;  wr_cycle[22217] = 1'b0;  addr_rom[22217]='h00001b24;  wr_data_rom[22217]='h00000000;
    rd_cycle[22218] = 1'b1;  wr_cycle[22218] = 1'b0;  addr_rom[22218]='h00001b28;  wr_data_rom[22218]='h00000000;
    rd_cycle[22219] = 1'b1;  wr_cycle[22219] = 1'b0;  addr_rom[22219]='h00001b2c;  wr_data_rom[22219]='h00000000;
    rd_cycle[22220] = 1'b1;  wr_cycle[22220] = 1'b0;  addr_rom[22220]='h00001b30;  wr_data_rom[22220]='h00000000;
    rd_cycle[22221] = 1'b1;  wr_cycle[22221] = 1'b0;  addr_rom[22221]='h00001b34;  wr_data_rom[22221]='h00000000;
    rd_cycle[22222] = 1'b1;  wr_cycle[22222] = 1'b0;  addr_rom[22222]='h00001b38;  wr_data_rom[22222]='h00000000;
    rd_cycle[22223] = 1'b1;  wr_cycle[22223] = 1'b0;  addr_rom[22223]='h00001b3c;  wr_data_rom[22223]='h00000000;
    rd_cycle[22224] = 1'b1;  wr_cycle[22224] = 1'b0;  addr_rom[22224]='h00001b40;  wr_data_rom[22224]='h00000000;
    rd_cycle[22225] = 1'b1;  wr_cycle[22225] = 1'b0;  addr_rom[22225]='h00001b44;  wr_data_rom[22225]='h00000000;
    rd_cycle[22226] = 1'b1;  wr_cycle[22226] = 1'b0;  addr_rom[22226]='h00001b48;  wr_data_rom[22226]='h00000000;
    rd_cycle[22227] = 1'b1;  wr_cycle[22227] = 1'b0;  addr_rom[22227]='h00001b4c;  wr_data_rom[22227]='h00000000;
    rd_cycle[22228] = 1'b1;  wr_cycle[22228] = 1'b0;  addr_rom[22228]='h00001b50;  wr_data_rom[22228]='h00000000;
    rd_cycle[22229] = 1'b1;  wr_cycle[22229] = 1'b0;  addr_rom[22229]='h00001b54;  wr_data_rom[22229]='h00000000;
    rd_cycle[22230] = 1'b1;  wr_cycle[22230] = 1'b0;  addr_rom[22230]='h00001b58;  wr_data_rom[22230]='h00000000;
    rd_cycle[22231] = 1'b1;  wr_cycle[22231] = 1'b0;  addr_rom[22231]='h00001b5c;  wr_data_rom[22231]='h00000000;
    rd_cycle[22232] = 1'b1;  wr_cycle[22232] = 1'b0;  addr_rom[22232]='h00001b60;  wr_data_rom[22232]='h00000000;
    rd_cycle[22233] = 1'b1;  wr_cycle[22233] = 1'b0;  addr_rom[22233]='h00001b64;  wr_data_rom[22233]='h00000000;
    rd_cycle[22234] = 1'b1;  wr_cycle[22234] = 1'b0;  addr_rom[22234]='h00001b68;  wr_data_rom[22234]='h00000000;
    rd_cycle[22235] = 1'b1;  wr_cycle[22235] = 1'b0;  addr_rom[22235]='h00001b6c;  wr_data_rom[22235]='h00000000;
    rd_cycle[22236] = 1'b1;  wr_cycle[22236] = 1'b0;  addr_rom[22236]='h00001b70;  wr_data_rom[22236]='h00000000;
    rd_cycle[22237] = 1'b1;  wr_cycle[22237] = 1'b0;  addr_rom[22237]='h00001b74;  wr_data_rom[22237]='h00000000;
    rd_cycle[22238] = 1'b1;  wr_cycle[22238] = 1'b0;  addr_rom[22238]='h00001b78;  wr_data_rom[22238]='h00000000;
    rd_cycle[22239] = 1'b1;  wr_cycle[22239] = 1'b0;  addr_rom[22239]='h00001b7c;  wr_data_rom[22239]='h00000000;
    rd_cycle[22240] = 1'b1;  wr_cycle[22240] = 1'b0;  addr_rom[22240]='h00001b80;  wr_data_rom[22240]='h00000000;
    rd_cycle[22241] = 1'b1;  wr_cycle[22241] = 1'b0;  addr_rom[22241]='h00001b84;  wr_data_rom[22241]='h00000000;
    rd_cycle[22242] = 1'b1;  wr_cycle[22242] = 1'b0;  addr_rom[22242]='h00001b88;  wr_data_rom[22242]='h00000000;
    rd_cycle[22243] = 1'b1;  wr_cycle[22243] = 1'b0;  addr_rom[22243]='h00001b8c;  wr_data_rom[22243]='h00000000;
    rd_cycle[22244] = 1'b1;  wr_cycle[22244] = 1'b0;  addr_rom[22244]='h00001b90;  wr_data_rom[22244]='h00000000;
    rd_cycle[22245] = 1'b1;  wr_cycle[22245] = 1'b0;  addr_rom[22245]='h00001b94;  wr_data_rom[22245]='h00000000;
    rd_cycle[22246] = 1'b1;  wr_cycle[22246] = 1'b0;  addr_rom[22246]='h00001b98;  wr_data_rom[22246]='h00000000;
    rd_cycle[22247] = 1'b1;  wr_cycle[22247] = 1'b0;  addr_rom[22247]='h00001b9c;  wr_data_rom[22247]='h00000000;
    rd_cycle[22248] = 1'b1;  wr_cycle[22248] = 1'b0;  addr_rom[22248]='h00001ba0;  wr_data_rom[22248]='h00000000;
    rd_cycle[22249] = 1'b1;  wr_cycle[22249] = 1'b0;  addr_rom[22249]='h00001ba4;  wr_data_rom[22249]='h00000000;
    rd_cycle[22250] = 1'b1;  wr_cycle[22250] = 1'b0;  addr_rom[22250]='h00001ba8;  wr_data_rom[22250]='h00000000;
    rd_cycle[22251] = 1'b1;  wr_cycle[22251] = 1'b0;  addr_rom[22251]='h00001bac;  wr_data_rom[22251]='h00000000;
    rd_cycle[22252] = 1'b1;  wr_cycle[22252] = 1'b0;  addr_rom[22252]='h00001bb0;  wr_data_rom[22252]='h00000000;
    rd_cycle[22253] = 1'b1;  wr_cycle[22253] = 1'b0;  addr_rom[22253]='h00001bb4;  wr_data_rom[22253]='h00000000;
    rd_cycle[22254] = 1'b1;  wr_cycle[22254] = 1'b0;  addr_rom[22254]='h00001bb8;  wr_data_rom[22254]='h00000000;
    rd_cycle[22255] = 1'b1;  wr_cycle[22255] = 1'b0;  addr_rom[22255]='h00001bbc;  wr_data_rom[22255]='h00000000;
    rd_cycle[22256] = 1'b1;  wr_cycle[22256] = 1'b0;  addr_rom[22256]='h00001bc0;  wr_data_rom[22256]='h00000000;
    rd_cycle[22257] = 1'b1;  wr_cycle[22257] = 1'b0;  addr_rom[22257]='h00001bc4;  wr_data_rom[22257]='h00000000;
    rd_cycle[22258] = 1'b1;  wr_cycle[22258] = 1'b0;  addr_rom[22258]='h00001bc8;  wr_data_rom[22258]='h00000000;
    rd_cycle[22259] = 1'b1;  wr_cycle[22259] = 1'b0;  addr_rom[22259]='h00001bcc;  wr_data_rom[22259]='h00000000;
    rd_cycle[22260] = 1'b1;  wr_cycle[22260] = 1'b0;  addr_rom[22260]='h00001bd0;  wr_data_rom[22260]='h00000000;
    rd_cycle[22261] = 1'b1;  wr_cycle[22261] = 1'b0;  addr_rom[22261]='h00001bd4;  wr_data_rom[22261]='h00000000;
    rd_cycle[22262] = 1'b1;  wr_cycle[22262] = 1'b0;  addr_rom[22262]='h00001bd8;  wr_data_rom[22262]='h00000000;
    rd_cycle[22263] = 1'b1;  wr_cycle[22263] = 1'b0;  addr_rom[22263]='h00001bdc;  wr_data_rom[22263]='h00000000;
    rd_cycle[22264] = 1'b1;  wr_cycle[22264] = 1'b0;  addr_rom[22264]='h00001be0;  wr_data_rom[22264]='h00000000;
    rd_cycle[22265] = 1'b1;  wr_cycle[22265] = 1'b0;  addr_rom[22265]='h00001be4;  wr_data_rom[22265]='h00000000;
    rd_cycle[22266] = 1'b1;  wr_cycle[22266] = 1'b0;  addr_rom[22266]='h00001be8;  wr_data_rom[22266]='h00000000;
    rd_cycle[22267] = 1'b1;  wr_cycle[22267] = 1'b0;  addr_rom[22267]='h00001bec;  wr_data_rom[22267]='h00000000;
    rd_cycle[22268] = 1'b1;  wr_cycle[22268] = 1'b0;  addr_rom[22268]='h00001bf0;  wr_data_rom[22268]='h00000000;
    rd_cycle[22269] = 1'b1;  wr_cycle[22269] = 1'b0;  addr_rom[22269]='h00001bf4;  wr_data_rom[22269]='h00000000;
    rd_cycle[22270] = 1'b1;  wr_cycle[22270] = 1'b0;  addr_rom[22270]='h00001bf8;  wr_data_rom[22270]='h00000000;
    rd_cycle[22271] = 1'b1;  wr_cycle[22271] = 1'b0;  addr_rom[22271]='h00001bfc;  wr_data_rom[22271]='h00000000;
    rd_cycle[22272] = 1'b1;  wr_cycle[22272] = 1'b0;  addr_rom[22272]='h00001c00;  wr_data_rom[22272]='h00000000;
    rd_cycle[22273] = 1'b1;  wr_cycle[22273] = 1'b0;  addr_rom[22273]='h00001c04;  wr_data_rom[22273]='h00000000;
    rd_cycle[22274] = 1'b1;  wr_cycle[22274] = 1'b0;  addr_rom[22274]='h00001c08;  wr_data_rom[22274]='h00000000;
    rd_cycle[22275] = 1'b1;  wr_cycle[22275] = 1'b0;  addr_rom[22275]='h00001c0c;  wr_data_rom[22275]='h00000000;
    rd_cycle[22276] = 1'b1;  wr_cycle[22276] = 1'b0;  addr_rom[22276]='h00001c10;  wr_data_rom[22276]='h00000000;
    rd_cycle[22277] = 1'b1;  wr_cycle[22277] = 1'b0;  addr_rom[22277]='h00001c14;  wr_data_rom[22277]='h00000000;
    rd_cycle[22278] = 1'b1;  wr_cycle[22278] = 1'b0;  addr_rom[22278]='h00001c18;  wr_data_rom[22278]='h00000000;
    rd_cycle[22279] = 1'b1;  wr_cycle[22279] = 1'b0;  addr_rom[22279]='h00001c1c;  wr_data_rom[22279]='h00000000;
    rd_cycle[22280] = 1'b1;  wr_cycle[22280] = 1'b0;  addr_rom[22280]='h00001c20;  wr_data_rom[22280]='h00000000;
    rd_cycle[22281] = 1'b1;  wr_cycle[22281] = 1'b0;  addr_rom[22281]='h00001c24;  wr_data_rom[22281]='h00000000;
    rd_cycle[22282] = 1'b1;  wr_cycle[22282] = 1'b0;  addr_rom[22282]='h00001c28;  wr_data_rom[22282]='h00000000;
    rd_cycle[22283] = 1'b1;  wr_cycle[22283] = 1'b0;  addr_rom[22283]='h00001c2c;  wr_data_rom[22283]='h00000000;
    rd_cycle[22284] = 1'b1;  wr_cycle[22284] = 1'b0;  addr_rom[22284]='h00001c30;  wr_data_rom[22284]='h00000000;
    rd_cycle[22285] = 1'b1;  wr_cycle[22285] = 1'b0;  addr_rom[22285]='h00001c34;  wr_data_rom[22285]='h00000000;
    rd_cycle[22286] = 1'b1;  wr_cycle[22286] = 1'b0;  addr_rom[22286]='h00001c38;  wr_data_rom[22286]='h00000000;
    rd_cycle[22287] = 1'b1;  wr_cycle[22287] = 1'b0;  addr_rom[22287]='h00001c3c;  wr_data_rom[22287]='h00000000;
    rd_cycle[22288] = 1'b1;  wr_cycle[22288] = 1'b0;  addr_rom[22288]='h00001c40;  wr_data_rom[22288]='h00000000;
    rd_cycle[22289] = 1'b1;  wr_cycle[22289] = 1'b0;  addr_rom[22289]='h00001c44;  wr_data_rom[22289]='h00000000;
    rd_cycle[22290] = 1'b1;  wr_cycle[22290] = 1'b0;  addr_rom[22290]='h00001c48;  wr_data_rom[22290]='h00000000;
    rd_cycle[22291] = 1'b1;  wr_cycle[22291] = 1'b0;  addr_rom[22291]='h00001c4c;  wr_data_rom[22291]='h00000000;
    rd_cycle[22292] = 1'b1;  wr_cycle[22292] = 1'b0;  addr_rom[22292]='h00001c50;  wr_data_rom[22292]='h00000000;
    rd_cycle[22293] = 1'b1;  wr_cycle[22293] = 1'b0;  addr_rom[22293]='h00001c54;  wr_data_rom[22293]='h00000000;
    rd_cycle[22294] = 1'b1;  wr_cycle[22294] = 1'b0;  addr_rom[22294]='h00001c58;  wr_data_rom[22294]='h00000000;
    rd_cycle[22295] = 1'b1;  wr_cycle[22295] = 1'b0;  addr_rom[22295]='h00001c5c;  wr_data_rom[22295]='h00000000;
    rd_cycle[22296] = 1'b1;  wr_cycle[22296] = 1'b0;  addr_rom[22296]='h00001c60;  wr_data_rom[22296]='h00000000;
    rd_cycle[22297] = 1'b1;  wr_cycle[22297] = 1'b0;  addr_rom[22297]='h00001c64;  wr_data_rom[22297]='h00000000;
    rd_cycle[22298] = 1'b1;  wr_cycle[22298] = 1'b0;  addr_rom[22298]='h00001c68;  wr_data_rom[22298]='h00000000;
    rd_cycle[22299] = 1'b1;  wr_cycle[22299] = 1'b0;  addr_rom[22299]='h00001c6c;  wr_data_rom[22299]='h00000000;
    rd_cycle[22300] = 1'b1;  wr_cycle[22300] = 1'b0;  addr_rom[22300]='h00001c70;  wr_data_rom[22300]='h00000000;
    rd_cycle[22301] = 1'b1;  wr_cycle[22301] = 1'b0;  addr_rom[22301]='h00001c74;  wr_data_rom[22301]='h00000000;
    rd_cycle[22302] = 1'b1;  wr_cycle[22302] = 1'b0;  addr_rom[22302]='h00001c78;  wr_data_rom[22302]='h00000000;
    rd_cycle[22303] = 1'b1;  wr_cycle[22303] = 1'b0;  addr_rom[22303]='h00001c7c;  wr_data_rom[22303]='h00000000;
    rd_cycle[22304] = 1'b1;  wr_cycle[22304] = 1'b0;  addr_rom[22304]='h00001c80;  wr_data_rom[22304]='h00000000;
    rd_cycle[22305] = 1'b1;  wr_cycle[22305] = 1'b0;  addr_rom[22305]='h00001c84;  wr_data_rom[22305]='h00000000;
    rd_cycle[22306] = 1'b1;  wr_cycle[22306] = 1'b0;  addr_rom[22306]='h00001c88;  wr_data_rom[22306]='h00000000;
    rd_cycle[22307] = 1'b1;  wr_cycle[22307] = 1'b0;  addr_rom[22307]='h00001c8c;  wr_data_rom[22307]='h00000000;
    rd_cycle[22308] = 1'b1;  wr_cycle[22308] = 1'b0;  addr_rom[22308]='h00001c90;  wr_data_rom[22308]='h00000000;
    rd_cycle[22309] = 1'b1;  wr_cycle[22309] = 1'b0;  addr_rom[22309]='h00001c94;  wr_data_rom[22309]='h00000000;
    rd_cycle[22310] = 1'b1;  wr_cycle[22310] = 1'b0;  addr_rom[22310]='h00001c98;  wr_data_rom[22310]='h00000000;
    rd_cycle[22311] = 1'b1;  wr_cycle[22311] = 1'b0;  addr_rom[22311]='h00001c9c;  wr_data_rom[22311]='h00000000;
    rd_cycle[22312] = 1'b1;  wr_cycle[22312] = 1'b0;  addr_rom[22312]='h00001ca0;  wr_data_rom[22312]='h00000000;
    rd_cycle[22313] = 1'b1;  wr_cycle[22313] = 1'b0;  addr_rom[22313]='h00001ca4;  wr_data_rom[22313]='h00000000;
    rd_cycle[22314] = 1'b1;  wr_cycle[22314] = 1'b0;  addr_rom[22314]='h00001ca8;  wr_data_rom[22314]='h00000000;
    rd_cycle[22315] = 1'b1;  wr_cycle[22315] = 1'b0;  addr_rom[22315]='h00001cac;  wr_data_rom[22315]='h00000000;
    rd_cycle[22316] = 1'b1;  wr_cycle[22316] = 1'b0;  addr_rom[22316]='h00001cb0;  wr_data_rom[22316]='h00000000;
    rd_cycle[22317] = 1'b1;  wr_cycle[22317] = 1'b0;  addr_rom[22317]='h00001cb4;  wr_data_rom[22317]='h00000000;
    rd_cycle[22318] = 1'b1;  wr_cycle[22318] = 1'b0;  addr_rom[22318]='h00001cb8;  wr_data_rom[22318]='h00000000;
    rd_cycle[22319] = 1'b1;  wr_cycle[22319] = 1'b0;  addr_rom[22319]='h00001cbc;  wr_data_rom[22319]='h00000000;
    rd_cycle[22320] = 1'b1;  wr_cycle[22320] = 1'b0;  addr_rom[22320]='h00001cc0;  wr_data_rom[22320]='h00000000;
    rd_cycle[22321] = 1'b1;  wr_cycle[22321] = 1'b0;  addr_rom[22321]='h00001cc4;  wr_data_rom[22321]='h00000000;
    rd_cycle[22322] = 1'b1;  wr_cycle[22322] = 1'b0;  addr_rom[22322]='h00001cc8;  wr_data_rom[22322]='h00000000;
    rd_cycle[22323] = 1'b1;  wr_cycle[22323] = 1'b0;  addr_rom[22323]='h00001ccc;  wr_data_rom[22323]='h00000000;
    rd_cycle[22324] = 1'b1;  wr_cycle[22324] = 1'b0;  addr_rom[22324]='h00001cd0;  wr_data_rom[22324]='h00000000;
    rd_cycle[22325] = 1'b1;  wr_cycle[22325] = 1'b0;  addr_rom[22325]='h00001cd4;  wr_data_rom[22325]='h00000000;
    rd_cycle[22326] = 1'b1;  wr_cycle[22326] = 1'b0;  addr_rom[22326]='h00001cd8;  wr_data_rom[22326]='h00000000;
    rd_cycle[22327] = 1'b1;  wr_cycle[22327] = 1'b0;  addr_rom[22327]='h00001cdc;  wr_data_rom[22327]='h00000000;
    rd_cycle[22328] = 1'b1;  wr_cycle[22328] = 1'b0;  addr_rom[22328]='h00001ce0;  wr_data_rom[22328]='h00000000;
    rd_cycle[22329] = 1'b1;  wr_cycle[22329] = 1'b0;  addr_rom[22329]='h00001ce4;  wr_data_rom[22329]='h00000000;
    rd_cycle[22330] = 1'b1;  wr_cycle[22330] = 1'b0;  addr_rom[22330]='h00001ce8;  wr_data_rom[22330]='h00000000;
    rd_cycle[22331] = 1'b1;  wr_cycle[22331] = 1'b0;  addr_rom[22331]='h00001cec;  wr_data_rom[22331]='h00000000;
    rd_cycle[22332] = 1'b1;  wr_cycle[22332] = 1'b0;  addr_rom[22332]='h00001cf0;  wr_data_rom[22332]='h00000000;
    rd_cycle[22333] = 1'b1;  wr_cycle[22333] = 1'b0;  addr_rom[22333]='h00001cf4;  wr_data_rom[22333]='h00000000;
    rd_cycle[22334] = 1'b1;  wr_cycle[22334] = 1'b0;  addr_rom[22334]='h00001cf8;  wr_data_rom[22334]='h00000000;
    rd_cycle[22335] = 1'b1;  wr_cycle[22335] = 1'b0;  addr_rom[22335]='h00001cfc;  wr_data_rom[22335]='h00000000;
    rd_cycle[22336] = 1'b1;  wr_cycle[22336] = 1'b0;  addr_rom[22336]='h00001d00;  wr_data_rom[22336]='h00000000;
    rd_cycle[22337] = 1'b1;  wr_cycle[22337] = 1'b0;  addr_rom[22337]='h00001d04;  wr_data_rom[22337]='h00000000;
    rd_cycle[22338] = 1'b1;  wr_cycle[22338] = 1'b0;  addr_rom[22338]='h00001d08;  wr_data_rom[22338]='h00000000;
    rd_cycle[22339] = 1'b1;  wr_cycle[22339] = 1'b0;  addr_rom[22339]='h00001d0c;  wr_data_rom[22339]='h00000000;
    rd_cycle[22340] = 1'b1;  wr_cycle[22340] = 1'b0;  addr_rom[22340]='h00001d10;  wr_data_rom[22340]='h00000000;
    rd_cycle[22341] = 1'b1;  wr_cycle[22341] = 1'b0;  addr_rom[22341]='h00001d14;  wr_data_rom[22341]='h00000000;
    rd_cycle[22342] = 1'b1;  wr_cycle[22342] = 1'b0;  addr_rom[22342]='h00001d18;  wr_data_rom[22342]='h00000000;
    rd_cycle[22343] = 1'b1;  wr_cycle[22343] = 1'b0;  addr_rom[22343]='h00001d1c;  wr_data_rom[22343]='h00000000;
    rd_cycle[22344] = 1'b1;  wr_cycle[22344] = 1'b0;  addr_rom[22344]='h00001d20;  wr_data_rom[22344]='h00000000;
    rd_cycle[22345] = 1'b1;  wr_cycle[22345] = 1'b0;  addr_rom[22345]='h00001d24;  wr_data_rom[22345]='h00000000;
    rd_cycle[22346] = 1'b1;  wr_cycle[22346] = 1'b0;  addr_rom[22346]='h00001d28;  wr_data_rom[22346]='h00000000;
    rd_cycle[22347] = 1'b1;  wr_cycle[22347] = 1'b0;  addr_rom[22347]='h00001d2c;  wr_data_rom[22347]='h00000000;
    rd_cycle[22348] = 1'b1;  wr_cycle[22348] = 1'b0;  addr_rom[22348]='h00001d30;  wr_data_rom[22348]='h00000000;
    rd_cycle[22349] = 1'b1;  wr_cycle[22349] = 1'b0;  addr_rom[22349]='h00001d34;  wr_data_rom[22349]='h00000000;
    rd_cycle[22350] = 1'b1;  wr_cycle[22350] = 1'b0;  addr_rom[22350]='h00001d38;  wr_data_rom[22350]='h00000000;
    rd_cycle[22351] = 1'b1;  wr_cycle[22351] = 1'b0;  addr_rom[22351]='h00001d3c;  wr_data_rom[22351]='h00000000;
    rd_cycle[22352] = 1'b1;  wr_cycle[22352] = 1'b0;  addr_rom[22352]='h00001d40;  wr_data_rom[22352]='h00000000;
    rd_cycle[22353] = 1'b1;  wr_cycle[22353] = 1'b0;  addr_rom[22353]='h00001d44;  wr_data_rom[22353]='h00000000;
    rd_cycle[22354] = 1'b1;  wr_cycle[22354] = 1'b0;  addr_rom[22354]='h00001d48;  wr_data_rom[22354]='h00000000;
    rd_cycle[22355] = 1'b1;  wr_cycle[22355] = 1'b0;  addr_rom[22355]='h00001d4c;  wr_data_rom[22355]='h00000000;
    rd_cycle[22356] = 1'b1;  wr_cycle[22356] = 1'b0;  addr_rom[22356]='h00001d50;  wr_data_rom[22356]='h00000000;
    rd_cycle[22357] = 1'b1;  wr_cycle[22357] = 1'b0;  addr_rom[22357]='h00001d54;  wr_data_rom[22357]='h00000000;
    rd_cycle[22358] = 1'b1;  wr_cycle[22358] = 1'b0;  addr_rom[22358]='h00001d58;  wr_data_rom[22358]='h00000000;
    rd_cycle[22359] = 1'b1;  wr_cycle[22359] = 1'b0;  addr_rom[22359]='h00001d5c;  wr_data_rom[22359]='h00000000;
    rd_cycle[22360] = 1'b1;  wr_cycle[22360] = 1'b0;  addr_rom[22360]='h00001d60;  wr_data_rom[22360]='h00000000;
    rd_cycle[22361] = 1'b1;  wr_cycle[22361] = 1'b0;  addr_rom[22361]='h00001d64;  wr_data_rom[22361]='h00000000;
    rd_cycle[22362] = 1'b1;  wr_cycle[22362] = 1'b0;  addr_rom[22362]='h00001d68;  wr_data_rom[22362]='h00000000;
    rd_cycle[22363] = 1'b1;  wr_cycle[22363] = 1'b0;  addr_rom[22363]='h00001d6c;  wr_data_rom[22363]='h00000000;
    rd_cycle[22364] = 1'b1;  wr_cycle[22364] = 1'b0;  addr_rom[22364]='h00001d70;  wr_data_rom[22364]='h00000000;
    rd_cycle[22365] = 1'b1;  wr_cycle[22365] = 1'b0;  addr_rom[22365]='h00001d74;  wr_data_rom[22365]='h00000000;
    rd_cycle[22366] = 1'b1;  wr_cycle[22366] = 1'b0;  addr_rom[22366]='h00001d78;  wr_data_rom[22366]='h00000000;
    rd_cycle[22367] = 1'b1;  wr_cycle[22367] = 1'b0;  addr_rom[22367]='h00001d7c;  wr_data_rom[22367]='h00000000;
    rd_cycle[22368] = 1'b1;  wr_cycle[22368] = 1'b0;  addr_rom[22368]='h00001d80;  wr_data_rom[22368]='h00000000;
    rd_cycle[22369] = 1'b1;  wr_cycle[22369] = 1'b0;  addr_rom[22369]='h00001d84;  wr_data_rom[22369]='h00000000;
    rd_cycle[22370] = 1'b1;  wr_cycle[22370] = 1'b0;  addr_rom[22370]='h00001d88;  wr_data_rom[22370]='h00000000;
    rd_cycle[22371] = 1'b1;  wr_cycle[22371] = 1'b0;  addr_rom[22371]='h00001d8c;  wr_data_rom[22371]='h00000000;
    rd_cycle[22372] = 1'b1;  wr_cycle[22372] = 1'b0;  addr_rom[22372]='h00001d90;  wr_data_rom[22372]='h00000000;
    rd_cycle[22373] = 1'b1;  wr_cycle[22373] = 1'b0;  addr_rom[22373]='h00001d94;  wr_data_rom[22373]='h00000000;
    rd_cycle[22374] = 1'b1;  wr_cycle[22374] = 1'b0;  addr_rom[22374]='h00001d98;  wr_data_rom[22374]='h00000000;
    rd_cycle[22375] = 1'b1;  wr_cycle[22375] = 1'b0;  addr_rom[22375]='h00001d9c;  wr_data_rom[22375]='h00000000;
    rd_cycle[22376] = 1'b1;  wr_cycle[22376] = 1'b0;  addr_rom[22376]='h00001da0;  wr_data_rom[22376]='h00000000;
    rd_cycle[22377] = 1'b1;  wr_cycle[22377] = 1'b0;  addr_rom[22377]='h00001da4;  wr_data_rom[22377]='h00000000;
    rd_cycle[22378] = 1'b1;  wr_cycle[22378] = 1'b0;  addr_rom[22378]='h00001da8;  wr_data_rom[22378]='h00000000;
    rd_cycle[22379] = 1'b1;  wr_cycle[22379] = 1'b0;  addr_rom[22379]='h00001dac;  wr_data_rom[22379]='h00000000;
    rd_cycle[22380] = 1'b1;  wr_cycle[22380] = 1'b0;  addr_rom[22380]='h00001db0;  wr_data_rom[22380]='h00000000;
    rd_cycle[22381] = 1'b1;  wr_cycle[22381] = 1'b0;  addr_rom[22381]='h00001db4;  wr_data_rom[22381]='h00000000;
    rd_cycle[22382] = 1'b1;  wr_cycle[22382] = 1'b0;  addr_rom[22382]='h00001db8;  wr_data_rom[22382]='h00000000;
    rd_cycle[22383] = 1'b1;  wr_cycle[22383] = 1'b0;  addr_rom[22383]='h00001dbc;  wr_data_rom[22383]='h00000000;
    rd_cycle[22384] = 1'b1;  wr_cycle[22384] = 1'b0;  addr_rom[22384]='h00001dc0;  wr_data_rom[22384]='h00000000;
    rd_cycle[22385] = 1'b1;  wr_cycle[22385] = 1'b0;  addr_rom[22385]='h00001dc4;  wr_data_rom[22385]='h00000000;
    rd_cycle[22386] = 1'b1;  wr_cycle[22386] = 1'b0;  addr_rom[22386]='h00001dc8;  wr_data_rom[22386]='h00000000;
    rd_cycle[22387] = 1'b1;  wr_cycle[22387] = 1'b0;  addr_rom[22387]='h00001dcc;  wr_data_rom[22387]='h00000000;
    rd_cycle[22388] = 1'b1;  wr_cycle[22388] = 1'b0;  addr_rom[22388]='h00001dd0;  wr_data_rom[22388]='h00000000;
    rd_cycle[22389] = 1'b1;  wr_cycle[22389] = 1'b0;  addr_rom[22389]='h00001dd4;  wr_data_rom[22389]='h00000000;
    rd_cycle[22390] = 1'b1;  wr_cycle[22390] = 1'b0;  addr_rom[22390]='h00001dd8;  wr_data_rom[22390]='h00000000;
    rd_cycle[22391] = 1'b1;  wr_cycle[22391] = 1'b0;  addr_rom[22391]='h00001ddc;  wr_data_rom[22391]='h00000000;
    rd_cycle[22392] = 1'b1;  wr_cycle[22392] = 1'b0;  addr_rom[22392]='h00001de0;  wr_data_rom[22392]='h00000000;
    rd_cycle[22393] = 1'b1;  wr_cycle[22393] = 1'b0;  addr_rom[22393]='h00001de4;  wr_data_rom[22393]='h00000000;
    rd_cycle[22394] = 1'b1;  wr_cycle[22394] = 1'b0;  addr_rom[22394]='h00001de8;  wr_data_rom[22394]='h00000000;
    rd_cycle[22395] = 1'b1;  wr_cycle[22395] = 1'b0;  addr_rom[22395]='h00001dec;  wr_data_rom[22395]='h00000000;
    rd_cycle[22396] = 1'b1;  wr_cycle[22396] = 1'b0;  addr_rom[22396]='h00001df0;  wr_data_rom[22396]='h00000000;
    rd_cycle[22397] = 1'b1;  wr_cycle[22397] = 1'b0;  addr_rom[22397]='h00001df4;  wr_data_rom[22397]='h00000000;
    rd_cycle[22398] = 1'b1;  wr_cycle[22398] = 1'b0;  addr_rom[22398]='h00001df8;  wr_data_rom[22398]='h00000000;
    rd_cycle[22399] = 1'b1;  wr_cycle[22399] = 1'b0;  addr_rom[22399]='h00001dfc;  wr_data_rom[22399]='h00000000;
    rd_cycle[22400] = 1'b1;  wr_cycle[22400] = 1'b0;  addr_rom[22400]='h00001e00;  wr_data_rom[22400]='h00000000;
    rd_cycle[22401] = 1'b1;  wr_cycle[22401] = 1'b0;  addr_rom[22401]='h00001e04;  wr_data_rom[22401]='h00000000;
    rd_cycle[22402] = 1'b1;  wr_cycle[22402] = 1'b0;  addr_rom[22402]='h00001e08;  wr_data_rom[22402]='h00000000;
    rd_cycle[22403] = 1'b1;  wr_cycle[22403] = 1'b0;  addr_rom[22403]='h00001e0c;  wr_data_rom[22403]='h00000000;
    rd_cycle[22404] = 1'b1;  wr_cycle[22404] = 1'b0;  addr_rom[22404]='h00001e10;  wr_data_rom[22404]='h00000000;
    rd_cycle[22405] = 1'b1;  wr_cycle[22405] = 1'b0;  addr_rom[22405]='h00001e14;  wr_data_rom[22405]='h00000000;
    rd_cycle[22406] = 1'b1;  wr_cycle[22406] = 1'b0;  addr_rom[22406]='h00001e18;  wr_data_rom[22406]='h00000000;
    rd_cycle[22407] = 1'b1;  wr_cycle[22407] = 1'b0;  addr_rom[22407]='h00001e1c;  wr_data_rom[22407]='h00000000;
    rd_cycle[22408] = 1'b1;  wr_cycle[22408] = 1'b0;  addr_rom[22408]='h00001e20;  wr_data_rom[22408]='h00000000;
    rd_cycle[22409] = 1'b1;  wr_cycle[22409] = 1'b0;  addr_rom[22409]='h00001e24;  wr_data_rom[22409]='h00000000;
    rd_cycle[22410] = 1'b1;  wr_cycle[22410] = 1'b0;  addr_rom[22410]='h00001e28;  wr_data_rom[22410]='h00000000;
    rd_cycle[22411] = 1'b1;  wr_cycle[22411] = 1'b0;  addr_rom[22411]='h00001e2c;  wr_data_rom[22411]='h00000000;
    rd_cycle[22412] = 1'b1;  wr_cycle[22412] = 1'b0;  addr_rom[22412]='h00001e30;  wr_data_rom[22412]='h00000000;
    rd_cycle[22413] = 1'b1;  wr_cycle[22413] = 1'b0;  addr_rom[22413]='h00001e34;  wr_data_rom[22413]='h00000000;
    rd_cycle[22414] = 1'b1;  wr_cycle[22414] = 1'b0;  addr_rom[22414]='h00001e38;  wr_data_rom[22414]='h00000000;
    rd_cycle[22415] = 1'b1;  wr_cycle[22415] = 1'b0;  addr_rom[22415]='h00001e3c;  wr_data_rom[22415]='h00000000;
    rd_cycle[22416] = 1'b1;  wr_cycle[22416] = 1'b0;  addr_rom[22416]='h00001e40;  wr_data_rom[22416]='h00000000;
    rd_cycle[22417] = 1'b1;  wr_cycle[22417] = 1'b0;  addr_rom[22417]='h00001e44;  wr_data_rom[22417]='h00000000;
    rd_cycle[22418] = 1'b1;  wr_cycle[22418] = 1'b0;  addr_rom[22418]='h00001e48;  wr_data_rom[22418]='h00000000;
    rd_cycle[22419] = 1'b1;  wr_cycle[22419] = 1'b0;  addr_rom[22419]='h00001e4c;  wr_data_rom[22419]='h00000000;
    rd_cycle[22420] = 1'b1;  wr_cycle[22420] = 1'b0;  addr_rom[22420]='h00001e50;  wr_data_rom[22420]='h00000000;
    rd_cycle[22421] = 1'b1;  wr_cycle[22421] = 1'b0;  addr_rom[22421]='h00001e54;  wr_data_rom[22421]='h00000000;
    rd_cycle[22422] = 1'b1;  wr_cycle[22422] = 1'b0;  addr_rom[22422]='h00001e58;  wr_data_rom[22422]='h00000000;
    rd_cycle[22423] = 1'b1;  wr_cycle[22423] = 1'b0;  addr_rom[22423]='h00001e5c;  wr_data_rom[22423]='h00000000;
    rd_cycle[22424] = 1'b1;  wr_cycle[22424] = 1'b0;  addr_rom[22424]='h00001e60;  wr_data_rom[22424]='h00000000;
    rd_cycle[22425] = 1'b1;  wr_cycle[22425] = 1'b0;  addr_rom[22425]='h00001e64;  wr_data_rom[22425]='h00000000;
    rd_cycle[22426] = 1'b1;  wr_cycle[22426] = 1'b0;  addr_rom[22426]='h00001e68;  wr_data_rom[22426]='h00000000;
    rd_cycle[22427] = 1'b1;  wr_cycle[22427] = 1'b0;  addr_rom[22427]='h00001e6c;  wr_data_rom[22427]='h00000000;
    rd_cycle[22428] = 1'b1;  wr_cycle[22428] = 1'b0;  addr_rom[22428]='h00001e70;  wr_data_rom[22428]='h00000000;
    rd_cycle[22429] = 1'b1;  wr_cycle[22429] = 1'b0;  addr_rom[22429]='h00001e74;  wr_data_rom[22429]='h00000000;
    rd_cycle[22430] = 1'b1;  wr_cycle[22430] = 1'b0;  addr_rom[22430]='h00001e78;  wr_data_rom[22430]='h00000000;
    rd_cycle[22431] = 1'b1;  wr_cycle[22431] = 1'b0;  addr_rom[22431]='h00001e7c;  wr_data_rom[22431]='h00000000;
    rd_cycle[22432] = 1'b1;  wr_cycle[22432] = 1'b0;  addr_rom[22432]='h00001e80;  wr_data_rom[22432]='h00000000;
    rd_cycle[22433] = 1'b1;  wr_cycle[22433] = 1'b0;  addr_rom[22433]='h00001e84;  wr_data_rom[22433]='h00000000;
    rd_cycle[22434] = 1'b1;  wr_cycle[22434] = 1'b0;  addr_rom[22434]='h00001e88;  wr_data_rom[22434]='h00000000;
    rd_cycle[22435] = 1'b1;  wr_cycle[22435] = 1'b0;  addr_rom[22435]='h00001e8c;  wr_data_rom[22435]='h00000000;
    rd_cycle[22436] = 1'b1;  wr_cycle[22436] = 1'b0;  addr_rom[22436]='h00001e90;  wr_data_rom[22436]='h00000000;
    rd_cycle[22437] = 1'b1;  wr_cycle[22437] = 1'b0;  addr_rom[22437]='h00001e94;  wr_data_rom[22437]='h00000000;
    rd_cycle[22438] = 1'b1;  wr_cycle[22438] = 1'b0;  addr_rom[22438]='h00001e98;  wr_data_rom[22438]='h00000000;
    rd_cycle[22439] = 1'b1;  wr_cycle[22439] = 1'b0;  addr_rom[22439]='h00001e9c;  wr_data_rom[22439]='h00000000;
    rd_cycle[22440] = 1'b1;  wr_cycle[22440] = 1'b0;  addr_rom[22440]='h00001ea0;  wr_data_rom[22440]='h00000000;
    rd_cycle[22441] = 1'b1;  wr_cycle[22441] = 1'b0;  addr_rom[22441]='h00001ea4;  wr_data_rom[22441]='h00000000;
    rd_cycle[22442] = 1'b1;  wr_cycle[22442] = 1'b0;  addr_rom[22442]='h00001ea8;  wr_data_rom[22442]='h00000000;
    rd_cycle[22443] = 1'b1;  wr_cycle[22443] = 1'b0;  addr_rom[22443]='h00001eac;  wr_data_rom[22443]='h00000000;
    rd_cycle[22444] = 1'b1;  wr_cycle[22444] = 1'b0;  addr_rom[22444]='h00001eb0;  wr_data_rom[22444]='h00000000;
    rd_cycle[22445] = 1'b1;  wr_cycle[22445] = 1'b0;  addr_rom[22445]='h00001eb4;  wr_data_rom[22445]='h00000000;
    rd_cycle[22446] = 1'b1;  wr_cycle[22446] = 1'b0;  addr_rom[22446]='h00001eb8;  wr_data_rom[22446]='h00000000;
    rd_cycle[22447] = 1'b1;  wr_cycle[22447] = 1'b0;  addr_rom[22447]='h00001ebc;  wr_data_rom[22447]='h00000000;
    rd_cycle[22448] = 1'b1;  wr_cycle[22448] = 1'b0;  addr_rom[22448]='h00001ec0;  wr_data_rom[22448]='h00000000;
    rd_cycle[22449] = 1'b1;  wr_cycle[22449] = 1'b0;  addr_rom[22449]='h00001ec4;  wr_data_rom[22449]='h00000000;
    rd_cycle[22450] = 1'b1;  wr_cycle[22450] = 1'b0;  addr_rom[22450]='h00001ec8;  wr_data_rom[22450]='h00000000;
    rd_cycle[22451] = 1'b1;  wr_cycle[22451] = 1'b0;  addr_rom[22451]='h00001ecc;  wr_data_rom[22451]='h00000000;
    rd_cycle[22452] = 1'b1;  wr_cycle[22452] = 1'b0;  addr_rom[22452]='h00001ed0;  wr_data_rom[22452]='h00000000;
    rd_cycle[22453] = 1'b1;  wr_cycle[22453] = 1'b0;  addr_rom[22453]='h00001ed4;  wr_data_rom[22453]='h00000000;
    rd_cycle[22454] = 1'b1;  wr_cycle[22454] = 1'b0;  addr_rom[22454]='h00001ed8;  wr_data_rom[22454]='h00000000;
    rd_cycle[22455] = 1'b1;  wr_cycle[22455] = 1'b0;  addr_rom[22455]='h00001edc;  wr_data_rom[22455]='h00000000;
    rd_cycle[22456] = 1'b1;  wr_cycle[22456] = 1'b0;  addr_rom[22456]='h00001ee0;  wr_data_rom[22456]='h00000000;
    rd_cycle[22457] = 1'b1;  wr_cycle[22457] = 1'b0;  addr_rom[22457]='h00001ee4;  wr_data_rom[22457]='h00000000;
    rd_cycle[22458] = 1'b1;  wr_cycle[22458] = 1'b0;  addr_rom[22458]='h00001ee8;  wr_data_rom[22458]='h00000000;
    rd_cycle[22459] = 1'b1;  wr_cycle[22459] = 1'b0;  addr_rom[22459]='h00001eec;  wr_data_rom[22459]='h00000000;
    rd_cycle[22460] = 1'b1;  wr_cycle[22460] = 1'b0;  addr_rom[22460]='h00001ef0;  wr_data_rom[22460]='h00000000;
    rd_cycle[22461] = 1'b1;  wr_cycle[22461] = 1'b0;  addr_rom[22461]='h00001ef4;  wr_data_rom[22461]='h00000000;
    rd_cycle[22462] = 1'b1;  wr_cycle[22462] = 1'b0;  addr_rom[22462]='h00001ef8;  wr_data_rom[22462]='h00000000;
    rd_cycle[22463] = 1'b1;  wr_cycle[22463] = 1'b0;  addr_rom[22463]='h00001efc;  wr_data_rom[22463]='h00000000;
    rd_cycle[22464] = 1'b1;  wr_cycle[22464] = 1'b0;  addr_rom[22464]='h00001f00;  wr_data_rom[22464]='h00000000;
    rd_cycle[22465] = 1'b1;  wr_cycle[22465] = 1'b0;  addr_rom[22465]='h00001f04;  wr_data_rom[22465]='h00000000;
    rd_cycle[22466] = 1'b1;  wr_cycle[22466] = 1'b0;  addr_rom[22466]='h00001f08;  wr_data_rom[22466]='h00000000;
    rd_cycle[22467] = 1'b1;  wr_cycle[22467] = 1'b0;  addr_rom[22467]='h00001f0c;  wr_data_rom[22467]='h00000000;
    rd_cycle[22468] = 1'b1;  wr_cycle[22468] = 1'b0;  addr_rom[22468]='h00001f10;  wr_data_rom[22468]='h00000000;
    rd_cycle[22469] = 1'b1;  wr_cycle[22469] = 1'b0;  addr_rom[22469]='h00001f14;  wr_data_rom[22469]='h00000000;
    rd_cycle[22470] = 1'b1;  wr_cycle[22470] = 1'b0;  addr_rom[22470]='h00001f18;  wr_data_rom[22470]='h00000000;
    rd_cycle[22471] = 1'b1;  wr_cycle[22471] = 1'b0;  addr_rom[22471]='h00001f1c;  wr_data_rom[22471]='h00000000;
    rd_cycle[22472] = 1'b1;  wr_cycle[22472] = 1'b0;  addr_rom[22472]='h00001f20;  wr_data_rom[22472]='h00000000;
    rd_cycle[22473] = 1'b1;  wr_cycle[22473] = 1'b0;  addr_rom[22473]='h00001f24;  wr_data_rom[22473]='h00000000;
    rd_cycle[22474] = 1'b1;  wr_cycle[22474] = 1'b0;  addr_rom[22474]='h00001f28;  wr_data_rom[22474]='h00000000;
    rd_cycle[22475] = 1'b1;  wr_cycle[22475] = 1'b0;  addr_rom[22475]='h00001f2c;  wr_data_rom[22475]='h00000000;
    rd_cycle[22476] = 1'b1;  wr_cycle[22476] = 1'b0;  addr_rom[22476]='h00001f30;  wr_data_rom[22476]='h00000000;
    rd_cycle[22477] = 1'b1;  wr_cycle[22477] = 1'b0;  addr_rom[22477]='h00001f34;  wr_data_rom[22477]='h00000000;
    rd_cycle[22478] = 1'b1;  wr_cycle[22478] = 1'b0;  addr_rom[22478]='h00001f38;  wr_data_rom[22478]='h00000000;
    rd_cycle[22479] = 1'b1;  wr_cycle[22479] = 1'b0;  addr_rom[22479]='h00001f3c;  wr_data_rom[22479]='h00000000;
    rd_cycle[22480] = 1'b1;  wr_cycle[22480] = 1'b0;  addr_rom[22480]='h00001f40;  wr_data_rom[22480]='h00000000;
    rd_cycle[22481] = 1'b1;  wr_cycle[22481] = 1'b0;  addr_rom[22481]='h00001f44;  wr_data_rom[22481]='h00000000;
    rd_cycle[22482] = 1'b1;  wr_cycle[22482] = 1'b0;  addr_rom[22482]='h00001f48;  wr_data_rom[22482]='h00000000;
    rd_cycle[22483] = 1'b1;  wr_cycle[22483] = 1'b0;  addr_rom[22483]='h00001f4c;  wr_data_rom[22483]='h00000000;
    rd_cycle[22484] = 1'b1;  wr_cycle[22484] = 1'b0;  addr_rom[22484]='h00001f50;  wr_data_rom[22484]='h00000000;
    rd_cycle[22485] = 1'b1;  wr_cycle[22485] = 1'b0;  addr_rom[22485]='h00001f54;  wr_data_rom[22485]='h00000000;
    rd_cycle[22486] = 1'b1;  wr_cycle[22486] = 1'b0;  addr_rom[22486]='h00001f58;  wr_data_rom[22486]='h00000000;
    rd_cycle[22487] = 1'b1;  wr_cycle[22487] = 1'b0;  addr_rom[22487]='h00001f5c;  wr_data_rom[22487]='h00000000;
    rd_cycle[22488] = 1'b1;  wr_cycle[22488] = 1'b0;  addr_rom[22488]='h00001f60;  wr_data_rom[22488]='h00000000;
    rd_cycle[22489] = 1'b1;  wr_cycle[22489] = 1'b0;  addr_rom[22489]='h00001f64;  wr_data_rom[22489]='h00000000;
    rd_cycle[22490] = 1'b1;  wr_cycle[22490] = 1'b0;  addr_rom[22490]='h00001f68;  wr_data_rom[22490]='h00000000;
    rd_cycle[22491] = 1'b1;  wr_cycle[22491] = 1'b0;  addr_rom[22491]='h00001f6c;  wr_data_rom[22491]='h00000000;
    rd_cycle[22492] = 1'b1;  wr_cycle[22492] = 1'b0;  addr_rom[22492]='h00001f70;  wr_data_rom[22492]='h00000000;
    rd_cycle[22493] = 1'b1;  wr_cycle[22493] = 1'b0;  addr_rom[22493]='h00001f74;  wr_data_rom[22493]='h00000000;
    rd_cycle[22494] = 1'b1;  wr_cycle[22494] = 1'b0;  addr_rom[22494]='h00001f78;  wr_data_rom[22494]='h00000000;
    rd_cycle[22495] = 1'b1;  wr_cycle[22495] = 1'b0;  addr_rom[22495]='h00001f7c;  wr_data_rom[22495]='h00000000;
    rd_cycle[22496] = 1'b1;  wr_cycle[22496] = 1'b0;  addr_rom[22496]='h00001f80;  wr_data_rom[22496]='h00000000;
    rd_cycle[22497] = 1'b1;  wr_cycle[22497] = 1'b0;  addr_rom[22497]='h00001f84;  wr_data_rom[22497]='h00000000;
    rd_cycle[22498] = 1'b1;  wr_cycle[22498] = 1'b0;  addr_rom[22498]='h00001f88;  wr_data_rom[22498]='h00000000;
    rd_cycle[22499] = 1'b1;  wr_cycle[22499] = 1'b0;  addr_rom[22499]='h00001f8c;  wr_data_rom[22499]='h00000000;
    rd_cycle[22500] = 1'b1;  wr_cycle[22500] = 1'b0;  addr_rom[22500]='h00001f90;  wr_data_rom[22500]='h00000000;
    rd_cycle[22501] = 1'b1;  wr_cycle[22501] = 1'b0;  addr_rom[22501]='h00001f94;  wr_data_rom[22501]='h00000000;
    rd_cycle[22502] = 1'b1;  wr_cycle[22502] = 1'b0;  addr_rom[22502]='h00001f98;  wr_data_rom[22502]='h00000000;
    rd_cycle[22503] = 1'b1;  wr_cycle[22503] = 1'b0;  addr_rom[22503]='h00001f9c;  wr_data_rom[22503]='h00000000;
    rd_cycle[22504] = 1'b1;  wr_cycle[22504] = 1'b0;  addr_rom[22504]='h00001fa0;  wr_data_rom[22504]='h00000000;
    rd_cycle[22505] = 1'b1;  wr_cycle[22505] = 1'b0;  addr_rom[22505]='h00001fa4;  wr_data_rom[22505]='h00000000;
    rd_cycle[22506] = 1'b1;  wr_cycle[22506] = 1'b0;  addr_rom[22506]='h00001fa8;  wr_data_rom[22506]='h00000000;
    rd_cycle[22507] = 1'b1;  wr_cycle[22507] = 1'b0;  addr_rom[22507]='h00001fac;  wr_data_rom[22507]='h00000000;
    rd_cycle[22508] = 1'b1;  wr_cycle[22508] = 1'b0;  addr_rom[22508]='h00001fb0;  wr_data_rom[22508]='h00000000;
    rd_cycle[22509] = 1'b1;  wr_cycle[22509] = 1'b0;  addr_rom[22509]='h00001fb4;  wr_data_rom[22509]='h00000000;
    rd_cycle[22510] = 1'b1;  wr_cycle[22510] = 1'b0;  addr_rom[22510]='h00001fb8;  wr_data_rom[22510]='h00000000;
    rd_cycle[22511] = 1'b1;  wr_cycle[22511] = 1'b0;  addr_rom[22511]='h00001fbc;  wr_data_rom[22511]='h00000000;
    rd_cycle[22512] = 1'b1;  wr_cycle[22512] = 1'b0;  addr_rom[22512]='h00001fc0;  wr_data_rom[22512]='h00000000;
    rd_cycle[22513] = 1'b1;  wr_cycle[22513] = 1'b0;  addr_rom[22513]='h00001fc4;  wr_data_rom[22513]='h00000000;
    rd_cycle[22514] = 1'b1;  wr_cycle[22514] = 1'b0;  addr_rom[22514]='h00001fc8;  wr_data_rom[22514]='h00000000;
    rd_cycle[22515] = 1'b1;  wr_cycle[22515] = 1'b0;  addr_rom[22515]='h00001fcc;  wr_data_rom[22515]='h00000000;
    rd_cycle[22516] = 1'b1;  wr_cycle[22516] = 1'b0;  addr_rom[22516]='h00001fd0;  wr_data_rom[22516]='h00000000;
    rd_cycle[22517] = 1'b1;  wr_cycle[22517] = 1'b0;  addr_rom[22517]='h00001fd4;  wr_data_rom[22517]='h00000000;
    rd_cycle[22518] = 1'b1;  wr_cycle[22518] = 1'b0;  addr_rom[22518]='h00001fd8;  wr_data_rom[22518]='h00000000;
    rd_cycle[22519] = 1'b1;  wr_cycle[22519] = 1'b0;  addr_rom[22519]='h00001fdc;  wr_data_rom[22519]='h00000000;
    rd_cycle[22520] = 1'b1;  wr_cycle[22520] = 1'b0;  addr_rom[22520]='h00001fe0;  wr_data_rom[22520]='h00000000;
    rd_cycle[22521] = 1'b1;  wr_cycle[22521] = 1'b0;  addr_rom[22521]='h00001fe4;  wr_data_rom[22521]='h00000000;
    rd_cycle[22522] = 1'b1;  wr_cycle[22522] = 1'b0;  addr_rom[22522]='h00001fe8;  wr_data_rom[22522]='h00000000;
    rd_cycle[22523] = 1'b1;  wr_cycle[22523] = 1'b0;  addr_rom[22523]='h00001fec;  wr_data_rom[22523]='h00000000;
    rd_cycle[22524] = 1'b1;  wr_cycle[22524] = 1'b0;  addr_rom[22524]='h00001ff0;  wr_data_rom[22524]='h00000000;
    rd_cycle[22525] = 1'b1;  wr_cycle[22525] = 1'b0;  addr_rom[22525]='h00001ff4;  wr_data_rom[22525]='h00000000;
    rd_cycle[22526] = 1'b1;  wr_cycle[22526] = 1'b0;  addr_rom[22526]='h00001ff8;  wr_data_rom[22526]='h00000000;
    rd_cycle[22527] = 1'b1;  wr_cycle[22527] = 1'b0;  addr_rom[22527]='h00001ffc;  wr_data_rom[22527]='h00000000;
    rd_cycle[22528] = 1'b1;  wr_cycle[22528] = 1'b0;  addr_rom[22528]='h00002000;  wr_data_rom[22528]='h00000000;
    rd_cycle[22529] = 1'b1;  wr_cycle[22529] = 1'b0;  addr_rom[22529]='h00002004;  wr_data_rom[22529]='h00000000;
    rd_cycle[22530] = 1'b1;  wr_cycle[22530] = 1'b0;  addr_rom[22530]='h00002008;  wr_data_rom[22530]='h00000000;
    rd_cycle[22531] = 1'b1;  wr_cycle[22531] = 1'b0;  addr_rom[22531]='h0000200c;  wr_data_rom[22531]='h00000000;
    rd_cycle[22532] = 1'b1;  wr_cycle[22532] = 1'b0;  addr_rom[22532]='h00002010;  wr_data_rom[22532]='h00000000;
    rd_cycle[22533] = 1'b1;  wr_cycle[22533] = 1'b0;  addr_rom[22533]='h00002014;  wr_data_rom[22533]='h00000000;
    rd_cycle[22534] = 1'b1;  wr_cycle[22534] = 1'b0;  addr_rom[22534]='h00002018;  wr_data_rom[22534]='h00000000;
    rd_cycle[22535] = 1'b1;  wr_cycle[22535] = 1'b0;  addr_rom[22535]='h0000201c;  wr_data_rom[22535]='h00000000;
    rd_cycle[22536] = 1'b1;  wr_cycle[22536] = 1'b0;  addr_rom[22536]='h00002020;  wr_data_rom[22536]='h00000000;
    rd_cycle[22537] = 1'b1;  wr_cycle[22537] = 1'b0;  addr_rom[22537]='h00002024;  wr_data_rom[22537]='h00000000;
    rd_cycle[22538] = 1'b1;  wr_cycle[22538] = 1'b0;  addr_rom[22538]='h00002028;  wr_data_rom[22538]='h00000000;
    rd_cycle[22539] = 1'b1;  wr_cycle[22539] = 1'b0;  addr_rom[22539]='h0000202c;  wr_data_rom[22539]='h00000000;
    rd_cycle[22540] = 1'b1;  wr_cycle[22540] = 1'b0;  addr_rom[22540]='h00002030;  wr_data_rom[22540]='h00000000;
    rd_cycle[22541] = 1'b1;  wr_cycle[22541] = 1'b0;  addr_rom[22541]='h00002034;  wr_data_rom[22541]='h00000000;
    rd_cycle[22542] = 1'b1;  wr_cycle[22542] = 1'b0;  addr_rom[22542]='h00002038;  wr_data_rom[22542]='h00000000;
    rd_cycle[22543] = 1'b1;  wr_cycle[22543] = 1'b0;  addr_rom[22543]='h0000203c;  wr_data_rom[22543]='h00000000;
    rd_cycle[22544] = 1'b1;  wr_cycle[22544] = 1'b0;  addr_rom[22544]='h00002040;  wr_data_rom[22544]='h00000000;
    rd_cycle[22545] = 1'b1;  wr_cycle[22545] = 1'b0;  addr_rom[22545]='h00002044;  wr_data_rom[22545]='h00000000;
    rd_cycle[22546] = 1'b1;  wr_cycle[22546] = 1'b0;  addr_rom[22546]='h00002048;  wr_data_rom[22546]='h00000000;
    rd_cycle[22547] = 1'b1;  wr_cycle[22547] = 1'b0;  addr_rom[22547]='h0000204c;  wr_data_rom[22547]='h00000000;
    rd_cycle[22548] = 1'b1;  wr_cycle[22548] = 1'b0;  addr_rom[22548]='h00002050;  wr_data_rom[22548]='h00000000;
    rd_cycle[22549] = 1'b1;  wr_cycle[22549] = 1'b0;  addr_rom[22549]='h00002054;  wr_data_rom[22549]='h00000000;
    rd_cycle[22550] = 1'b1;  wr_cycle[22550] = 1'b0;  addr_rom[22550]='h00002058;  wr_data_rom[22550]='h00000000;
    rd_cycle[22551] = 1'b1;  wr_cycle[22551] = 1'b0;  addr_rom[22551]='h0000205c;  wr_data_rom[22551]='h00000000;
    rd_cycle[22552] = 1'b1;  wr_cycle[22552] = 1'b0;  addr_rom[22552]='h00002060;  wr_data_rom[22552]='h00000000;
    rd_cycle[22553] = 1'b1;  wr_cycle[22553] = 1'b0;  addr_rom[22553]='h00002064;  wr_data_rom[22553]='h00000000;
    rd_cycle[22554] = 1'b1;  wr_cycle[22554] = 1'b0;  addr_rom[22554]='h00002068;  wr_data_rom[22554]='h00000000;
    rd_cycle[22555] = 1'b1;  wr_cycle[22555] = 1'b0;  addr_rom[22555]='h0000206c;  wr_data_rom[22555]='h00000000;
    rd_cycle[22556] = 1'b1;  wr_cycle[22556] = 1'b0;  addr_rom[22556]='h00002070;  wr_data_rom[22556]='h00000000;
    rd_cycle[22557] = 1'b1;  wr_cycle[22557] = 1'b0;  addr_rom[22557]='h00002074;  wr_data_rom[22557]='h00000000;
    rd_cycle[22558] = 1'b1;  wr_cycle[22558] = 1'b0;  addr_rom[22558]='h00002078;  wr_data_rom[22558]='h00000000;
    rd_cycle[22559] = 1'b1;  wr_cycle[22559] = 1'b0;  addr_rom[22559]='h0000207c;  wr_data_rom[22559]='h00000000;
    rd_cycle[22560] = 1'b1;  wr_cycle[22560] = 1'b0;  addr_rom[22560]='h00002080;  wr_data_rom[22560]='h00000000;
    rd_cycle[22561] = 1'b1;  wr_cycle[22561] = 1'b0;  addr_rom[22561]='h00002084;  wr_data_rom[22561]='h00000000;
    rd_cycle[22562] = 1'b1;  wr_cycle[22562] = 1'b0;  addr_rom[22562]='h00002088;  wr_data_rom[22562]='h00000000;
    rd_cycle[22563] = 1'b1;  wr_cycle[22563] = 1'b0;  addr_rom[22563]='h0000208c;  wr_data_rom[22563]='h00000000;
    rd_cycle[22564] = 1'b1;  wr_cycle[22564] = 1'b0;  addr_rom[22564]='h00002090;  wr_data_rom[22564]='h00000000;
    rd_cycle[22565] = 1'b1;  wr_cycle[22565] = 1'b0;  addr_rom[22565]='h00002094;  wr_data_rom[22565]='h00000000;
    rd_cycle[22566] = 1'b1;  wr_cycle[22566] = 1'b0;  addr_rom[22566]='h00002098;  wr_data_rom[22566]='h00000000;
    rd_cycle[22567] = 1'b1;  wr_cycle[22567] = 1'b0;  addr_rom[22567]='h0000209c;  wr_data_rom[22567]='h00000000;
    rd_cycle[22568] = 1'b1;  wr_cycle[22568] = 1'b0;  addr_rom[22568]='h000020a0;  wr_data_rom[22568]='h00000000;
    rd_cycle[22569] = 1'b1;  wr_cycle[22569] = 1'b0;  addr_rom[22569]='h000020a4;  wr_data_rom[22569]='h00000000;
    rd_cycle[22570] = 1'b1;  wr_cycle[22570] = 1'b0;  addr_rom[22570]='h000020a8;  wr_data_rom[22570]='h00000000;
    rd_cycle[22571] = 1'b1;  wr_cycle[22571] = 1'b0;  addr_rom[22571]='h000020ac;  wr_data_rom[22571]='h00000000;
    rd_cycle[22572] = 1'b1;  wr_cycle[22572] = 1'b0;  addr_rom[22572]='h000020b0;  wr_data_rom[22572]='h00000000;
    rd_cycle[22573] = 1'b1;  wr_cycle[22573] = 1'b0;  addr_rom[22573]='h000020b4;  wr_data_rom[22573]='h00000000;
    rd_cycle[22574] = 1'b1;  wr_cycle[22574] = 1'b0;  addr_rom[22574]='h000020b8;  wr_data_rom[22574]='h00000000;
    rd_cycle[22575] = 1'b1;  wr_cycle[22575] = 1'b0;  addr_rom[22575]='h000020bc;  wr_data_rom[22575]='h00000000;
    rd_cycle[22576] = 1'b1;  wr_cycle[22576] = 1'b0;  addr_rom[22576]='h000020c0;  wr_data_rom[22576]='h00000000;
    rd_cycle[22577] = 1'b1;  wr_cycle[22577] = 1'b0;  addr_rom[22577]='h000020c4;  wr_data_rom[22577]='h00000000;
    rd_cycle[22578] = 1'b1;  wr_cycle[22578] = 1'b0;  addr_rom[22578]='h000020c8;  wr_data_rom[22578]='h00000000;
    rd_cycle[22579] = 1'b1;  wr_cycle[22579] = 1'b0;  addr_rom[22579]='h000020cc;  wr_data_rom[22579]='h00000000;
    rd_cycle[22580] = 1'b1;  wr_cycle[22580] = 1'b0;  addr_rom[22580]='h000020d0;  wr_data_rom[22580]='h00000000;
    rd_cycle[22581] = 1'b1;  wr_cycle[22581] = 1'b0;  addr_rom[22581]='h000020d4;  wr_data_rom[22581]='h00000000;
    rd_cycle[22582] = 1'b1;  wr_cycle[22582] = 1'b0;  addr_rom[22582]='h000020d8;  wr_data_rom[22582]='h00000000;
    rd_cycle[22583] = 1'b1;  wr_cycle[22583] = 1'b0;  addr_rom[22583]='h000020dc;  wr_data_rom[22583]='h00000000;
    rd_cycle[22584] = 1'b1;  wr_cycle[22584] = 1'b0;  addr_rom[22584]='h000020e0;  wr_data_rom[22584]='h00000000;
    rd_cycle[22585] = 1'b1;  wr_cycle[22585] = 1'b0;  addr_rom[22585]='h000020e4;  wr_data_rom[22585]='h00000000;
    rd_cycle[22586] = 1'b1;  wr_cycle[22586] = 1'b0;  addr_rom[22586]='h000020e8;  wr_data_rom[22586]='h00000000;
    rd_cycle[22587] = 1'b1;  wr_cycle[22587] = 1'b0;  addr_rom[22587]='h000020ec;  wr_data_rom[22587]='h00000000;
    rd_cycle[22588] = 1'b1;  wr_cycle[22588] = 1'b0;  addr_rom[22588]='h000020f0;  wr_data_rom[22588]='h00000000;
    rd_cycle[22589] = 1'b1;  wr_cycle[22589] = 1'b0;  addr_rom[22589]='h000020f4;  wr_data_rom[22589]='h00000000;
    rd_cycle[22590] = 1'b1;  wr_cycle[22590] = 1'b0;  addr_rom[22590]='h000020f8;  wr_data_rom[22590]='h00000000;
    rd_cycle[22591] = 1'b1;  wr_cycle[22591] = 1'b0;  addr_rom[22591]='h000020fc;  wr_data_rom[22591]='h00000000;
    rd_cycle[22592] = 1'b1;  wr_cycle[22592] = 1'b0;  addr_rom[22592]='h00002100;  wr_data_rom[22592]='h00000000;
    rd_cycle[22593] = 1'b1;  wr_cycle[22593] = 1'b0;  addr_rom[22593]='h00002104;  wr_data_rom[22593]='h00000000;
    rd_cycle[22594] = 1'b1;  wr_cycle[22594] = 1'b0;  addr_rom[22594]='h00002108;  wr_data_rom[22594]='h00000000;
    rd_cycle[22595] = 1'b1;  wr_cycle[22595] = 1'b0;  addr_rom[22595]='h0000210c;  wr_data_rom[22595]='h00000000;
    rd_cycle[22596] = 1'b1;  wr_cycle[22596] = 1'b0;  addr_rom[22596]='h00002110;  wr_data_rom[22596]='h00000000;
    rd_cycle[22597] = 1'b1;  wr_cycle[22597] = 1'b0;  addr_rom[22597]='h00002114;  wr_data_rom[22597]='h00000000;
    rd_cycle[22598] = 1'b1;  wr_cycle[22598] = 1'b0;  addr_rom[22598]='h00002118;  wr_data_rom[22598]='h00000000;
    rd_cycle[22599] = 1'b1;  wr_cycle[22599] = 1'b0;  addr_rom[22599]='h0000211c;  wr_data_rom[22599]='h00000000;
    rd_cycle[22600] = 1'b1;  wr_cycle[22600] = 1'b0;  addr_rom[22600]='h00002120;  wr_data_rom[22600]='h00000000;
    rd_cycle[22601] = 1'b1;  wr_cycle[22601] = 1'b0;  addr_rom[22601]='h00002124;  wr_data_rom[22601]='h00000000;
    rd_cycle[22602] = 1'b1;  wr_cycle[22602] = 1'b0;  addr_rom[22602]='h00002128;  wr_data_rom[22602]='h00000000;
    rd_cycle[22603] = 1'b1;  wr_cycle[22603] = 1'b0;  addr_rom[22603]='h0000212c;  wr_data_rom[22603]='h00000000;
    rd_cycle[22604] = 1'b1;  wr_cycle[22604] = 1'b0;  addr_rom[22604]='h00002130;  wr_data_rom[22604]='h00000000;
    rd_cycle[22605] = 1'b1;  wr_cycle[22605] = 1'b0;  addr_rom[22605]='h00002134;  wr_data_rom[22605]='h00000000;
    rd_cycle[22606] = 1'b1;  wr_cycle[22606] = 1'b0;  addr_rom[22606]='h00002138;  wr_data_rom[22606]='h00000000;
    rd_cycle[22607] = 1'b1;  wr_cycle[22607] = 1'b0;  addr_rom[22607]='h0000213c;  wr_data_rom[22607]='h00000000;
    rd_cycle[22608] = 1'b1;  wr_cycle[22608] = 1'b0;  addr_rom[22608]='h00002140;  wr_data_rom[22608]='h00000000;
    rd_cycle[22609] = 1'b1;  wr_cycle[22609] = 1'b0;  addr_rom[22609]='h00002144;  wr_data_rom[22609]='h00000000;
    rd_cycle[22610] = 1'b1;  wr_cycle[22610] = 1'b0;  addr_rom[22610]='h00002148;  wr_data_rom[22610]='h00000000;
    rd_cycle[22611] = 1'b1;  wr_cycle[22611] = 1'b0;  addr_rom[22611]='h0000214c;  wr_data_rom[22611]='h00000000;
    rd_cycle[22612] = 1'b1;  wr_cycle[22612] = 1'b0;  addr_rom[22612]='h00002150;  wr_data_rom[22612]='h00000000;
    rd_cycle[22613] = 1'b1;  wr_cycle[22613] = 1'b0;  addr_rom[22613]='h00002154;  wr_data_rom[22613]='h00000000;
    rd_cycle[22614] = 1'b1;  wr_cycle[22614] = 1'b0;  addr_rom[22614]='h00002158;  wr_data_rom[22614]='h00000000;
    rd_cycle[22615] = 1'b1;  wr_cycle[22615] = 1'b0;  addr_rom[22615]='h0000215c;  wr_data_rom[22615]='h00000000;
    rd_cycle[22616] = 1'b1;  wr_cycle[22616] = 1'b0;  addr_rom[22616]='h00002160;  wr_data_rom[22616]='h00000000;
    rd_cycle[22617] = 1'b1;  wr_cycle[22617] = 1'b0;  addr_rom[22617]='h00002164;  wr_data_rom[22617]='h00000000;
    rd_cycle[22618] = 1'b1;  wr_cycle[22618] = 1'b0;  addr_rom[22618]='h00002168;  wr_data_rom[22618]='h00000000;
    rd_cycle[22619] = 1'b1;  wr_cycle[22619] = 1'b0;  addr_rom[22619]='h0000216c;  wr_data_rom[22619]='h00000000;
    rd_cycle[22620] = 1'b1;  wr_cycle[22620] = 1'b0;  addr_rom[22620]='h00002170;  wr_data_rom[22620]='h00000000;
    rd_cycle[22621] = 1'b1;  wr_cycle[22621] = 1'b0;  addr_rom[22621]='h00002174;  wr_data_rom[22621]='h00000000;
    rd_cycle[22622] = 1'b1;  wr_cycle[22622] = 1'b0;  addr_rom[22622]='h00002178;  wr_data_rom[22622]='h00000000;
    rd_cycle[22623] = 1'b1;  wr_cycle[22623] = 1'b0;  addr_rom[22623]='h0000217c;  wr_data_rom[22623]='h00000000;
    rd_cycle[22624] = 1'b1;  wr_cycle[22624] = 1'b0;  addr_rom[22624]='h00002180;  wr_data_rom[22624]='h00000000;
    rd_cycle[22625] = 1'b1;  wr_cycle[22625] = 1'b0;  addr_rom[22625]='h00002184;  wr_data_rom[22625]='h00000000;
    rd_cycle[22626] = 1'b1;  wr_cycle[22626] = 1'b0;  addr_rom[22626]='h00002188;  wr_data_rom[22626]='h00000000;
    rd_cycle[22627] = 1'b1;  wr_cycle[22627] = 1'b0;  addr_rom[22627]='h0000218c;  wr_data_rom[22627]='h00000000;
    rd_cycle[22628] = 1'b1;  wr_cycle[22628] = 1'b0;  addr_rom[22628]='h00002190;  wr_data_rom[22628]='h00000000;
    rd_cycle[22629] = 1'b1;  wr_cycle[22629] = 1'b0;  addr_rom[22629]='h00002194;  wr_data_rom[22629]='h00000000;
    rd_cycle[22630] = 1'b1;  wr_cycle[22630] = 1'b0;  addr_rom[22630]='h00002198;  wr_data_rom[22630]='h00000000;
    rd_cycle[22631] = 1'b1;  wr_cycle[22631] = 1'b0;  addr_rom[22631]='h0000219c;  wr_data_rom[22631]='h00000000;
    rd_cycle[22632] = 1'b1;  wr_cycle[22632] = 1'b0;  addr_rom[22632]='h000021a0;  wr_data_rom[22632]='h00000000;
    rd_cycle[22633] = 1'b1;  wr_cycle[22633] = 1'b0;  addr_rom[22633]='h000021a4;  wr_data_rom[22633]='h00000000;
    rd_cycle[22634] = 1'b1;  wr_cycle[22634] = 1'b0;  addr_rom[22634]='h000021a8;  wr_data_rom[22634]='h00000000;
    rd_cycle[22635] = 1'b1;  wr_cycle[22635] = 1'b0;  addr_rom[22635]='h000021ac;  wr_data_rom[22635]='h00000000;
    rd_cycle[22636] = 1'b1;  wr_cycle[22636] = 1'b0;  addr_rom[22636]='h000021b0;  wr_data_rom[22636]='h00000000;
    rd_cycle[22637] = 1'b1;  wr_cycle[22637] = 1'b0;  addr_rom[22637]='h000021b4;  wr_data_rom[22637]='h00000000;
    rd_cycle[22638] = 1'b1;  wr_cycle[22638] = 1'b0;  addr_rom[22638]='h000021b8;  wr_data_rom[22638]='h00000000;
    rd_cycle[22639] = 1'b1;  wr_cycle[22639] = 1'b0;  addr_rom[22639]='h000021bc;  wr_data_rom[22639]='h00000000;
    rd_cycle[22640] = 1'b1;  wr_cycle[22640] = 1'b0;  addr_rom[22640]='h000021c0;  wr_data_rom[22640]='h00000000;
    rd_cycle[22641] = 1'b1;  wr_cycle[22641] = 1'b0;  addr_rom[22641]='h000021c4;  wr_data_rom[22641]='h00000000;
    rd_cycle[22642] = 1'b1;  wr_cycle[22642] = 1'b0;  addr_rom[22642]='h000021c8;  wr_data_rom[22642]='h00000000;
    rd_cycle[22643] = 1'b1;  wr_cycle[22643] = 1'b0;  addr_rom[22643]='h000021cc;  wr_data_rom[22643]='h00000000;
    rd_cycle[22644] = 1'b1;  wr_cycle[22644] = 1'b0;  addr_rom[22644]='h000021d0;  wr_data_rom[22644]='h00000000;
    rd_cycle[22645] = 1'b1;  wr_cycle[22645] = 1'b0;  addr_rom[22645]='h000021d4;  wr_data_rom[22645]='h00000000;
    rd_cycle[22646] = 1'b1;  wr_cycle[22646] = 1'b0;  addr_rom[22646]='h000021d8;  wr_data_rom[22646]='h00000000;
    rd_cycle[22647] = 1'b1;  wr_cycle[22647] = 1'b0;  addr_rom[22647]='h000021dc;  wr_data_rom[22647]='h00000000;
    rd_cycle[22648] = 1'b1;  wr_cycle[22648] = 1'b0;  addr_rom[22648]='h000021e0;  wr_data_rom[22648]='h00000000;
    rd_cycle[22649] = 1'b1;  wr_cycle[22649] = 1'b0;  addr_rom[22649]='h000021e4;  wr_data_rom[22649]='h00000000;
    rd_cycle[22650] = 1'b1;  wr_cycle[22650] = 1'b0;  addr_rom[22650]='h000021e8;  wr_data_rom[22650]='h00000000;
    rd_cycle[22651] = 1'b1;  wr_cycle[22651] = 1'b0;  addr_rom[22651]='h000021ec;  wr_data_rom[22651]='h00000000;
    rd_cycle[22652] = 1'b1;  wr_cycle[22652] = 1'b0;  addr_rom[22652]='h000021f0;  wr_data_rom[22652]='h00000000;
    rd_cycle[22653] = 1'b1;  wr_cycle[22653] = 1'b0;  addr_rom[22653]='h000021f4;  wr_data_rom[22653]='h00000000;
    rd_cycle[22654] = 1'b1;  wr_cycle[22654] = 1'b0;  addr_rom[22654]='h000021f8;  wr_data_rom[22654]='h00000000;
    rd_cycle[22655] = 1'b1;  wr_cycle[22655] = 1'b0;  addr_rom[22655]='h000021fc;  wr_data_rom[22655]='h00000000;
    rd_cycle[22656] = 1'b1;  wr_cycle[22656] = 1'b0;  addr_rom[22656]='h00002200;  wr_data_rom[22656]='h00000000;
    rd_cycle[22657] = 1'b1;  wr_cycle[22657] = 1'b0;  addr_rom[22657]='h00002204;  wr_data_rom[22657]='h00000000;
    rd_cycle[22658] = 1'b1;  wr_cycle[22658] = 1'b0;  addr_rom[22658]='h00002208;  wr_data_rom[22658]='h00000000;
    rd_cycle[22659] = 1'b1;  wr_cycle[22659] = 1'b0;  addr_rom[22659]='h0000220c;  wr_data_rom[22659]='h00000000;
    rd_cycle[22660] = 1'b1;  wr_cycle[22660] = 1'b0;  addr_rom[22660]='h00002210;  wr_data_rom[22660]='h00000000;
    rd_cycle[22661] = 1'b1;  wr_cycle[22661] = 1'b0;  addr_rom[22661]='h00002214;  wr_data_rom[22661]='h00000000;
    rd_cycle[22662] = 1'b1;  wr_cycle[22662] = 1'b0;  addr_rom[22662]='h00002218;  wr_data_rom[22662]='h00000000;
    rd_cycle[22663] = 1'b1;  wr_cycle[22663] = 1'b0;  addr_rom[22663]='h0000221c;  wr_data_rom[22663]='h00000000;
    rd_cycle[22664] = 1'b1;  wr_cycle[22664] = 1'b0;  addr_rom[22664]='h00002220;  wr_data_rom[22664]='h00000000;
    rd_cycle[22665] = 1'b1;  wr_cycle[22665] = 1'b0;  addr_rom[22665]='h00002224;  wr_data_rom[22665]='h00000000;
    rd_cycle[22666] = 1'b1;  wr_cycle[22666] = 1'b0;  addr_rom[22666]='h00002228;  wr_data_rom[22666]='h00000000;
    rd_cycle[22667] = 1'b1;  wr_cycle[22667] = 1'b0;  addr_rom[22667]='h0000222c;  wr_data_rom[22667]='h00000000;
    rd_cycle[22668] = 1'b1;  wr_cycle[22668] = 1'b0;  addr_rom[22668]='h00002230;  wr_data_rom[22668]='h00000000;
    rd_cycle[22669] = 1'b1;  wr_cycle[22669] = 1'b0;  addr_rom[22669]='h00002234;  wr_data_rom[22669]='h00000000;
    rd_cycle[22670] = 1'b1;  wr_cycle[22670] = 1'b0;  addr_rom[22670]='h00002238;  wr_data_rom[22670]='h00000000;
    rd_cycle[22671] = 1'b1;  wr_cycle[22671] = 1'b0;  addr_rom[22671]='h0000223c;  wr_data_rom[22671]='h00000000;
    rd_cycle[22672] = 1'b1;  wr_cycle[22672] = 1'b0;  addr_rom[22672]='h00002240;  wr_data_rom[22672]='h00000000;
    rd_cycle[22673] = 1'b1;  wr_cycle[22673] = 1'b0;  addr_rom[22673]='h00002244;  wr_data_rom[22673]='h00000000;
    rd_cycle[22674] = 1'b1;  wr_cycle[22674] = 1'b0;  addr_rom[22674]='h00002248;  wr_data_rom[22674]='h00000000;
    rd_cycle[22675] = 1'b1;  wr_cycle[22675] = 1'b0;  addr_rom[22675]='h0000224c;  wr_data_rom[22675]='h00000000;
    rd_cycle[22676] = 1'b1;  wr_cycle[22676] = 1'b0;  addr_rom[22676]='h00002250;  wr_data_rom[22676]='h00000000;
    rd_cycle[22677] = 1'b1;  wr_cycle[22677] = 1'b0;  addr_rom[22677]='h00002254;  wr_data_rom[22677]='h00000000;
    rd_cycle[22678] = 1'b1;  wr_cycle[22678] = 1'b0;  addr_rom[22678]='h00002258;  wr_data_rom[22678]='h00000000;
    rd_cycle[22679] = 1'b1;  wr_cycle[22679] = 1'b0;  addr_rom[22679]='h0000225c;  wr_data_rom[22679]='h00000000;
    rd_cycle[22680] = 1'b1;  wr_cycle[22680] = 1'b0;  addr_rom[22680]='h00002260;  wr_data_rom[22680]='h00000000;
    rd_cycle[22681] = 1'b1;  wr_cycle[22681] = 1'b0;  addr_rom[22681]='h00002264;  wr_data_rom[22681]='h00000000;
    rd_cycle[22682] = 1'b1;  wr_cycle[22682] = 1'b0;  addr_rom[22682]='h00002268;  wr_data_rom[22682]='h00000000;
    rd_cycle[22683] = 1'b1;  wr_cycle[22683] = 1'b0;  addr_rom[22683]='h0000226c;  wr_data_rom[22683]='h00000000;
    rd_cycle[22684] = 1'b1;  wr_cycle[22684] = 1'b0;  addr_rom[22684]='h00002270;  wr_data_rom[22684]='h00000000;
    rd_cycle[22685] = 1'b1;  wr_cycle[22685] = 1'b0;  addr_rom[22685]='h00002274;  wr_data_rom[22685]='h00000000;
    rd_cycle[22686] = 1'b1;  wr_cycle[22686] = 1'b0;  addr_rom[22686]='h00002278;  wr_data_rom[22686]='h00000000;
    rd_cycle[22687] = 1'b1;  wr_cycle[22687] = 1'b0;  addr_rom[22687]='h0000227c;  wr_data_rom[22687]='h00000000;
    rd_cycle[22688] = 1'b1;  wr_cycle[22688] = 1'b0;  addr_rom[22688]='h00002280;  wr_data_rom[22688]='h00000000;
    rd_cycle[22689] = 1'b1;  wr_cycle[22689] = 1'b0;  addr_rom[22689]='h00002284;  wr_data_rom[22689]='h00000000;
    rd_cycle[22690] = 1'b1;  wr_cycle[22690] = 1'b0;  addr_rom[22690]='h00002288;  wr_data_rom[22690]='h00000000;
    rd_cycle[22691] = 1'b1;  wr_cycle[22691] = 1'b0;  addr_rom[22691]='h0000228c;  wr_data_rom[22691]='h00000000;
    rd_cycle[22692] = 1'b1;  wr_cycle[22692] = 1'b0;  addr_rom[22692]='h00002290;  wr_data_rom[22692]='h00000000;
    rd_cycle[22693] = 1'b1;  wr_cycle[22693] = 1'b0;  addr_rom[22693]='h00002294;  wr_data_rom[22693]='h00000000;
    rd_cycle[22694] = 1'b1;  wr_cycle[22694] = 1'b0;  addr_rom[22694]='h00002298;  wr_data_rom[22694]='h00000000;
    rd_cycle[22695] = 1'b1;  wr_cycle[22695] = 1'b0;  addr_rom[22695]='h0000229c;  wr_data_rom[22695]='h00000000;
    rd_cycle[22696] = 1'b1;  wr_cycle[22696] = 1'b0;  addr_rom[22696]='h000022a0;  wr_data_rom[22696]='h00000000;
    rd_cycle[22697] = 1'b1;  wr_cycle[22697] = 1'b0;  addr_rom[22697]='h000022a4;  wr_data_rom[22697]='h00000000;
    rd_cycle[22698] = 1'b1;  wr_cycle[22698] = 1'b0;  addr_rom[22698]='h000022a8;  wr_data_rom[22698]='h00000000;
    rd_cycle[22699] = 1'b1;  wr_cycle[22699] = 1'b0;  addr_rom[22699]='h000022ac;  wr_data_rom[22699]='h00000000;
    rd_cycle[22700] = 1'b1;  wr_cycle[22700] = 1'b0;  addr_rom[22700]='h000022b0;  wr_data_rom[22700]='h00000000;
    rd_cycle[22701] = 1'b1;  wr_cycle[22701] = 1'b0;  addr_rom[22701]='h000022b4;  wr_data_rom[22701]='h00000000;
    rd_cycle[22702] = 1'b1;  wr_cycle[22702] = 1'b0;  addr_rom[22702]='h000022b8;  wr_data_rom[22702]='h00000000;
    rd_cycle[22703] = 1'b1;  wr_cycle[22703] = 1'b0;  addr_rom[22703]='h000022bc;  wr_data_rom[22703]='h00000000;
    rd_cycle[22704] = 1'b1;  wr_cycle[22704] = 1'b0;  addr_rom[22704]='h000022c0;  wr_data_rom[22704]='h00000000;
    rd_cycle[22705] = 1'b1;  wr_cycle[22705] = 1'b0;  addr_rom[22705]='h000022c4;  wr_data_rom[22705]='h00000000;
    rd_cycle[22706] = 1'b1;  wr_cycle[22706] = 1'b0;  addr_rom[22706]='h000022c8;  wr_data_rom[22706]='h00000000;
    rd_cycle[22707] = 1'b1;  wr_cycle[22707] = 1'b0;  addr_rom[22707]='h000022cc;  wr_data_rom[22707]='h00000000;
    rd_cycle[22708] = 1'b1;  wr_cycle[22708] = 1'b0;  addr_rom[22708]='h000022d0;  wr_data_rom[22708]='h00000000;
    rd_cycle[22709] = 1'b1;  wr_cycle[22709] = 1'b0;  addr_rom[22709]='h000022d4;  wr_data_rom[22709]='h00000000;
    rd_cycle[22710] = 1'b1;  wr_cycle[22710] = 1'b0;  addr_rom[22710]='h000022d8;  wr_data_rom[22710]='h00000000;
    rd_cycle[22711] = 1'b1;  wr_cycle[22711] = 1'b0;  addr_rom[22711]='h000022dc;  wr_data_rom[22711]='h00000000;
    rd_cycle[22712] = 1'b1;  wr_cycle[22712] = 1'b0;  addr_rom[22712]='h000022e0;  wr_data_rom[22712]='h00000000;
    rd_cycle[22713] = 1'b1;  wr_cycle[22713] = 1'b0;  addr_rom[22713]='h000022e4;  wr_data_rom[22713]='h00000000;
    rd_cycle[22714] = 1'b1;  wr_cycle[22714] = 1'b0;  addr_rom[22714]='h000022e8;  wr_data_rom[22714]='h00000000;
    rd_cycle[22715] = 1'b1;  wr_cycle[22715] = 1'b0;  addr_rom[22715]='h000022ec;  wr_data_rom[22715]='h00000000;
    rd_cycle[22716] = 1'b1;  wr_cycle[22716] = 1'b0;  addr_rom[22716]='h000022f0;  wr_data_rom[22716]='h00000000;
    rd_cycle[22717] = 1'b1;  wr_cycle[22717] = 1'b0;  addr_rom[22717]='h000022f4;  wr_data_rom[22717]='h00000000;
    rd_cycle[22718] = 1'b1;  wr_cycle[22718] = 1'b0;  addr_rom[22718]='h000022f8;  wr_data_rom[22718]='h00000000;
    rd_cycle[22719] = 1'b1;  wr_cycle[22719] = 1'b0;  addr_rom[22719]='h000022fc;  wr_data_rom[22719]='h00000000;
    rd_cycle[22720] = 1'b1;  wr_cycle[22720] = 1'b0;  addr_rom[22720]='h00002300;  wr_data_rom[22720]='h00000000;
    rd_cycle[22721] = 1'b1;  wr_cycle[22721] = 1'b0;  addr_rom[22721]='h00002304;  wr_data_rom[22721]='h00000000;
    rd_cycle[22722] = 1'b1;  wr_cycle[22722] = 1'b0;  addr_rom[22722]='h00002308;  wr_data_rom[22722]='h00000000;
    rd_cycle[22723] = 1'b1;  wr_cycle[22723] = 1'b0;  addr_rom[22723]='h0000230c;  wr_data_rom[22723]='h00000000;
    rd_cycle[22724] = 1'b1;  wr_cycle[22724] = 1'b0;  addr_rom[22724]='h00002310;  wr_data_rom[22724]='h00000000;
    rd_cycle[22725] = 1'b1;  wr_cycle[22725] = 1'b0;  addr_rom[22725]='h00002314;  wr_data_rom[22725]='h00000000;
    rd_cycle[22726] = 1'b1;  wr_cycle[22726] = 1'b0;  addr_rom[22726]='h00002318;  wr_data_rom[22726]='h00000000;
    rd_cycle[22727] = 1'b1;  wr_cycle[22727] = 1'b0;  addr_rom[22727]='h0000231c;  wr_data_rom[22727]='h00000000;
    rd_cycle[22728] = 1'b1;  wr_cycle[22728] = 1'b0;  addr_rom[22728]='h00002320;  wr_data_rom[22728]='h00000000;
    rd_cycle[22729] = 1'b1;  wr_cycle[22729] = 1'b0;  addr_rom[22729]='h00002324;  wr_data_rom[22729]='h00000000;
    rd_cycle[22730] = 1'b1;  wr_cycle[22730] = 1'b0;  addr_rom[22730]='h00002328;  wr_data_rom[22730]='h00000000;
    rd_cycle[22731] = 1'b1;  wr_cycle[22731] = 1'b0;  addr_rom[22731]='h0000232c;  wr_data_rom[22731]='h00000000;
    rd_cycle[22732] = 1'b1;  wr_cycle[22732] = 1'b0;  addr_rom[22732]='h00002330;  wr_data_rom[22732]='h00000000;
    rd_cycle[22733] = 1'b1;  wr_cycle[22733] = 1'b0;  addr_rom[22733]='h00002334;  wr_data_rom[22733]='h00000000;
    rd_cycle[22734] = 1'b1;  wr_cycle[22734] = 1'b0;  addr_rom[22734]='h00002338;  wr_data_rom[22734]='h00000000;
    rd_cycle[22735] = 1'b1;  wr_cycle[22735] = 1'b0;  addr_rom[22735]='h0000233c;  wr_data_rom[22735]='h00000000;
    rd_cycle[22736] = 1'b1;  wr_cycle[22736] = 1'b0;  addr_rom[22736]='h00002340;  wr_data_rom[22736]='h00000000;
    rd_cycle[22737] = 1'b1;  wr_cycle[22737] = 1'b0;  addr_rom[22737]='h00002344;  wr_data_rom[22737]='h00000000;
    rd_cycle[22738] = 1'b1;  wr_cycle[22738] = 1'b0;  addr_rom[22738]='h00002348;  wr_data_rom[22738]='h00000000;
    rd_cycle[22739] = 1'b1;  wr_cycle[22739] = 1'b0;  addr_rom[22739]='h0000234c;  wr_data_rom[22739]='h00000000;
    rd_cycle[22740] = 1'b1;  wr_cycle[22740] = 1'b0;  addr_rom[22740]='h00002350;  wr_data_rom[22740]='h00000000;
    rd_cycle[22741] = 1'b1;  wr_cycle[22741] = 1'b0;  addr_rom[22741]='h00002354;  wr_data_rom[22741]='h00000000;
    rd_cycle[22742] = 1'b1;  wr_cycle[22742] = 1'b0;  addr_rom[22742]='h00002358;  wr_data_rom[22742]='h00000000;
    rd_cycle[22743] = 1'b1;  wr_cycle[22743] = 1'b0;  addr_rom[22743]='h0000235c;  wr_data_rom[22743]='h00000000;
    rd_cycle[22744] = 1'b1;  wr_cycle[22744] = 1'b0;  addr_rom[22744]='h00002360;  wr_data_rom[22744]='h00000000;
    rd_cycle[22745] = 1'b1;  wr_cycle[22745] = 1'b0;  addr_rom[22745]='h00002364;  wr_data_rom[22745]='h00000000;
    rd_cycle[22746] = 1'b1;  wr_cycle[22746] = 1'b0;  addr_rom[22746]='h00002368;  wr_data_rom[22746]='h00000000;
    rd_cycle[22747] = 1'b1;  wr_cycle[22747] = 1'b0;  addr_rom[22747]='h0000236c;  wr_data_rom[22747]='h00000000;
    rd_cycle[22748] = 1'b1;  wr_cycle[22748] = 1'b0;  addr_rom[22748]='h00002370;  wr_data_rom[22748]='h00000000;
    rd_cycle[22749] = 1'b1;  wr_cycle[22749] = 1'b0;  addr_rom[22749]='h00002374;  wr_data_rom[22749]='h00000000;
    rd_cycle[22750] = 1'b1;  wr_cycle[22750] = 1'b0;  addr_rom[22750]='h00002378;  wr_data_rom[22750]='h00000000;
    rd_cycle[22751] = 1'b1;  wr_cycle[22751] = 1'b0;  addr_rom[22751]='h0000237c;  wr_data_rom[22751]='h00000000;
    rd_cycle[22752] = 1'b1;  wr_cycle[22752] = 1'b0;  addr_rom[22752]='h00002380;  wr_data_rom[22752]='h00000000;
    rd_cycle[22753] = 1'b1;  wr_cycle[22753] = 1'b0;  addr_rom[22753]='h00002384;  wr_data_rom[22753]='h00000000;
    rd_cycle[22754] = 1'b1;  wr_cycle[22754] = 1'b0;  addr_rom[22754]='h00002388;  wr_data_rom[22754]='h00000000;
    rd_cycle[22755] = 1'b1;  wr_cycle[22755] = 1'b0;  addr_rom[22755]='h0000238c;  wr_data_rom[22755]='h00000000;
    rd_cycle[22756] = 1'b1;  wr_cycle[22756] = 1'b0;  addr_rom[22756]='h00002390;  wr_data_rom[22756]='h00000000;
    rd_cycle[22757] = 1'b1;  wr_cycle[22757] = 1'b0;  addr_rom[22757]='h00002394;  wr_data_rom[22757]='h00000000;
    rd_cycle[22758] = 1'b1;  wr_cycle[22758] = 1'b0;  addr_rom[22758]='h00002398;  wr_data_rom[22758]='h00000000;
    rd_cycle[22759] = 1'b1;  wr_cycle[22759] = 1'b0;  addr_rom[22759]='h0000239c;  wr_data_rom[22759]='h00000000;
    rd_cycle[22760] = 1'b1;  wr_cycle[22760] = 1'b0;  addr_rom[22760]='h000023a0;  wr_data_rom[22760]='h00000000;
    rd_cycle[22761] = 1'b1;  wr_cycle[22761] = 1'b0;  addr_rom[22761]='h000023a4;  wr_data_rom[22761]='h00000000;
    rd_cycle[22762] = 1'b1;  wr_cycle[22762] = 1'b0;  addr_rom[22762]='h000023a8;  wr_data_rom[22762]='h00000000;
    rd_cycle[22763] = 1'b1;  wr_cycle[22763] = 1'b0;  addr_rom[22763]='h000023ac;  wr_data_rom[22763]='h00000000;
    rd_cycle[22764] = 1'b1;  wr_cycle[22764] = 1'b0;  addr_rom[22764]='h000023b0;  wr_data_rom[22764]='h00000000;
    rd_cycle[22765] = 1'b1;  wr_cycle[22765] = 1'b0;  addr_rom[22765]='h000023b4;  wr_data_rom[22765]='h00000000;
    rd_cycle[22766] = 1'b1;  wr_cycle[22766] = 1'b0;  addr_rom[22766]='h000023b8;  wr_data_rom[22766]='h00000000;
    rd_cycle[22767] = 1'b1;  wr_cycle[22767] = 1'b0;  addr_rom[22767]='h000023bc;  wr_data_rom[22767]='h00000000;
    rd_cycle[22768] = 1'b1;  wr_cycle[22768] = 1'b0;  addr_rom[22768]='h000023c0;  wr_data_rom[22768]='h00000000;
    rd_cycle[22769] = 1'b1;  wr_cycle[22769] = 1'b0;  addr_rom[22769]='h000023c4;  wr_data_rom[22769]='h00000000;
    rd_cycle[22770] = 1'b1;  wr_cycle[22770] = 1'b0;  addr_rom[22770]='h000023c8;  wr_data_rom[22770]='h00000000;
    rd_cycle[22771] = 1'b1;  wr_cycle[22771] = 1'b0;  addr_rom[22771]='h000023cc;  wr_data_rom[22771]='h00000000;
    rd_cycle[22772] = 1'b1;  wr_cycle[22772] = 1'b0;  addr_rom[22772]='h000023d0;  wr_data_rom[22772]='h00000000;
    rd_cycle[22773] = 1'b1;  wr_cycle[22773] = 1'b0;  addr_rom[22773]='h000023d4;  wr_data_rom[22773]='h00000000;
    rd_cycle[22774] = 1'b1;  wr_cycle[22774] = 1'b0;  addr_rom[22774]='h000023d8;  wr_data_rom[22774]='h00000000;
    rd_cycle[22775] = 1'b1;  wr_cycle[22775] = 1'b0;  addr_rom[22775]='h000023dc;  wr_data_rom[22775]='h00000000;
    rd_cycle[22776] = 1'b1;  wr_cycle[22776] = 1'b0;  addr_rom[22776]='h000023e0;  wr_data_rom[22776]='h00000000;
    rd_cycle[22777] = 1'b1;  wr_cycle[22777] = 1'b0;  addr_rom[22777]='h000023e4;  wr_data_rom[22777]='h00000000;
    rd_cycle[22778] = 1'b1;  wr_cycle[22778] = 1'b0;  addr_rom[22778]='h000023e8;  wr_data_rom[22778]='h00000000;
    rd_cycle[22779] = 1'b1;  wr_cycle[22779] = 1'b0;  addr_rom[22779]='h000023ec;  wr_data_rom[22779]='h00000000;
    rd_cycle[22780] = 1'b1;  wr_cycle[22780] = 1'b0;  addr_rom[22780]='h000023f0;  wr_data_rom[22780]='h00000000;
    rd_cycle[22781] = 1'b1;  wr_cycle[22781] = 1'b0;  addr_rom[22781]='h000023f4;  wr_data_rom[22781]='h00000000;
    rd_cycle[22782] = 1'b1;  wr_cycle[22782] = 1'b0;  addr_rom[22782]='h000023f8;  wr_data_rom[22782]='h00000000;
    rd_cycle[22783] = 1'b1;  wr_cycle[22783] = 1'b0;  addr_rom[22783]='h000023fc;  wr_data_rom[22783]='h00000000;
    rd_cycle[22784] = 1'b1;  wr_cycle[22784] = 1'b0;  addr_rom[22784]='h00002400;  wr_data_rom[22784]='h00000000;
    rd_cycle[22785] = 1'b1;  wr_cycle[22785] = 1'b0;  addr_rom[22785]='h00002404;  wr_data_rom[22785]='h00000000;
    rd_cycle[22786] = 1'b1;  wr_cycle[22786] = 1'b0;  addr_rom[22786]='h00002408;  wr_data_rom[22786]='h00000000;
    rd_cycle[22787] = 1'b1;  wr_cycle[22787] = 1'b0;  addr_rom[22787]='h0000240c;  wr_data_rom[22787]='h00000000;
    rd_cycle[22788] = 1'b1;  wr_cycle[22788] = 1'b0;  addr_rom[22788]='h00002410;  wr_data_rom[22788]='h00000000;
    rd_cycle[22789] = 1'b1;  wr_cycle[22789] = 1'b0;  addr_rom[22789]='h00002414;  wr_data_rom[22789]='h00000000;
    rd_cycle[22790] = 1'b1;  wr_cycle[22790] = 1'b0;  addr_rom[22790]='h00002418;  wr_data_rom[22790]='h00000000;
    rd_cycle[22791] = 1'b1;  wr_cycle[22791] = 1'b0;  addr_rom[22791]='h0000241c;  wr_data_rom[22791]='h00000000;
    rd_cycle[22792] = 1'b1;  wr_cycle[22792] = 1'b0;  addr_rom[22792]='h00002420;  wr_data_rom[22792]='h00000000;
    rd_cycle[22793] = 1'b1;  wr_cycle[22793] = 1'b0;  addr_rom[22793]='h00002424;  wr_data_rom[22793]='h00000000;
    rd_cycle[22794] = 1'b1;  wr_cycle[22794] = 1'b0;  addr_rom[22794]='h00002428;  wr_data_rom[22794]='h00000000;
    rd_cycle[22795] = 1'b1;  wr_cycle[22795] = 1'b0;  addr_rom[22795]='h0000242c;  wr_data_rom[22795]='h00000000;
    rd_cycle[22796] = 1'b1;  wr_cycle[22796] = 1'b0;  addr_rom[22796]='h00002430;  wr_data_rom[22796]='h00000000;
    rd_cycle[22797] = 1'b1;  wr_cycle[22797] = 1'b0;  addr_rom[22797]='h00002434;  wr_data_rom[22797]='h00000000;
    rd_cycle[22798] = 1'b1;  wr_cycle[22798] = 1'b0;  addr_rom[22798]='h00002438;  wr_data_rom[22798]='h00000000;
    rd_cycle[22799] = 1'b1;  wr_cycle[22799] = 1'b0;  addr_rom[22799]='h0000243c;  wr_data_rom[22799]='h00000000;
    rd_cycle[22800] = 1'b1;  wr_cycle[22800] = 1'b0;  addr_rom[22800]='h00002440;  wr_data_rom[22800]='h00000000;
    rd_cycle[22801] = 1'b1;  wr_cycle[22801] = 1'b0;  addr_rom[22801]='h00002444;  wr_data_rom[22801]='h00000000;
    rd_cycle[22802] = 1'b1;  wr_cycle[22802] = 1'b0;  addr_rom[22802]='h00002448;  wr_data_rom[22802]='h00000000;
    rd_cycle[22803] = 1'b1;  wr_cycle[22803] = 1'b0;  addr_rom[22803]='h0000244c;  wr_data_rom[22803]='h00000000;
    rd_cycle[22804] = 1'b1;  wr_cycle[22804] = 1'b0;  addr_rom[22804]='h00002450;  wr_data_rom[22804]='h00000000;
    rd_cycle[22805] = 1'b1;  wr_cycle[22805] = 1'b0;  addr_rom[22805]='h00002454;  wr_data_rom[22805]='h00000000;
    rd_cycle[22806] = 1'b1;  wr_cycle[22806] = 1'b0;  addr_rom[22806]='h00002458;  wr_data_rom[22806]='h00000000;
    rd_cycle[22807] = 1'b1;  wr_cycle[22807] = 1'b0;  addr_rom[22807]='h0000245c;  wr_data_rom[22807]='h00000000;
    rd_cycle[22808] = 1'b1;  wr_cycle[22808] = 1'b0;  addr_rom[22808]='h00002460;  wr_data_rom[22808]='h00000000;
    rd_cycle[22809] = 1'b1;  wr_cycle[22809] = 1'b0;  addr_rom[22809]='h00002464;  wr_data_rom[22809]='h00000000;
    rd_cycle[22810] = 1'b1;  wr_cycle[22810] = 1'b0;  addr_rom[22810]='h00002468;  wr_data_rom[22810]='h00000000;
    rd_cycle[22811] = 1'b1;  wr_cycle[22811] = 1'b0;  addr_rom[22811]='h0000246c;  wr_data_rom[22811]='h00000000;
    rd_cycle[22812] = 1'b1;  wr_cycle[22812] = 1'b0;  addr_rom[22812]='h00002470;  wr_data_rom[22812]='h00000000;
    rd_cycle[22813] = 1'b1;  wr_cycle[22813] = 1'b0;  addr_rom[22813]='h00002474;  wr_data_rom[22813]='h00000000;
    rd_cycle[22814] = 1'b1;  wr_cycle[22814] = 1'b0;  addr_rom[22814]='h00002478;  wr_data_rom[22814]='h00000000;
    rd_cycle[22815] = 1'b1;  wr_cycle[22815] = 1'b0;  addr_rom[22815]='h0000247c;  wr_data_rom[22815]='h00000000;
    rd_cycle[22816] = 1'b1;  wr_cycle[22816] = 1'b0;  addr_rom[22816]='h00002480;  wr_data_rom[22816]='h00000000;
    rd_cycle[22817] = 1'b1;  wr_cycle[22817] = 1'b0;  addr_rom[22817]='h00002484;  wr_data_rom[22817]='h00000000;
    rd_cycle[22818] = 1'b1;  wr_cycle[22818] = 1'b0;  addr_rom[22818]='h00002488;  wr_data_rom[22818]='h00000000;
    rd_cycle[22819] = 1'b1;  wr_cycle[22819] = 1'b0;  addr_rom[22819]='h0000248c;  wr_data_rom[22819]='h00000000;
    rd_cycle[22820] = 1'b1;  wr_cycle[22820] = 1'b0;  addr_rom[22820]='h00002490;  wr_data_rom[22820]='h00000000;
    rd_cycle[22821] = 1'b1;  wr_cycle[22821] = 1'b0;  addr_rom[22821]='h00002494;  wr_data_rom[22821]='h00000000;
    rd_cycle[22822] = 1'b1;  wr_cycle[22822] = 1'b0;  addr_rom[22822]='h00002498;  wr_data_rom[22822]='h00000000;
    rd_cycle[22823] = 1'b1;  wr_cycle[22823] = 1'b0;  addr_rom[22823]='h0000249c;  wr_data_rom[22823]='h00000000;
    rd_cycle[22824] = 1'b1;  wr_cycle[22824] = 1'b0;  addr_rom[22824]='h000024a0;  wr_data_rom[22824]='h00000000;
    rd_cycle[22825] = 1'b1;  wr_cycle[22825] = 1'b0;  addr_rom[22825]='h000024a4;  wr_data_rom[22825]='h00000000;
    rd_cycle[22826] = 1'b1;  wr_cycle[22826] = 1'b0;  addr_rom[22826]='h000024a8;  wr_data_rom[22826]='h00000000;
    rd_cycle[22827] = 1'b1;  wr_cycle[22827] = 1'b0;  addr_rom[22827]='h000024ac;  wr_data_rom[22827]='h00000000;
    rd_cycle[22828] = 1'b1;  wr_cycle[22828] = 1'b0;  addr_rom[22828]='h000024b0;  wr_data_rom[22828]='h00000000;
    rd_cycle[22829] = 1'b1;  wr_cycle[22829] = 1'b0;  addr_rom[22829]='h000024b4;  wr_data_rom[22829]='h00000000;
    rd_cycle[22830] = 1'b1;  wr_cycle[22830] = 1'b0;  addr_rom[22830]='h000024b8;  wr_data_rom[22830]='h00000000;
    rd_cycle[22831] = 1'b1;  wr_cycle[22831] = 1'b0;  addr_rom[22831]='h000024bc;  wr_data_rom[22831]='h00000000;
    rd_cycle[22832] = 1'b1;  wr_cycle[22832] = 1'b0;  addr_rom[22832]='h000024c0;  wr_data_rom[22832]='h00000000;
    rd_cycle[22833] = 1'b1;  wr_cycle[22833] = 1'b0;  addr_rom[22833]='h000024c4;  wr_data_rom[22833]='h00000000;
    rd_cycle[22834] = 1'b1;  wr_cycle[22834] = 1'b0;  addr_rom[22834]='h000024c8;  wr_data_rom[22834]='h00000000;
    rd_cycle[22835] = 1'b1;  wr_cycle[22835] = 1'b0;  addr_rom[22835]='h000024cc;  wr_data_rom[22835]='h00000000;
    rd_cycle[22836] = 1'b1;  wr_cycle[22836] = 1'b0;  addr_rom[22836]='h000024d0;  wr_data_rom[22836]='h00000000;
    rd_cycle[22837] = 1'b1;  wr_cycle[22837] = 1'b0;  addr_rom[22837]='h000024d4;  wr_data_rom[22837]='h00000000;
    rd_cycle[22838] = 1'b1;  wr_cycle[22838] = 1'b0;  addr_rom[22838]='h000024d8;  wr_data_rom[22838]='h00000000;
    rd_cycle[22839] = 1'b1;  wr_cycle[22839] = 1'b0;  addr_rom[22839]='h000024dc;  wr_data_rom[22839]='h00000000;
    rd_cycle[22840] = 1'b1;  wr_cycle[22840] = 1'b0;  addr_rom[22840]='h000024e0;  wr_data_rom[22840]='h00000000;
    rd_cycle[22841] = 1'b1;  wr_cycle[22841] = 1'b0;  addr_rom[22841]='h000024e4;  wr_data_rom[22841]='h00000000;
    rd_cycle[22842] = 1'b1;  wr_cycle[22842] = 1'b0;  addr_rom[22842]='h000024e8;  wr_data_rom[22842]='h00000000;
    rd_cycle[22843] = 1'b1;  wr_cycle[22843] = 1'b0;  addr_rom[22843]='h000024ec;  wr_data_rom[22843]='h00000000;
    rd_cycle[22844] = 1'b1;  wr_cycle[22844] = 1'b0;  addr_rom[22844]='h000024f0;  wr_data_rom[22844]='h00000000;
    rd_cycle[22845] = 1'b1;  wr_cycle[22845] = 1'b0;  addr_rom[22845]='h000024f4;  wr_data_rom[22845]='h00000000;
    rd_cycle[22846] = 1'b1;  wr_cycle[22846] = 1'b0;  addr_rom[22846]='h000024f8;  wr_data_rom[22846]='h00000000;
    rd_cycle[22847] = 1'b1;  wr_cycle[22847] = 1'b0;  addr_rom[22847]='h000024fc;  wr_data_rom[22847]='h00000000;
    rd_cycle[22848] = 1'b1;  wr_cycle[22848] = 1'b0;  addr_rom[22848]='h00002500;  wr_data_rom[22848]='h00000000;
    rd_cycle[22849] = 1'b1;  wr_cycle[22849] = 1'b0;  addr_rom[22849]='h00002504;  wr_data_rom[22849]='h00000000;
    rd_cycle[22850] = 1'b1;  wr_cycle[22850] = 1'b0;  addr_rom[22850]='h00002508;  wr_data_rom[22850]='h00000000;
    rd_cycle[22851] = 1'b1;  wr_cycle[22851] = 1'b0;  addr_rom[22851]='h0000250c;  wr_data_rom[22851]='h00000000;
    rd_cycle[22852] = 1'b1;  wr_cycle[22852] = 1'b0;  addr_rom[22852]='h00002510;  wr_data_rom[22852]='h00000000;
    rd_cycle[22853] = 1'b1;  wr_cycle[22853] = 1'b0;  addr_rom[22853]='h00002514;  wr_data_rom[22853]='h00000000;
    rd_cycle[22854] = 1'b1;  wr_cycle[22854] = 1'b0;  addr_rom[22854]='h00002518;  wr_data_rom[22854]='h00000000;
    rd_cycle[22855] = 1'b1;  wr_cycle[22855] = 1'b0;  addr_rom[22855]='h0000251c;  wr_data_rom[22855]='h00000000;
    rd_cycle[22856] = 1'b1;  wr_cycle[22856] = 1'b0;  addr_rom[22856]='h00002520;  wr_data_rom[22856]='h00000000;
    rd_cycle[22857] = 1'b1;  wr_cycle[22857] = 1'b0;  addr_rom[22857]='h00002524;  wr_data_rom[22857]='h00000000;
    rd_cycle[22858] = 1'b1;  wr_cycle[22858] = 1'b0;  addr_rom[22858]='h00002528;  wr_data_rom[22858]='h00000000;
    rd_cycle[22859] = 1'b1;  wr_cycle[22859] = 1'b0;  addr_rom[22859]='h0000252c;  wr_data_rom[22859]='h00000000;
    rd_cycle[22860] = 1'b1;  wr_cycle[22860] = 1'b0;  addr_rom[22860]='h00002530;  wr_data_rom[22860]='h00000000;
    rd_cycle[22861] = 1'b1;  wr_cycle[22861] = 1'b0;  addr_rom[22861]='h00002534;  wr_data_rom[22861]='h00000000;
    rd_cycle[22862] = 1'b1;  wr_cycle[22862] = 1'b0;  addr_rom[22862]='h00002538;  wr_data_rom[22862]='h00000000;
    rd_cycle[22863] = 1'b1;  wr_cycle[22863] = 1'b0;  addr_rom[22863]='h0000253c;  wr_data_rom[22863]='h00000000;
    rd_cycle[22864] = 1'b1;  wr_cycle[22864] = 1'b0;  addr_rom[22864]='h00002540;  wr_data_rom[22864]='h00000000;
    rd_cycle[22865] = 1'b1;  wr_cycle[22865] = 1'b0;  addr_rom[22865]='h00002544;  wr_data_rom[22865]='h00000000;
    rd_cycle[22866] = 1'b1;  wr_cycle[22866] = 1'b0;  addr_rom[22866]='h00002548;  wr_data_rom[22866]='h00000000;
    rd_cycle[22867] = 1'b1;  wr_cycle[22867] = 1'b0;  addr_rom[22867]='h0000254c;  wr_data_rom[22867]='h00000000;
    rd_cycle[22868] = 1'b1;  wr_cycle[22868] = 1'b0;  addr_rom[22868]='h00002550;  wr_data_rom[22868]='h00000000;
    rd_cycle[22869] = 1'b1;  wr_cycle[22869] = 1'b0;  addr_rom[22869]='h00002554;  wr_data_rom[22869]='h00000000;
    rd_cycle[22870] = 1'b1;  wr_cycle[22870] = 1'b0;  addr_rom[22870]='h00002558;  wr_data_rom[22870]='h00000000;
    rd_cycle[22871] = 1'b1;  wr_cycle[22871] = 1'b0;  addr_rom[22871]='h0000255c;  wr_data_rom[22871]='h00000000;
    rd_cycle[22872] = 1'b1;  wr_cycle[22872] = 1'b0;  addr_rom[22872]='h00002560;  wr_data_rom[22872]='h00000000;
    rd_cycle[22873] = 1'b1;  wr_cycle[22873] = 1'b0;  addr_rom[22873]='h00002564;  wr_data_rom[22873]='h00000000;
    rd_cycle[22874] = 1'b1;  wr_cycle[22874] = 1'b0;  addr_rom[22874]='h00002568;  wr_data_rom[22874]='h00000000;
    rd_cycle[22875] = 1'b1;  wr_cycle[22875] = 1'b0;  addr_rom[22875]='h0000256c;  wr_data_rom[22875]='h00000000;
    rd_cycle[22876] = 1'b1;  wr_cycle[22876] = 1'b0;  addr_rom[22876]='h00002570;  wr_data_rom[22876]='h00000000;
    rd_cycle[22877] = 1'b1;  wr_cycle[22877] = 1'b0;  addr_rom[22877]='h00002574;  wr_data_rom[22877]='h00000000;
    rd_cycle[22878] = 1'b1;  wr_cycle[22878] = 1'b0;  addr_rom[22878]='h00002578;  wr_data_rom[22878]='h00000000;
    rd_cycle[22879] = 1'b1;  wr_cycle[22879] = 1'b0;  addr_rom[22879]='h0000257c;  wr_data_rom[22879]='h00000000;
    rd_cycle[22880] = 1'b1;  wr_cycle[22880] = 1'b0;  addr_rom[22880]='h00002580;  wr_data_rom[22880]='h00000000;
    rd_cycle[22881] = 1'b1;  wr_cycle[22881] = 1'b0;  addr_rom[22881]='h00002584;  wr_data_rom[22881]='h00000000;
    rd_cycle[22882] = 1'b1;  wr_cycle[22882] = 1'b0;  addr_rom[22882]='h00002588;  wr_data_rom[22882]='h00000000;
    rd_cycle[22883] = 1'b1;  wr_cycle[22883] = 1'b0;  addr_rom[22883]='h0000258c;  wr_data_rom[22883]='h00000000;
    rd_cycle[22884] = 1'b1;  wr_cycle[22884] = 1'b0;  addr_rom[22884]='h00002590;  wr_data_rom[22884]='h00000000;
    rd_cycle[22885] = 1'b1;  wr_cycle[22885] = 1'b0;  addr_rom[22885]='h00002594;  wr_data_rom[22885]='h00000000;
    rd_cycle[22886] = 1'b1;  wr_cycle[22886] = 1'b0;  addr_rom[22886]='h00002598;  wr_data_rom[22886]='h00000000;
    rd_cycle[22887] = 1'b1;  wr_cycle[22887] = 1'b0;  addr_rom[22887]='h0000259c;  wr_data_rom[22887]='h00000000;
    rd_cycle[22888] = 1'b1;  wr_cycle[22888] = 1'b0;  addr_rom[22888]='h000025a0;  wr_data_rom[22888]='h00000000;
    rd_cycle[22889] = 1'b1;  wr_cycle[22889] = 1'b0;  addr_rom[22889]='h000025a4;  wr_data_rom[22889]='h00000000;
    rd_cycle[22890] = 1'b1;  wr_cycle[22890] = 1'b0;  addr_rom[22890]='h000025a8;  wr_data_rom[22890]='h00000000;
    rd_cycle[22891] = 1'b1;  wr_cycle[22891] = 1'b0;  addr_rom[22891]='h000025ac;  wr_data_rom[22891]='h00000000;
    rd_cycle[22892] = 1'b1;  wr_cycle[22892] = 1'b0;  addr_rom[22892]='h000025b0;  wr_data_rom[22892]='h00000000;
    rd_cycle[22893] = 1'b1;  wr_cycle[22893] = 1'b0;  addr_rom[22893]='h000025b4;  wr_data_rom[22893]='h00000000;
    rd_cycle[22894] = 1'b1;  wr_cycle[22894] = 1'b0;  addr_rom[22894]='h000025b8;  wr_data_rom[22894]='h00000000;
    rd_cycle[22895] = 1'b1;  wr_cycle[22895] = 1'b0;  addr_rom[22895]='h000025bc;  wr_data_rom[22895]='h00000000;
    rd_cycle[22896] = 1'b1;  wr_cycle[22896] = 1'b0;  addr_rom[22896]='h000025c0;  wr_data_rom[22896]='h00000000;
    rd_cycle[22897] = 1'b1;  wr_cycle[22897] = 1'b0;  addr_rom[22897]='h000025c4;  wr_data_rom[22897]='h00000000;
    rd_cycle[22898] = 1'b1;  wr_cycle[22898] = 1'b0;  addr_rom[22898]='h000025c8;  wr_data_rom[22898]='h00000000;
    rd_cycle[22899] = 1'b1;  wr_cycle[22899] = 1'b0;  addr_rom[22899]='h000025cc;  wr_data_rom[22899]='h00000000;
    rd_cycle[22900] = 1'b1;  wr_cycle[22900] = 1'b0;  addr_rom[22900]='h000025d0;  wr_data_rom[22900]='h00000000;
    rd_cycle[22901] = 1'b1;  wr_cycle[22901] = 1'b0;  addr_rom[22901]='h000025d4;  wr_data_rom[22901]='h00000000;
    rd_cycle[22902] = 1'b1;  wr_cycle[22902] = 1'b0;  addr_rom[22902]='h000025d8;  wr_data_rom[22902]='h00000000;
    rd_cycle[22903] = 1'b1;  wr_cycle[22903] = 1'b0;  addr_rom[22903]='h000025dc;  wr_data_rom[22903]='h00000000;
    rd_cycle[22904] = 1'b1;  wr_cycle[22904] = 1'b0;  addr_rom[22904]='h000025e0;  wr_data_rom[22904]='h00000000;
    rd_cycle[22905] = 1'b1;  wr_cycle[22905] = 1'b0;  addr_rom[22905]='h000025e4;  wr_data_rom[22905]='h00000000;
    rd_cycle[22906] = 1'b1;  wr_cycle[22906] = 1'b0;  addr_rom[22906]='h000025e8;  wr_data_rom[22906]='h00000000;
    rd_cycle[22907] = 1'b1;  wr_cycle[22907] = 1'b0;  addr_rom[22907]='h000025ec;  wr_data_rom[22907]='h00000000;
    rd_cycle[22908] = 1'b1;  wr_cycle[22908] = 1'b0;  addr_rom[22908]='h000025f0;  wr_data_rom[22908]='h00000000;
    rd_cycle[22909] = 1'b1;  wr_cycle[22909] = 1'b0;  addr_rom[22909]='h000025f4;  wr_data_rom[22909]='h00000000;
    rd_cycle[22910] = 1'b1;  wr_cycle[22910] = 1'b0;  addr_rom[22910]='h000025f8;  wr_data_rom[22910]='h00000000;
    rd_cycle[22911] = 1'b1;  wr_cycle[22911] = 1'b0;  addr_rom[22911]='h000025fc;  wr_data_rom[22911]='h00000000;
    rd_cycle[22912] = 1'b1;  wr_cycle[22912] = 1'b0;  addr_rom[22912]='h00002600;  wr_data_rom[22912]='h00000000;
    rd_cycle[22913] = 1'b1;  wr_cycle[22913] = 1'b0;  addr_rom[22913]='h00002604;  wr_data_rom[22913]='h00000000;
    rd_cycle[22914] = 1'b1;  wr_cycle[22914] = 1'b0;  addr_rom[22914]='h00002608;  wr_data_rom[22914]='h00000000;
    rd_cycle[22915] = 1'b1;  wr_cycle[22915] = 1'b0;  addr_rom[22915]='h0000260c;  wr_data_rom[22915]='h00000000;
    rd_cycle[22916] = 1'b1;  wr_cycle[22916] = 1'b0;  addr_rom[22916]='h00002610;  wr_data_rom[22916]='h00000000;
    rd_cycle[22917] = 1'b1;  wr_cycle[22917] = 1'b0;  addr_rom[22917]='h00002614;  wr_data_rom[22917]='h00000000;
    rd_cycle[22918] = 1'b1;  wr_cycle[22918] = 1'b0;  addr_rom[22918]='h00002618;  wr_data_rom[22918]='h00000000;
    rd_cycle[22919] = 1'b1;  wr_cycle[22919] = 1'b0;  addr_rom[22919]='h0000261c;  wr_data_rom[22919]='h00000000;
    rd_cycle[22920] = 1'b1;  wr_cycle[22920] = 1'b0;  addr_rom[22920]='h00002620;  wr_data_rom[22920]='h00000000;
    rd_cycle[22921] = 1'b1;  wr_cycle[22921] = 1'b0;  addr_rom[22921]='h00002624;  wr_data_rom[22921]='h00000000;
    rd_cycle[22922] = 1'b1;  wr_cycle[22922] = 1'b0;  addr_rom[22922]='h00002628;  wr_data_rom[22922]='h00000000;
    rd_cycle[22923] = 1'b1;  wr_cycle[22923] = 1'b0;  addr_rom[22923]='h0000262c;  wr_data_rom[22923]='h00000000;
    rd_cycle[22924] = 1'b1;  wr_cycle[22924] = 1'b0;  addr_rom[22924]='h00002630;  wr_data_rom[22924]='h00000000;
    rd_cycle[22925] = 1'b1;  wr_cycle[22925] = 1'b0;  addr_rom[22925]='h00002634;  wr_data_rom[22925]='h00000000;
    rd_cycle[22926] = 1'b1;  wr_cycle[22926] = 1'b0;  addr_rom[22926]='h00002638;  wr_data_rom[22926]='h00000000;
    rd_cycle[22927] = 1'b1;  wr_cycle[22927] = 1'b0;  addr_rom[22927]='h0000263c;  wr_data_rom[22927]='h00000000;
    rd_cycle[22928] = 1'b1;  wr_cycle[22928] = 1'b0;  addr_rom[22928]='h00002640;  wr_data_rom[22928]='h00000000;
    rd_cycle[22929] = 1'b1;  wr_cycle[22929] = 1'b0;  addr_rom[22929]='h00002644;  wr_data_rom[22929]='h00000000;
    rd_cycle[22930] = 1'b1;  wr_cycle[22930] = 1'b0;  addr_rom[22930]='h00002648;  wr_data_rom[22930]='h00000000;
    rd_cycle[22931] = 1'b1;  wr_cycle[22931] = 1'b0;  addr_rom[22931]='h0000264c;  wr_data_rom[22931]='h00000000;
    rd_cycle[22932] = 1'b1;  wr_cycle[22932] = 1'b0;  addr_rom[22932]='h00002650;  wr_data_rom[22932]='h00000000;
    rd_cycle[22933] = 1'b1;  wr_cycle[22933] = 1'b0;  addr_rom[22933]='h00002654;  wr_data_rom[22933]='h00000000;
    rd_cycle[22934] = 1'b1;  wr_cycle[22934] = 1'b0;  addr_rom[22934]='h00002658;  wr_data_rom[22934]='h00000000;
    rd_cycle[22935] = 1'b1;  wr_cycle[22935] = 1'b0;  addr_rom[22935]='h0000265c;  wr_data_rom[22935]='h00000000;
    rd_cycle[22936] = 1'b1;  wr_cycle[22936] = 1'b0;  addr_rom[22936]='h00002660;  wr_data_rom[22936]='h00000000;
    rd_cycle[22937] = 1'b1;  wr_cycle[22937] = 1'b0;  addr_rom[22937]='h00002664;  wr_data_rom[22937]='h00000000;
    rd_cycle[22938] = 1'b1;  wr_cycle[22938] = 1'b0;  addr_rom[22938]='h00002668;  wr_data_rom[22938]='h00000000;
    rd_cycle[22939] = 1'b1;  wr_cycle[22939] = 1'b0;  addr_rom[22939]='h0000266c;  wr_data_rom[22939]='h00000000;
    rd_cycle[22940] = 1'b1;  wr_cycle[22940] = 1'b0;  addr_rom[22940]='h00002670;  wr_data_rom[22940]='h00000000;
    rd_cycle[22941] = 1'b1;  wr_cycle[22941] = 1'b0;  addr_rom[22941]='h00002674;  wr_data_rom[22941]='h00000000;
    rd_cycle[22942] = 1'b1;  wr_cycle[22942] = 1'b0;  addr_rom[22942]='h00002678;  wr_data_rom[22942]='h00000000;
    rd_cycle[22943] = 1'b1;  wr_cycle[22943] = 1'b0;  addr_rom[22943]='h0000267c;  wr_data_rom[22943]='h00000000;
    rd_cycle[22944] = 1'b1;  wr_cycle[22944] = 1'b0;  addr_rom[22944]='h00002680;  wr_data_rom[22944]='h00000000;
    rd_cycle[22945] = 1'b1;  wr_cycle[22945] = 1'b0;  addr_rom[22945]='h00002684;  wr_data_rom[22945]='h00000000;
    rd_cycle[22946] = 1'b1;  wr_cycle[22946] = 1'b0;  addr_rom[22946]='h00002688;  wr_data_rom[22946]='h00000000;
    rd_cycle[22947] = 1'b1;  wr_cycle[22947] = 1'b0;  addr_rom[22947]='h0000268c;  wr_data_rom[22947]='h00000000;
    rd_cycle[22948] = 1'b1;  wr_cycle[22948] = 1'b0;  addr_rom[22948]='h00002690;  wr_data_rom[22948]='h00000000;
    rd_cycle[22949] = 1'b1;  wr_cycle[22949] = 1'b0;  addr_rom[22949]='h00002694;  wr_data_rom[22949]='h00000000;
    rd_cycle[22950] = 1'b1;  wr_cycle[22950] = 1'b0;  addr_rom[22950]='h00002698;  wr_data_rom[22950]='h00000000;
    rd_cycle[22951] = 1'b1;  wr_cycle[22951] = 1'b0;  addr_rom[22951]='h0000269c;  wr_data_rom[22951]='h00000000;
    rd_cycle[22952] = 1'b1;  wr_cycle[22952] = 1'b0;  addr_rom[22952]='h000026a0;  wr_data_rom[22952]='h00000000;
    rd_cycle[22953] = 1'b1;  wr_cycle[22953] = 1'b0;  addr_rom[22953]='h000026a4;  wr_data_rom[22953]='h00000000;
    rd_cycle[22954] = 1'b1;  wr_cycle[22954] = 1'b0;  addr_rom[22954]='h000026a8;  wr_data_rom[22954]='h00000000;
    rd_cycle[22955] = 1'b1;  wr_cycle[22955] = 1'b0;  addr_rom[22955]='h000026ac;  wr_data_rom[22955]='h00000000;
    rd_cycle[22956] = 1'b1;  wr_cycle[22956] = 1'b0;  addr_rom[22956]='h000026b0;  wr_data_rom[22956]='h00000000;
    rd_cycle[22957] = 1'b1;  wr_cycle[22957] = 1'b0;  addr_rom[22957]='h000026b4;  wr_data_rom[22957]='h00000000;
    rd_cycle[22958] = 1'b1;  wr_cycle[22958] = 1'b0;  addr_rom[22958]='h000026b8;  wr_data_rom[22958]='h00000000;
    rd_cycle[22959] = 1'b1;  wr_cycle[22959] = 1'b0;  addr_rom[22959]='h000026bc;  wr_data_rom[22959]='h00000000;
    rd_cycle[22960] = 1'b1;  wr_cycle[22960] = 1'b0;  addr_rom[22960]='h000026c0;  wr_data_rom[22960]='h00000000;
    rd_cycle[22961] = 1'b1;  wr_cycle[22961] = 1'b0;  addr_rom[22961]='h000026c4;  wr_data_rom[22961]='h00000000;
    rd_cycle[22962] = 1'b1;  wr_cycle[22962] = 1'b0;  addr_rom[22962]='h000026c8;  wr_data_rom[22962]='h00000000;
    rd_cycle[22963] = 1'b1;  wr_cycle[22963] = 1'b0;  addr_rom[22963]='h000026cc;  wr_data_rom[22963]='h00000000;
    rd_cycle[22964] = 1'b1;  wr_cycle[22964] = 1'b0;  addr_rom[22964]='h000026d0;  wr_data_rom[22964]='h00000000;
    rd_cycle[22965] = 1'b1;  wr_cycle[22965] = 1'b0;  addr_rom[22965]='h000026d4;  wr_data_rom[22965]='h00000000;
    rd_cycle[22966] = 1'b1;  wr_cycle[22966] = 1'b0;  addr_rom[22966]='h000026d8;  wr_data_rom[22966]='h00000000;
    rd_cycle[22967] = 1'b1;  wr_cycle[22967] = 1'b0;  addr_rom[22967]='h000026dc;  wr_data_rom[22967]='h00000000;
    rd_cycle[22968] = 1'b1;  wr_cycle[22968] = 1'b0;  addr_rom[22968]='h000026e0;  wr_data_rom[22968]='h00000000;
    rd_cycle[22969] = 1'b1;  wr_cycle[22969] = 1'b0;  addr_rom[22969]='h000026e4;  wr_data_rom[22969]='h00000000;
    rd_cycle[22970] = 1'b1;  wr_cycle[22970] = 1'b0;  addr_rom[22970]='h000026e8;  wr_data_rom[22970]='h00000000;
    rd_cycle[22971] = 1'b1;  wr_cycle[22971] = 1'b0;  addr_rom[22971]='h000026ec;  wr_data_rom[22971]='h00000000;
    rd_cycle[22972] = 1'b1;  wr_cycle[22972] = 1'b0;  addr_rom[22972]='h000026f0;  wr_data_rom[22972]='h00000000;
    rd_cycle[22973] = 1'b1;  wr_cycle[22973] = 1'b0;  addr_rom[22973]='h000026f4;  wr_data_rom[22973]='h00000000;
    rd_cycle[22974] = 1'b1;  wr_cycle[22974] = 1'b0;  addr_rom[22974]='h000026f8;  wr_data_rom[22974]='h00000000;
    rd_cycle[22975] = 1'b1;  wr_cycle[22975] = 1'b0;  addr_rom[22975]='h000026fc;  wr_data_rom[22975]='h00000000;
    rd_cycle[22976] = 1'b1;  wr_cycle[22976] = 1'b0;  addr_rom[22976]='h00002700;  wr_data_rom[22976]='h00000000;
    rd_cycle[22977] = 1'b1;  wr_cycle[22977] = 1'b0;  addr_rom[22977]='h00002704;  wr_data_rom[22977]='h00000000;
    rd_cycle[22978] = 1'b1;  wr_cycle[22978] = 1'b0;  addr_rom[22978]='h00002708;  wr_data_rom[22978]='h00000000;
    rd_cycle[22979] = 1'b1;  wr_cycle[22979] = 1'b0;  addr_rom[22979]='h0000270c;  wr_data_rom[22979]='h00000000;
    rd_cycle[22980] = 1'b1;  wr_cycle[22980] = 1'b0;  addr_rom[22980]='h00002710;  wr_data_rom[22980]='h00000000;
    rd_cycle[22981] = 1'b1;  wr_cycle[22981] = 1'b0;  addr_rom[22981]='h00002714;  wr_data_rom[22981]='h00000000;
    rd_cycle[22982] = 1'b1;  wr_cycle[22982] = 1'b0;  addr_rom[22982]='h00002718;  wr_data_rom[22982]='h00000000;
    rd_cycle[22983] = 1'b1;  wr_cycle[22983] = 1'b0;  addr_rom[22983]='h0000271c;  wr_data_rom[22983]='h00000000;
    rd_cycle[22984] = 1'b1;  wr_cycle[22984] = 1'b0;  addr_rom[22984]='h00002720;  wr_data_rom[22984]='h00000000;
    rd_cycle[22985] = 1'b1;  wr_cycle[22985] = 1'b0;  addr_rom[22985]='h00002724;  wr_data_rom[22985]='h00000000;
    rd_cycle[22986] = 1'b1;  wr_cycle[22986] = 1'b0;  addr_rom[22986]='h00002728;  wr_data_rom[22986]='h00000000;
    rd_cycle[22987] = 1'b1;  wr_cycle[22987] = 1'b0;  addr_rom[22987]='h0000272c;  wr_data_rom[22987]='h00000000;
    rd_cycle[22988] = 1'b1;  wr_cycle[22988] = 1'b0;  addr_rom[22988]='h00002730;  wr_data_rom[22988]='h00000000;
    rd_cycle[22989] = 1'b1;  wr_cycle[22989] = 1'b0;  addr_rom[22989]='h00002734;  wr_data_rom[22989]='h00000000;
    rd_cycle[22990] = 1'b1;  wr_cycle[22990] = 1'b0;  addr_rom[22990]='h00002738;  wr_data_rom[22990]='h00000000;
    rd_cycle[22991] = 1'b1;  wr_cycle[22991] = 1'b0;  addr_rom[22991]='h0000273c;  wr_data_rom[22991]='h00000000;
    rd_cycle[22992] = 1'b1;  wr_cycle[22992] = 1'b0;  addr_rom[22992]='h00002740;  wr_data_rom[22992]='h00000000;
    rd_cycle[22993] = 1'b1;  wr_cycle[22993] = 1'b0;  addr_rom[22993]='h00002744;  wr_data_rom[22993]='h00000000;
    rd_cycle[22994] = 1'b1;  wr_cycle[22994] = 1'b0;  addr_rom[22994]='h00002748;  wr_data_rom[22994]='h00000000;
    rd_cycle[22995] = 1'b1;  wr_cycle[22995] = 1'b0;  addr_rom[22995]='h0000274c;  wr_data_rom[22995]='h00000000;
    rd_cycle[22996] = 1'b1;  wr_cycle[22996] = 1'b0;  addr_rom[22996]='h00002750;  wr_data_rom[22996]='h00000000;
    rd_cycle[22997] = 1'b1;  wr_cycle[22997] = 1'b0;  addr_rom[22997]='h00002754;  wr_data_rom[22997]='h00000000;
    rd_cycle[22998] = 1'b1;  wr_cycle[22998] = 1'b0;  addr_rom[22998]='h00002758;  wr_data_rom[22998]='h00000000;
    rd_cycle[22999] = 1'b1;  wr_cycle[22999] = 1'b0;  addr_rom[22999]='h0000275c;  wr_data_rom[22999]='h00000000;
    rd_cycle[23000] = 1'b1;  wr_cycle[23000] = 1'b0;  addr_rom[23000]='h00002760;  wr_data_rom[23000]='h00000000;
    rd_cycle[23001] = 1'b1;  wr_cycle[23001] = 1'b0;  addr_rom[23001]='h00002764;  wr_data_rom[23001]='h00000000;
    rd_cycle[23002] = 1'b1;  wr_cycle[23002] = 1'b0;  addr_rom[23002]='h00002768;  wr_data_rom[23002]='h00000000;
    rd_cycle[23003] = 1'b1;  wr_cycle[23003] = 1'b0;  addr_rom[23003]='h0000276c;  wr_data_rom[23003]='h00000000;
    rd_cycle[23004] = 1'b1;  wr_cycle[23004] = 1'b0;  addr_rom[23004]='h00002770;  wr_data_rom[23004]='h00000000;
    rd_cycle[23005] = 1'b1;  wr_cycle[23005] = 1'b0;  addr_rom[23005]='h00002774;  wr_data_rom[23005]='h00000000;
    rd_cycle[23006] = 1'b1;  wr_cycle[23006] = 1'b0;  addr_rom[23006]='h00002778;  wr_data_rom[23006]='h00000000;
    rd_cycle[23007] = 1'b1;  wr_cycle[23007] = 1'b0;  addr_rom[23007]='h0000277c;  wr_data_rom[23007]='h00000000;
    rd_cycle[23008] = 1'b1;  wr_cycle[23008] = 1'b0;  addr_rom[23008]='h00002780;  wr_data_rom[23008]='h00000000;
    rd_cycle[23009] = 1'b1;  wr_cycle[23009] = 1'b0;  addr_rom[23009]='h00002784;  wr_data_rom[23009]='h00000000;
    rd_cycle[23010] = 1'b1;  wr_cycle[23010] = 1'b0;  addr_rom[23010]='h00002788;  wr_data_rom[23010]='h00000000;
    rd_cycle[23011] = 1'b1;  wr_cycle[23011] = 1'b0;  addr_rom[23011]='h0000278c;  wr_data_rom[23011]='h00000000;
    rd_cycle[23012] = 1'b1;  wr_cycle[23012] = 1'b0;  addr_rom[23012]='h00002790;  wr_data_rom[23012]='h00000000;
    rd_cycle[23013] = 1'b1;  wr_cycle[23013] = 1'b0;  addr_rom[23013]='h00002794;  wr_data_rom[23013]='h00000000;
    rd_cycle[23014] = 1'b1;  wr_cycle[23014] = 1'b0;  addr_rom[23014]='h00002798;  wr_data_rom[23014]='h00000000;
    rd_cycle[23015] = 1'b1;  wr_cycle[23015] = 1'b0;  addr_rom[23015]='h0000279c;  wr_data_rom[23015]='h00000000;
    rd_cycle[23016] = 1'b1;  wr_cycle[23016] = 1'b0;  addr_rom[23016]='h000027a0;  wr_data_rom[23016]='h00000000;
    rd_cycle[23017] = 1'b1;  wr_cycle[23017] = 1'b0;  addr_rom[23017]='h000027a4;  wr_data_rom[23017]='h00000000;
    rd_cycle[23018] = 1'b1;  wr_cycle[23018] = 1'b0;  addr_rom[23018]='h000027a8;  wr_data_rom[23018]='h00000000;
    rd_cycle[23019] = 1'b1;  wr_cycle[23019] = 1'b0;  addr_rom[23019]='h000027ac;  wr_data_rom[23019]='h00000000;
    rd_cycle[23020] = 1'b1;  wr_cycle[23020] = 1'b0;  addr_rom[23020]='h000027b0;  wr_data_rom[23020]='h00000000;
    rd_cycle[23021] = 1'b1;  wr_cycle[23021] = 1'b0;  addr_rom[23021]='h000027b4;  wr_data_rom[23021]='h00000000;
    rd_cycle[23022] = 1'b1;  wr_cycle[23022] = 1'b0;  addr_rom[23022]='h000027b8;  wr_data_rom[23022]='h00000000;
    rd_cycle[23023] = 1'b1;  wr_cycle[23023] = 1'b0;  addr_rom[23023]='h000027bc;  wr_data_rom[23023]='h00000000;
    rd_cycle[23024] = 1'b1;  wr_cycle[23024] = 1'b0;  addr_rom[23024]='h000027c0;  wr_data_rom[23024]='h00000000;
    rd_cycle[23025] = 1'b1;  wr_cycle[23025] = 1'b0;  addr_rom[23025]='h000027c4;  wr_data_rom[23025]='h00000000;
    rd_cycle[23026] = 1'b1;  wr_cycle[23026] = 1'b0;  addr_rom[23026]='h000027c8;  wr_data_rom[23026]='h00000000;
    rd_cycle[23027] = 1'b1;  wr_cycle[23027] = 1'b0;  addr_rom[23027]='h000027cc;  wr_data_rom[23027]='h00000000;
    rd_cycle[23028] = 1'b1;  wr_cycle[23028] = 1'b0;  addr_rom[23028]='h000027d0;  wr_data_rom[23028]='h00000000;
    rd_cycle[23029] = 1'b1;  wr_cycle[23029] = 1'b0;  addr_rom[23029]='h000027d4;  wr_data_rom[23029]='h00000000;
    rd_cycle[23030] = 1'b1;  wr_cycle[23030] = 1'b0;  addr_rom[23030]='h000027d8;  wr_data_rom[23030]='h00000000;
    rd_cycle[23031] = 1'b1;  wr_cycle[23031] = 1'b0;  addr_rom[23031]='h000027dc;  wr_data_rom[23031]='h00000000;
    rd_cycle[23032] = 1'b1;  wr_cycle[23032] = 1'b0;  addr_rom[23032]='h000027e0;  wr_data_rom[23032]='h00000000;
    rd_cycle[23033] = 1'b1;  wr_cycle[23033] = 1'b0;  addr_rom[23033]='h000027e4;  wr_data_rom[23033]='h00000000;
    rd_cycle[23034] = 1'b1;  wr_cycle[23034] = 1'b0;  addr_rom[23034]='h000027e8;  wr_data_rom[23034]='h00000000;
    rd_cycle[23035] = 1'b1;  wr_cycle[23035] = 1'b0;  addr_rom[23035]='h000027ec;  wr_data_rom[23035]='h00000000;
    rd_cycle[23036] = 1'b1;  wr_cycle[23036] = 1'b0;  addr_rom[23036]='h000027f0;  wr_data_rom[23036]='h00000000;
    rd_cycle[23037] = 1'b1;  wr_cycle[23037] = 1'b0;  addr_rom[23037]='h000027f4;  wr_data_rom[23037]='h00000000;
    rd_cycle[23038] = 1'b1;  wr_cycle[23038] = 1'b0;  addr_rom[23038]='h000027f8;  wr_data_rom[23038]='h00000000;
    rd_cycle[23039] = 1'b1;  wr_cycle[23039] = 1'b0;  addr_rom[23039]='h000027fc;  wr_data_rom[23039]='h00000000;
    rd_cycle[23040] = 1'b1;  wr_cycle[23040] = 1'b0;  addr_rom[23040]='h00002800;  wr_data_rom[23040]='h00000000;
    rd_cycle[23041] = 1'b1;  wr_cycle[23041] = 1'b0;  addr_rom[23041]='h00002804;  wr_data_rom[23041]='h00000000;
    rd_cycle[23042] = 1'b1;  wr_cycle[23042] = 1'b0;  addr_rom[23042]='h00002808;  wr_data_rom[23042]='h00000000;
    rd_cycle[23043] = 1'b1;  wr_cycle[23043] = 1'b0;  addr_rom[23043]='h0000280c;  wr_data_rom[23043]='h00000000;
    rd_cycle[23044] = 1'b1;  wr_cycle[23044] = 1'b0;  addr_rom[23044]='h00002810;  wr_data_rom[23044]='h00000000;
    rd_cycle[23045] = 1'b1;  wr_cycle[23045] = 1'b0;  addr_rom[23045]='h00002814;  wr_data_rom[23045]='h00000000;
    rd_cycle[23046] = 1'b1;  wr_cycle[23046] = 1'b0;  addr_rom[23046]='h00002818;  wr_data_rom[23046]='h00000000;
    rd_cycle[23047] = 1'b1;  wr_cycle[23047] = 1'b0;  addr_rom[23047]='h0000281c;  wr_data_rom[23047]='h00000000;
    rd_cycle[23048] = 1'b1;  wr_cycle[23048] = 1'b0;  addr_rom[23048]='h00002820;  wr_data_rom[23048]='h00000000;
    rd_cycle[23049] = 1'b1;  wr_cycle[23049] = 1'b0;  addr_rom[23049]='h00002824;  wr_data_rom[23049]='h00000000;
    rd_cycle[23050] = 1'b1;  wr_cycle[23050] = 1'b0;  addr_rom[23050]='h00002828;  wr_data_rom[23050]='h00000000;
    rd_cycle[23051] = 1'b1;  wr_cycle[23051] = 1'b0;  addr_rom[23051]='h0000282c;  wr_data_rom[23051]='h00000000;
    rd_cycle[23052] = 1'b1;  wr_cycle[23052] = 1'b0;  addr_rom[23052]='h00002830;  wr_data_rom[23052]='h00000000;
    rd_cycle[23053] = 1'b1;  wr_cycle[23053] = 1'b0;  addr_rom[23053]='h00002834;  wr_data_rom[23053]='h00000000;
    rd_cycle[23054] = 1'b1;  wr_cycle[23054] = 1'b0;  addr_rom[23054]='h00002838;  wr_data_rom[23054]='h00000000;
    rd_cycle[23055] = 1'b1;  wr_cycle[23055] = 1'b0;  addr_rom[23055]='h0000283c;  wr_data_rom[23055]='h00000000;
    rd_cycle[23056] = 1'b1;  wr_cycle[23056] = 1'b0;  addr_rom[23056]='h00002840;  wr_data_rom[23056]='h00000000;
    rd_cycle[23057] = 1'b1;  wr_cycle[23057] = 1'b0;  addr_rom[23057]='h00002844;  wr_data_rom[23057]='h00000000;
    rd_cycle[23058] = 1'b1;  wr_cycle[23058] = 1'b0;  addr_rom[23058]='h00002848;  wr_data_rom[23058]='h00000000;
    rd_cycle[23059] = 1'b1;  wr_cycle[23059] = 1'b0;  addr_rom[23059]='h0000284c;  wr_data_rom[23059]='h00000000;
    rd_cycle[23060] = 1'b1;  wr_cycle[23060] = 1'b0;  addr_rom[23060]='h00002850;  wr_data_rom[23060]='h00000000;
    rd_cycle[23061] = 1'b1;  wr_cycle[23061] = 1'b0;  addr_rom[23061]='h00002854;  wr_data_rom[23061]='h00000000;
    rd_cycle[23062] = 1'b1;  wr_cycle[23062] = 1'b0;  addr_rom[23062]='h00002858;  wr_data_rom[23062]='h00000000;
    rd_cycle[23063] = 1'b1;  wr_cycle[23063] = 1'b0;  addr_rom[23063]='h0000285c;  wr_data_rom[23063]='h00000000;
    rd_cycle[23064] = 1'b1;  wr_cycle[23064] = 1'b0;  addr_rom[23064]='h00002860;  wr_data_rom[23064]='h00000000;
    rd_cycle[23065] = 1'b1;  wr_cycle[23065] = 1'b0;  addr_rom[23065]='h00002864;  wr_data_rom[23065]='h00000000;
    rd_cycle[23066] = 1'b1;  wr_cycle[23066] = 1'b0;  addr_rom[23066]='h00002868;  wr_data_rom[23066]='h00000000;
    rd_cycle[23067] = 1'b1;  wr_cycle[23067] = 1'b0;  addr_rom[23067]='h0000286c;  wr_data_rom[23067]='h00000000;
    rd_cycle[23068] = 1'b1;  wr_cycle[23068] = 1'b0;  addr_rom[23068]='h00002870;  wr_data_rom[23068]='h00000000;
    rd_cycle[23069] = 1'b1;  wr_cycle[23069] = 1'b0;  addr_rom[23069]='h00002874;  wr_data_rom[23069]='h00000000;
    rd_cycle[23070] = 1'b1;  wr_cycle[23070] = 1'b0;  addr_rom[23070]='h00002878;  wr_data_rom[23070]='h00000000;
    rd_cycle[23071] = 1'b1;  wr_cycle[23071] = 1'b0;  addr_rom[23071]='h0000287c;  wr_data_rom[23071]='h00000000;
    rd_cycle[23072] = 1'b1;  wr_cycle[23072] = 1'b0;  addr_rom[23072]='h00002880;  wr_data_rom[23072]='h00000000;
    rd_cycle[23073] = 1'b1;  wr_cycle[23073] = 1'b0;  addr_rom[23073]='h00002884;  wr_data_rom[23073]='h00000000;
    rd_cycle[23074] = 1'b1;  wr_cycle[23074] = 1'b0;  addr_rom[23074]='h00002888;  wr_data_rom[23074]='h00000000;
    rd_cycle[23075] = 1'b1;  wr_cycle[23075] = 1'b0;  addr_rom[23075]='h0000288c;  wr_data_rom[23075]='h00000000;
    rd_cycle[23076] = 1'b1;  wr_cycle[23076] = 1'b0;  addr_rom[23076]='h00002890;  wr_data_rom[23076]='h00000000;
    rd_cycle[23077] = 1'b1;  wr_cycle[23077] = 1'b0;  addr_rom[23077]='h00002894;  wr_data_rom[23077]='h00000000;
    rd_cycle[23078] = 1'b1;  wr_cycle[23078] = 1'b0;  addr_rom[23078]='h00002898;  wr_data_rom[23078]='h00000000;
    rd_cycle[23079] = 1'b1;  wr_cycle[23079] = 1'b0;  addr_rom[23079]='h0000289c;  wr_data_rom[23079]='h00000000;
    rd_cycle[23080] = 1'b1;  wr_cycle[23080] = 1'b0;  addr_rom[23080]='h000028a0;  wr_data_rom[23080]='h00000000;
    rd_cycle[23081] = 1'b1;  wr_cycle[23081] = 1'b0;  addr_rom[23081]='h000028a4;  wr_data_rom[23081]='h00000000;
    rd_cycle[23082] = 1'b1;  wr_cycle[23082] = 1'b0;  addr_rom[23082]='h000028a8;  wr_data_rom[23082]='h00000000;
    rd_cycle[23083] = 1'b1;  wr_cycle[23083] = 1'b0;  addr_rom[23083]='h000028ac;  wr_data_rom[23083]='h00000000;
    rd_cycle[23084] = 1'b1;  wr_cycle[23084] = 1'b0;  addr_rom[23084]='h000028b0;  wr_data_rom[23084]='h00000000;
    rd_cycle[23085] = 1'b1;  wr_cycle[23085] = 1'b0;  addr_rom[23085]='h000028b4;  wr_data_rom[23085]='h00000000;
    rd_cycle[23086] = 1'b1;  wr_cycle[23086] = 1'b0;  addr_rom[23086]='h000028b8;  wr_data_rom[23086]='h00000000;
    rd_cycle[23087] = 1'b1;  wr_cycle[23087] = 1'b0;  addr_rom[23087]='h000028bc;  wr_data_rom[23087]='h00000000;
    rd_cycle[23088] = 1'b1;  wr_cycle[23088] = 1'b0;  addr_rom[23088]='h000028c0;  wr_data_rom[23088]='h00000000;
    rd_cycle[23089] = 1'b1;  wr_cycle[23089] = 1'b0;  addr_rom[23089]='h000028c4;  wr_data_rom[23089]='h00000000;
    rd_cycle[23090] = 1'b1;  wr_cycle[23090] = 1'b0;  addr_rom[23090]='h000028c8;  wr_data_rom[23090]='h00000000;
    rd_cycle[23091] = 1'b1;  wr_cycle[23091] = 1'b0;  addr_rom[23091]='h000028cc;  wr_data_rom[23091]='h00000000;
    rd_cycle[23092] = 1'b1;  wr_cycle[23092] = 1'b0;  addr_rom[23092]='h000028d0;  wr_data_rom[23092]='h00000000;
    rd_cycle[23093] = 1'b1;  wr_cycle[23093] = 1'b0;  addr_rom[23093]='h000028d4;  wr_data_rom[23093]='h00000000;
    rd_cycle[23094] = 1'b1;  wr_cycle[23094] = 1'b0;  addr_rom[23094]='h000028d8;  wr_data_rom[23094]='h00000000;
    rd_cycle[23095] = 1'b1;  wr_cycle[23095] = 1'b0;  addr_rom[23095]='h000028dc;  wr_data_rom[23095]='h00000000;
    rd_cycle[23096] = 1'b1;  wr_cycle[23096] = 1'b0;  addr_rom[23096]='h000028e0;  wr_data_rom[23096]='h00000000;
    rd_cycle[23097] = 1'b1;  wr_cycle[23097] = 1'b0;  addr_rom[23097]='h000028e4;  wr_data_rom[23097]='h00000000;
    rd_cycle[23098] = 1'b1;  wr_cycle[23098] = 1'b0;  addr_rom[23098]='h000028e8;  wr_data_rom[23098]='h00000000;
    rd_cycle[23099] = 1'b1;  wr_cycle[23099] = 1'b0;  addr_rom[23099]='h000028ec;  wr_data_rom[23099]='h00000000;
    rd_cycle[23100] = 1'b1;  wr_cycle[23100] = 1'b0;  addr_rom[23100]='h000028f0;  wr_data_rom[23100]='h00000000;
    rd_cycle[23101] = 1'b1;  wr_cycle[23101] = 1'b0;  addr_rom[23101]='h000028f4;  wr_data_rom[23101]='h00000000;
    rd_cycle[23102] = 1'b1;  wr_cycle[23102] = 1'b0;  addr_rom[23102]='h000028f8;  wr_data_rom[23102]='h00000000;
    rd_cycle[23103] = 1'b1;  wr_cycle[23103] = 1'b0;  addr_rom[23103]='h000028fc;  wr_data_rom[23103]='h00000000;
    rd_cycle[23104] = 1'b1;  wr_cycle[23104] = 1'b0;  addr_rom[23104]='h00002900;  wr_data_rom[23104]='h00000000;
    rd_cycle[23105] = 1'b1;  wr_cycle[23105] = 1'b0;  addr_rom[23105]='h00002904;  wr_data_rom[23105]='h00000000;
    rd_cycle[23106] = 1'b1;  wr_cycle[23106] = 1'b0;  addr_rom[23106]='h00002908;  wr_data_rom[23106]='h00000000;
    rd_cycle[23107] = 1'b1;  wr_cycle[23107] = 1'b0;  addr_rom[23107]='h0000290c;  wr_data_rom[23107]='h00000000;
    rd_cycle[23108] = 1'b1;  wr_cycle[23108] = 1'b0;  addr_rom[23108]='h00002910;  wr_data_rom[23108]='h00000000;
    rd_cycle[23109] = 1'b1;  wr_cycle[23109] = 1'b0;  addr_rom[23109]='h00002914;  wr_data_rom[23109]='h00000000;
    rd_cycle[23110] = 1'b1;  wr_cycle[23110] = 1'b0;  addr_rom[23110]='h00002918;  wr_data_rom[23110]='h00000000;
    rd_cycle[23111] = 1'b1;  wr_cycle[23111] = 1'b0;  addr_rom[23111]='h0000291c;  wr_data_rom[23111]='h00000000;
    rd_cycle[23112] = 1'b1;  wr_cycle[23112] = 1'b0;  addr_rom[23112]='h00002920;  wr_data_rom[23112]='h00000000;
    rd_cycle[23113] = 1'b1;  wr_cycle[23113] = 1'b0;  addr_rom[23113]='h00002924;  wr_data_rom[23113]='h00000000;
    rd_cycle[23114] = 1'b1;  wr_cycle[23114] = 1'b0;  addr_rom[23114]='h00002928;  wr_data_rom[23114]='h00000000;
    rd_cycle[23115] = 1'b1;  wr_cycle[23115] = 1'b0;  addr_rom[23115]='h0000292c;  wr_data_rom[23115]='h00000000;
    rd_cycle[23116] = 1'b1;  wr_cycle[23116] = 1'b0;  addr_rom[23116]='h00002930;  wr_data_rom[23116]='h00000000;
    rd_cycle[23117] = 1'b1;  wr_cycle[23117] = 1'b0;  addr_rom[23117]='h00002934;  wr_data_rom[23117]='h00000000;
    rd_cycle[23118] = 1'b1;  wr_cycle[23118] = 1'b0;  addr_rom[23118]='h00002938;  wr_data_rom[23118]='h00000000;
    rd_cycle[23119] = 1'b1;  wr_cycle[23119] = 1'b0;  addr_rom[23119]='h0000293c;  wr_data_rom[23119]='h00000000;
    rd_cycle[23120] = 1'b1;  wr_cycle[23120] = 1'b0;  addr_rom[23120]='h00002940;  wr_data_rom[23120]='h00000000;
    rd_cycle[23121] = 1'b1;  wr_cycle[23121] = 1'b0;  addr_rom[23121]='h00002944;  wr_data_rom[23121]='h00000000;
    rd_cycle[23122] = 1'b1;  wr_cycle[23122] = 1'b0;  addr_rom[23122]='h00002948;  wr_data_rom[23122]='h00000000;
    rd_cycle[23123] = 1'b1;  wr_cycle[23123] = 1'b0;  addr_rom[23123]='h0000294c;  wr_data_rom[23123]='h00000000;
    rd_cycle[23124] = 1'b1;  wr_cycle[23124] = 1'b0;  addr_rom[23124]='h00002950;  wr_data_rom[23124]='h00000000;
    rd_cycle[23125] = 1'b1;  wr_cycle[23125] = 1'b0;  addr_rom[23125]='h00002954;  wr_data_rom[23125]='h00000000;
    rd_cycle[23126] = 1'b1;  wr_cycle[23126] = 1'b0;  addr_rom[23126]='h00002958;  wr_data_rom[23126]='h00000000;
    rd_cycle[23127] = 1'b1;  wr_cycle[23127] = 1'b0;  addr_rom[23127]='h0000295c;  wr_data_rom[23127]='h00000000;
    rd_cycle[23128] = 1'b1;  wr_cycle[23128] = 1'b0;  addr_rom[23128]='h00002960;  wr_data_rom[23128]='h00000000;
    rd_cycle[23129] = 1'b1;  wr_cycle[23129] = 1'b0;  addr_rom[23129]='h00002964;  wr_data_rom[23129]='h00000000;
    rd_cycle[23130] = 1'b1;  wr_cycle[23130] = 1'b0;  addr_rom[23130]='h00002968;  wr_data_rom[23130]='h00000000;
    rd_cycle[23131] = 1'b1;  wr_cycle[23131] = 1'b0;  addr_rom[23131]='h0000296c;  wr_data_rom[23131]='h00000000;
    rd_cycle[23132] = 1'b1;  wr_cycle[23132] = 1'b0;  addr_rom[23132]='h00002970;  wr_data_rom[23132]='h00000000;
    rd_cycle[23133] = 1'b1;  wr_cycle[23133] = 1'b0;  addr_rom[23133]='h00002974;  wr_data_rom[23133]='h00000000;
    rd_cycle[23134] = 1'b1;  wr_cycle[23134] = 1'b0;  addr_rom[23134]='h00002978;  wr_data_rom[23134]='h00000000;
    rd_cycle[23135] = 1'b1;  wr_cycle[23135] = 1'b0;  addr_rom[23135]='h0000297c;  wr_data_rom[23135]='h00000000;
    rd_cycle[23136] = 1'b1;  wr_cycle[23136] = 1'b0;  addr_rom[23136]='h00002980;  wr_data_rom[23136]='h00000000;
    rd_cycle[23137] = 1'b1;  wr_cycle[23137] = 1'b0;  addr_rom[23137]='h00002984;  wr_data_rom[23137]='h00000000;
    rd_cycle[23138] = 1'b1;  wr_cycle[23138] = 1'b0;  addr_rom[23138]='h00002988;  wr_data_rom[23138]='h00000000;
    rd_cycle[23139] = 1'b1;  wr_cycle[23139] = 1'b0;  addr_rom[23139]='h0000298c;  wr_data_rom[23139]='h00000000;
    rd_cycle[23140] = 1'b1;  wr_cycle[23140] = 1'b0;  addr_rom[23140]='h00002990;  wr_data_rom[23140]='h00000000;
    rd_cycle[23141] = 1'b1;  wr_cycle[23141] = 1'b0;  addr_rom[23141]='h00002994;  wr_data_rom[23141]='h00000000;
    rd_cycle[23142] = 1'b1;  wr_cycle[23142] = 1'b0;  addr_rom[23142]='h00002998;  wr_data_rom[23142]='h00000000;
    rd_cycle[23143] = 1'b1;  wr_cycle[23143] = 1'b0;  addr_rom[23143]='h0000299c;  wr_data_rom[23143]='h00000000;
    rd_cycle[23144] = 1'b1;  wr_cycle[23144] = 1'b0;  addr_rom[23144]='h000029a0;  wr_data_rom[23144]='h00000000;
    rd_cycle[23145] = 1'b1;  wr_cycle[23145] = 1'b0;  addr_rom[23145]='h000029a4;  wr_data_rom[23145]='h00000000;
    rd_cycle[23146] = 1'b1;  wr_cycle[23146] = 1'b0;  addr_rom[23146]='h000029a8;  wr_data_rom[23146]='h00000000;
    rd_cycle[23147] = 1'b1;  wr_cycle[23147] = 1'b0;  addr_rom[23147]='h000029ac;  wr_data_rom[23147]='h00000000;
    rd_cycle[23148] = 1'b1;  wr_cycle[23148] = 1'b0;  addr_rom[23148]='h000029b0;  wr_data_rom[23148]='h00000000;
    rd_cycle[23149] = 1'b1;  wr_cycle[23149] = 1'b0;  addr_rom[23149]='h000029b4;  wr_data_rom[23149]='h00000000;
    rd_cycle[23150] = 1'b1;  wr_cycle[23150] = 1'b0;  addr_rom[23150]='h000029b8;  wr_data_rom[23150]='h00000000;
    rd_cycle[23151] = 1'b1;  wr_cycle[23151] = 1'b0;  addr_rom[23151]='h000029bc;  wr_data_rom[23151]='h00000000;
    rd_cycle[23152] = 1'b1;  wr_cycle[23152] = 1'b0;  addr_rom[23152]='h000029c0;  wr_data_rom[23152]='h00000000;
    rd_cycle[23153] = 1'b1;  wr_cycle[23153] = 1'b0;  addr_rom[23153]='h000029c4;  wr_data_rom[23153]='h00000000;
    rd_cycle[23154] = 1'b1;  wr_cycle[23154] = 1'b0;  addr_rom[23154]='h000029c8;  wr_data_rom[23154]='h00000000;
    rd_cycle[23155] = 1'b1;  wr_cycle[23155] = 1'b0;  addr_rom[23155]='h000029cc;  wr_data_rom[23155]='h00000000;
    rd_cycle[23156] = 1'b1;  wr_cycle[23156] = 1'b0;  addr_rom[23156]='h000029d0;  wr_data_rom[23156]='h00000000;
    rd_cycle[23157] = 1'b1;  wr_cycle[23157] = 1'b0;  addr_rom[23157]='h000029d4;  wr_data_rom[23157]='h00000000;
    rd_cycle[23158] = 1'b1;  wr_cycle[23158] = 1'b0;  addr_rom[23158]='h000029d8;  wr_data_rom[23158]='h00000000;
    rd_cycle[23159] = 1'b1;  wr_cycle[23159] = 1'b0;  addr_rom[23159]='h000029dc;  wr_data_rom[23159]='h00000000;
    rd_cycle[23160] = 1'b1;  wr_cycle[23160] = 1'b0;  addr_rom[23160]='h000029e0;  wr_data_rom[23160]='h00000000;
    rd_cycle[23161] = 1'b1;  wr_cycle[23161] = 1'b0;  addr_rom[23161]='h000029e4;  wr_data_rom[23161]='h00000000;
    rd_cycle[23162] = 1'b1;  wr_cycle[23162] = 1'b0;  addr_rom[23162]='h000029e8;  wr_data_rom[23162]='h00000000;
    rd_cycle[23163] = 1'b1;  wr_cycle[23163] = 1'b0;  addr_rom[23163]='h000029ec;  wr_data_rom[23163]='h00000000;
    rd_cycle[23164] = 1'b1;  wr_cycle[23164] = 1'b0;  addr_rom[23164]='h000029f0;  wr_data_rom[23164]='h00000000;
    rd_cycle[23165] = 1'b1;  wr_cycle[23165] = 1'b0;  addr_rom[23165]='h000029f4;  wr_data_rom[23165]='h00000000;
    rd_cycle[23166] = 1'b1;  wr_cycle[23166] = 1'b0;  addr_rom[23166]='h000029f8;  wr_data_rom[23166]='h00000000;
    rd_cycle[23167] = 1'b1;  wr_cycle[23167] = 1'b0;  addr_rom[23167]='h000029fc;  wr_data_rom[23167]='h00000000;
    rd_cycle[23168] = 1'b1;  wr_cycle[23168] = 1'b0;  addr_rom[23168]='h00002a00;  wr_data_rom[23168]='h00000000;
    rd_cycle[23169] = 1'b1;  wr_cycle[23169] = 1'b0;  addr_rom[23169]='h00002a04;  wr_data_rom[23169]='h00000000;
    rd_cycle[23170] = 1'b1;  wr_cycle[23170] = 1'b0;  addr_rom[23170]='h00002a08;  wr_data_rom[23170]='h00000000;
    rd_cycle[23171] = 1'b1;  wr_cycle[23171] = 1'b0;  addr_rom[23171]='h00002a0c;  wr_data_rom[23171]='h00000000;
    rd_cycle[23172] = 1'b1;  wr_cycle[23172] = 1'b0;  addr_rom[23172]='h00002a10;  wr_data_rom[23172]='h00000000;
    rd_cycle[23173] = 1'b1;  wr_cycle[23173] = 1'b0;  addr_rom[23173]='h00002a14;  wr_data_rom[23173]='h00000000;
    rd_cycle[23174] = 1'b1;  wr_cycle[23174] = 1'b0;  addr_rom[23174]='h00002a18;  wr_data_rom[23174]='h00000000;
    rd_cycle[23175] = 1'b1;  wr_cycle[23175] = 1'b0;  addr_rom[23175]='h00002a1c;  wr_data_rom[23175]='h00000000;
    rd_cycle[23176] = 1'b1;  wr_cycle[23176] = 1'b0;  addr_rom[23176]='h00002a20;  wr_data_rom[23176]='h00000000;
    rd_cycle[23177] = 1'b1;  wr_cycle[23177] = 1'b0;  addr_rom[23177]='h00002a24;  wr_data_rom[23177]='h00000000;
    rd_cycle[23178] = 1'b1;  wr_cycle[23178] = 1'b0;  addr_rom[23178]='h00002a28;  wr_data_rom[23178]='h00000000;
    rd_cycle[23179] = 1'b1;  wr_cycle[23179] = 1'b0;  addr_rom[23179]='h00002a2c;  wr_data_rom[23179]='h00000000;
    rd_cycle[23180] = 1'b1;  wr_cycle[23180] = 1'b0;  addr_rom[23180]='h00002a30;  wr_data_rom[23180]='h00000000;
    rd_cycle[23181] = 1'b1;  wr_cycle[23181] = 1'b0;  addr_rom[23181]='h00002a34;  wr_data_rom[23181]='h00000000;
    rd_cycle[23182] = 1'b1;  wr_cycle[23182] = 1'b0;  addr_rom[23182]='h00002a38;  wr_data_rom[23182]='h00000000;
    rd_cycle[23183] = 1'b1;  wr_cycle[23183] = 1'b0;  addr_rom[23183]='h00002a3c;  wr_data_rom[23183]='h00000000;
    rd_cycle[23184] = 1'b1;  wr_cycle[23184] = 1'b0;  addr_rom[23184]='h00002a40;  wr_data_rom[23184]='h00000000;
    rd_cycle[23185] = 1'b1;  wr_cycle[23185] = 1'b0;  addr_rom[23185]='h00002a44;  wr_data_rom[23185]='h00000000;
    rd_cycle[23186] = 1'b1;  wr_cycle[23186] = 1'b0;  addr_rom[23186]='h00002a48;  wr_data_rom[23186]='h00000000;
    rd_cycle[23187] = 1'b1;  wr_cycle[23187] = 1'b0;  addr_rom[23187]='h00002a4c;  wr_data_rom[23187]='h00000000;
    rd_cycle[23188] = 1'b1;  wr_cycle[23188] = 1'b0;  addr_rom[23188]='h00002a50;  wr_data_rom[23188]='h00000000;
    rd_cycle[23189] = 1'b1;  wr_cycle[23189] = 1'b0;  addr_rom[23189]='h00002a54;  wr_data_rom[23189]='h00000000;
    rd_cycle[23190] = 1'b1;  wr_cycle[23190] = 1'b0;  addr_rom[23190]='h00002a58;  wr_data_rom[23190]='h00000000;
    rd_cycle[23191] = 1'b1;  wr_cycle[23191] = 1'b0;  addr_rom[23191]='h00002a5c;  wr_data_rom[23191]='h00000000;
    rd_cycle[23192] = 1'b1;  wr_cycle[23192] = 1'b0;  addr_rom[23192]='h00002a60;  wr_data_rom[23192]='h00000000;
    rd_cycle[23193] = 1'b1;  wr_cycle[23193] = 1'b0;  addr_rom[23193]='h00002a64;  wr_data_rom[23193]='h00000000;
    rd_cycle[23194] = 1'b1;  wr_cycle[23194] = 1'b0;  addr_rom[23194]='h00002a68;  wr_data_rom[23194]='h00000000;
    rd_cycle[23195] = 1'b1;  wr_cycle[23195] = 1'b0;  addr_rom[23195]='h00002a6c;  wr_data_rom[23195]='h00000000;
    rd_cycle[23196] = 1'b1;  wr_cycle[23196] = 1'b0;  addr_rom[23196]='h00002a70;  wr_data_rom[23196]='h00000000;
    rd_cycle[23197] = 1'b1;  wr_cycle[23197] = 1'b0;  addr_rom[23197]='h00002a74;  wr_data_rom[23197]='h00000000;
    rd_cycle[23198] = 1'b1;  wr_cycle[23198] = 1'b0;  addr_rom[23198]='h00002a78;  wr_data_rom[23198]='h00000000;
    rd_cycle[23199] = 1'b1;  wr_cycle[23199] = 1'b0;  addr_rom[23199]='h00002a7c;  wr_data_rom[23199]='h00000000;
    rd_cycle[23200] = 1'b1;  wr_cycle[23200] = 1'b0;  addr_rom[23200]='h00002a80;  wr_data_rom[23200]='h00000000;
    rd_cycle[23201] = 1'b1;  wr_cycle[23201] = 1'b0;  addr_rom[23201]='h00002a84;  wr_data_rom[23201]='h00000000;
    rd_cycle[23202] = 1'b1;  wr_cycle[23202] = 1'b0;  addr_rom[23202]='h00002a88;  wr_data_rom[23202]='h00000000;
    rd_cycle[23203] = 1'b1;  wr_cycle[23203] = 1'b0;  addr_rom[23203]='h00002a8c;  wr_data_rom[23203]='h00000000;
    rd_cycle[23204] = 1'b1;  wr_cycle[23204] = 1'b0;  addr_rom[23204]='h00002a90;  wr_data_rom[23204]='h00000000;
    rd_cycle[23205] = 1'b1;  wr_cycle[23205] = 1'b0;  addr_rom[23205]='h00002a94;  wr_data_rom[23205]='h00000000;
    rd_cycle[23206] = 1'b1;  wr_cycle[23206] = 1'b0;  addr_rom[23206]='h00002a98;  wr_data_rom[23206]='h00000000;
    rd_cycle[23207] = 1'b1;  wr_cycle[23207] = 1'b0;  addr_rom[23207]='h00002a9c;  wr_data_rom[23207]='h00000000;
    rd_cycle[23208] = 1'b1;  wr_cycle[23208] = 1'b0;  addr_rom[23208]='h00002aa0;  wr_data_rom[23208]='h00000000;
    rd_cycle[23209] = 1'b1;  wr_cycle[23209] = 1'b0;  addr_rom[23209]='h00002aa4;  wr_data_rom[23209]='h00000000;
    rd_cycle[23210] = 1'b1;  wr_cycle[23210] = 1'b0;  addr_rom[23210]='h00002aa8;  wr_data_rom[23210]='h00000000;
    rd_cycle[23211] = 1'b1;  wr_cycle[23211] = 1'b0;  addr_rom[23211]='h00002aac;  wr_data_rom[23211]='h00000000;
    rd_cycle[23212] = 1'b1;  wr_cycle[23212] = 1'b0;  addr_rom[23212]='h00002ab0;  wr_data_rom[23212]='h00000000;
    rd_cycle[23213] = 1'b1;  wr_cycle[23213] = 1'b0;  addr_rom[23213]='h00002ab4;  wr_data_rom[23213]='h00000000;
    rd_cycle[23214] = 1'b1;  wr_cycle[23214] = 1'b0;  addr_rom[23214]='h00002ab8;  wr_data_rom[23214]='h00000000;
    rd_cycle[23215] = 1'b1;  wr_cycle[23215] = 1'b0;  addr_rom[23215]='h00002abc;  wr_data_rom[23215]='h00000000;
    rd_cycle[23216] = 1'b1;  wr_cycle[23216] = 1'b0;  addr_rom[23216]='h00002ac0;  wr_data_rom[23216]='h00000000;
    rd_cycle[23217] = 1'b1;  wr_cycle[23217] = 1'b0;  addr_rom[23217]='h00002ac4;  wr_data_rom[23217]='h00000000;
    rd_cycle[23218] = 1'b1;  wr_cycle[23218] = 1'b0;  addr_rom[23218]='h00002ac8;  wr_data_rom[23218]='h00000000;
    rd_cycle[23219] = 1'b1;  wr_cycle[23219] = 1'b0;  addr_rom[23219]='h00002acc;  wr_data_rom[23219]='h00000000;
    rd_cycle[23220] = 1'b1;  wr_cycle[23220] = 1'b0;  addr_rom[23220]='h00002ad0;  wr_data_rom[23220]='h00000000;
    rd_cycle[23221] = 1'b1;  wr_cycle[23221] = 1'b0;  addr_rom[23221]='h00002ad4;  wr_data_rom[23221]='h00000000;
    rd_cycle[23222] = 1'b1;  wr_cycle[23222] = 1'b0;  addr_rom[23222]='h00002ad8;  wr_data_rom[23222]='h00000000;
    rd_cycle[23223] = 1'b1;  wr_cycle[23223] = 1'b0;  addr_rom[23223]='h00002adc;  wr_data_rom[23223]='h00000000;
    rd_cycle[23224] = 1'b1;  wr_cycle[23224] = 1'b0;  addr_rom[23224]='h00002ae0;  wr_data_rom[23224]='h00000000;
    rd_cycle[23225] = 1'b1;  wr_cycle[23225] = 1'b0;  addr_rom[23225]='h00002ae4;  wr_data_rom[23225]='h00000000;
    rd_cycle[23226] = 1'b1;  wr_cycle[23226] = 1'b0;  addr_rom[23226]='h00002ae8;  wr_data_rom[23226]='h00000000;
    rd_cycle[23227] = 1'b1;  wr_cycle[23227] = 1'b0;  addr_rom[23227]='h00002aec;  wr_data_rom[23227]='h00000000;
    rd_cycle[23228] = 1'b1;  wr_cycle[23228] = 1'b0;  addr_rom[23228]='h00002af0;  wr_data_rom[23228]='h00000000;
    rd_cycle[23229] = 1'b1;  wr_cycle[23229] = 1'b0;  addr_rom[23229]='h00002af4;  wr_data_rom[23229]='h00000000;
    rd_cycle[23230] = 1'b1;  wr_cycle[23230] = 1'b0;  addr_rom[23230]='h00002af8;  wr_data_rom[23230]='h00000000;
    rd_cycle[23231] = 1'b1;  wr_cycle[23231] = 1'b0;  addr_rom[23231]='h00002afc;  wr_data_rom[23231]='h00000000;
    rd_cycle[23232] = 1'b1;  wr_cycle[23232] = 1'b0;  addr_rom[23232]='h00002b00;  wr_data_rom[23232]='h00000000;
    rd_cycle[23233] = 1'b1;  wr_cycle[23233] = 1'b0;  addr_rom[23233]='h00002b04;  wr_data_rom[23233]='h00000000;
    rd_cycle[23234] = 1'b1;  wr_cycle[23234] = 1'b0;  addr_rom[23234]='h00002b08;  wr_data_rom[23234]='h00000000;
    rd_cycle[23235] = 1'b1;  wr_cycle[23235] = 1'b0;  addr_rom[23235]='h00002b0c;  wr_data_rom[23235]='h00000000;
    rd_cycle[23236] = 1'b1;  wr_cycle[23236] = 1'b0;  addr_rom[23236]='h00002b10;  wr_data_rom[23236]='h00000000;
    rd_cycle[23237] = 1'b1;  wr_cycle[23237] = 1'b0;  addr_rom[23237]='h00002b14;  wr_data_rom[23237]='h00000000;
    rd_cycle[23238] = 1'b1;  wr_cycle[23238] = 1'b0;  addr_rom[23238]='h00002b18;  wr_data_rom[23238]='h00000000;
    rd_cycle[23239] = 1'b1;  wr_cycle[23239] = 1'b0;  addr_rom[23239]='h00002b1c;  wr_data_rom[23239]='h00000000;
    rd_cycle[23240] = 1'b1;  wr_cycle[23240] = 1'b0;  addr_rom[23240]='h00002b20;  wr_data_rom[23240]='h00000000;
    rd_cycle[23241] = 1'b1;  wr_cycle[23241] = 1'b0;  addr_rom[23241]='h00002b24;  wr_data_rom[23241]='h00000000;
    rd_cycle[23242] = 1'b1;  wr_cycle[23242] = 1'b0;  addr_rom[23242]='h00002b28;  wr_data_rom[23242]='h00000000;
    rd_cycle[23243] = 1'b1;  wr_cycle[23243] = 1'b0;  addr_rom[23243]='h00002b2c;  wr_data_rom[23243]='h00000000;
    rd_cycle[23244] = 1'b1;  wr_cycle[23244] = 1'b0;  addr_rom[23244]='h00002b30;  wr_data_rom[23244]='h00000000;
    rd_cycle[23245] = 1'b1;  wr_cycle[23245] = 1'b0;  addr_rom[23245]='h00002b34;  wr_data_rom[23245]='h00000000;
    rd_cycle[23246] = 1'b1;  wr_cycle[23246] = 1'b0;  addr_rom[23246]='h00002b38;  wr_data_rom[23246]='h00000000;
    rd_cycle[23247] = 1'b1;  wr_cycle[23247] = 1'b0;  addr_rom[23247]='h00002b3c;  wr_data_rom[23247]='h00000000;
    rd_cycle[23248] = 1'b1;  wr_cycle[23248] = 1'b0;  addr_rom[23248]='h00002b40;  wr_data_rom[23248]='h00000000;
    rd_cycle[23249] = 1'b1;  wr_cycle[23249] = 1'b0;  addr_rom[23249]='h00002b44;  wr_data_rom[23249]='h00000000;
    rd_cycle[23250] = 1'b1;  wr_cycle[23250] = 1'b0;  addr_rom[23250]='h00002b48;  wr_data_rom[23250]='h00000000;
    rd_cycle[23251] = 1'b1;  wr_cycle[23251] = 1'b0;  addr_rom[23251]='h00002b4c;  wr_data_rom[23251]='h00000000;
    rd_cycle[23252] = 1'b1;  wr_cycle[23252] = 1'b0;  addr_rom[23252]='h00002b50;  wr_data_rom[23252]='h00000000;
    rd_cycle[23253] = 1'b1;  wr_cycle[23253] = 1'b0;  addr_rom[23253]='h00002b54;  wr_data_rom[23253]='h00000000;
    rd_cycle[23254] = 1'b1;  wr_cycle[23254] = 1'b0;  addr_rom[23254]='h00002b58;  wr_data_rom[23254]='h00000000;
    rd_cycle[23255] = 1'b1;  wr_cycle[23255] = 1'b0;  addr_rom[23255]='h00002b5c;  wr_data_rom[23255]='h00000000;
    rd_cycle[23256] = 1'b1;  wr_cycle[23256] = 1'b0;  addr_rom[23256]='h00002b60;  wr_data_rom[23256]='h00000000;
    rd_cycle[23257] = 1'b1;  wr_cycle[23257] = 1'b0;  addr_rom[23257]='h00002b64;  wr_data_rom[23257]='h00000000;
    rd_cycle[23258] = 1'b1;  wr_cycle[23258] = 1'b0;  addr_rom[23258]='h00002b68;  wr_data_rom[23258]='h00000000;
    rd_cycle[23259] = 1'b1;  wr_cycle[23259] = 1'b0;  addr_rom[23259]='h00002b6c;  wr_data_rom[23259]='h00000000;
    rd_cycle[23260] = 1'b1;  wr_cycle[23260] = 1'b0;  addr_rom[23260]='h00002b70;  wr_data_rom[23260]='h00000000;
    rd_cycle[23261] = 1'b1;  wr_cycle[23261] = 1'b0;  addr_rom[23261]='h00002b74;  wr_data_rom[23261]='h00000000;
    rd_cycle[23262] = 1'b1;  wr_cycle[23262] = 1'b0;  addr_rom[23262]='h00002b78;  wr_data_rom[23262]='h00000000;
    rd_cycle[23263] = 1'b1;  wr_cycle[23263] = 1'b0;  addr_rom[23263]='h00002b7c;  wr_data_rom[23263]='h00000000;
    rd_cycle[23264] = 1'b1;  wr_cycle[23264] = 1'b0;  addr_rom[23264]='h00002b80;  wr_data_rom[23264]='h00000000;
    rd_cycle[23265] = 1'b1;  wr_cycle[23265] = 1'b0;  addr_rom[23265]='h00002b84;  wr_data_rom[23265]='h00000000;
    rd_cycle[23266] = 1'b1;  wr_cycle[23266] = 1'b0;  addr_rom[23266]='h00002b88;  wr_data_rom[23266]='h00000000;
    rd_cycle[23267] = 1'b1;  wr_cycle[23267] = 1'b0;  addr_rom[23267]='h00002b8c;  wr_data_rom[23267]='h00000000;
    rd_cycle[23268] = 1'b1;  wr_cycle[23268] = 1'b0;  addr_rom[23268]='h00002b90;  wr_data_rom[23268]='h00000000;
    rd_cycle[23269] = 1'b1;  wr_cycle[23269] = 1'b0;  addr_rom[23269]='h00002b94;  wr_data_rom[23269]='h00000000;
    rd_cycle[23270] = 1'b1;  wr_cycle[23270] = 1'b0;  addr_rom[23270]='h00002b98;  wr_data_rom[23270]='h00000000;
    rd_cycle[23271] = 1'b1;  wr_cycle[23271] = 1'b0;  addr_rom[23271]='h00002b9c;  wr_data_rom[23271]='h00000000;
    rd_cycle[23272] = 1'b1;  wr_cycle[23272] = 1'b0;  addr_rom[23272]='h00002ba0;  wr_data_rom[23272]='h00000000;
    rd_cycle[23273] = 1'b1;  wr_cycle[23273] = 1'b0;  addr_rom[23273]='h00002ba4;  wr_data_rom[23273]='h00000000;
    rd_cycle[23274] = 1'b1;  wr_cycle[23274] = 1'b0;  addr_rom[23274]='h00002ba8;  wr_data_rom[23274]='h00000000;
    rd_cycle[23275] = 1'b1;  wr_cycle[23275] = 1'b0;  addr_rom[23275]='h00002bac;  wr_data_rom[23275]='h00000000;
    rd_cycle[23276] = 1'b1;  wr_cycle[23276] = 1'b0;  addr_rom[23276]='h00002bb0;  wr_data_rom[23276]='h00000000;
    rd_cycle[23277] = 1'b1;  wr_cycle[23277] = 1'b0;  addr_rom[23277]='h00002bb4;  wr_data_rom[23277]='h00000000;
    rd_cycle[23278] = 1'b1;  wr_cycle[23278] = 1'b0;  addr_rom[23278]='h00002bb8;  wr_data_rom[23278]='h00000000;
    rd_cycle[23279] = 1'b1;  wr_cycle[23279] = 1'b0;  addr_rom[23279]='h00002bbc;  wr_data_rom[23279]='h00000000;
    rd_cycle[23280] = 1'b1;  wr_cycle[23280] = 1'b0;  addr_rom[23280]='h00002bc0;  wr_data_rom[23280]='h00000000;
    rd_cycle[23281] = 1'b1;  wr_cycle[23281] = 1'b0;  addr_rom[23281]='h00002bc4;  wr_data_rom[23281]='h00000000;
    rd_cycle[23282] = 1'b1;  wr_cycle[23282] = 1'b0;  addr_rom[23282]='h00002bc8;  wr_data_rom[23282]='h00000000;
    rd_cycle[23283] = 1'b1;  wr_cycle[23283] = 1'b0;  addr_rom[23283]='h00002bcc;  wr_data_rom[23283]='h00000000;
    rd_cycle[23284] = 1'b1;  wr_cycle[23284] = 1'b0;  addr_rom[23284]='h00002bd0;  wr_data_rom[23284]='h00000000;
    rd_cycle[23285] = 1'b1;  wr_cycle[23285] = 1'b0;  addr_rom[23285]='h00002bd4;  wr_data_rom[23285]='h00000000;
    rd_cycle[23286] = 1'b1;  wr_cycle[23286] = 1'b0;  addr_rom[23286]='h00002bd8;  wr_data_rom[23286]='h00000000;
    rd_cycle[23287] = 1'b1;  wr_cycle[23287] = 1'b0;  addr_rom[23287]='h00002bdc;  wr_data_rom[23287]='h00000000;
    rd_cycle[23288] = 1'b1;  wr_cycle[23288] = 1'b0;  addr_rom[23288]='h00002be0;  wr_data_rom[23288]='h00000000;
    rd_cycle[23289] = 1'b1;  wr_cycle[23289] = 1'b0;  addr_rom[23289]='h00002be4;  wr_data_rom[23289]='h00000000;
    rd_cycle[23290] = 1'b1;  wr_cycle[23290] = 1'b0;  addr_rom[23290]='h00002be8;  wr_data_rom[23290]='h00000000;
    rd_cycle[23291] = 1'b1;  wr_cycle[23291] = 1'b0;  addr_rom[23291]='h00002bec;  wr_data_rom[23291]='h00000000;
    rd_cycle[23292] = 1'b1;  wr_cycle[23292] = 1'b0;  addr_rom[23292]='h00002bf0;  wr_data_rom[23292]='h00000000;
    rd_cycle[23293] = 1'b1;  wr_cycle[23293] = 1'b0;  addr_rom[23293]='h00002bf4;  wr_data_rom[23293]='h00000000;
    rd_cycle[23294] = 1'b1;  wr_cycle[23294] = 1'b0;  addr_rom[23294]='h00002bf8;  wr_data_rom[23294]='h00000000;
    rd_cycle[23295] = 1'b1;  wr_cycle[23295] = 1'b0;  addr_rom[23295]='h00002bfc;  wr_data_rom[23295]='h00000000;
    rd_cycle[23296] = 1'b1;  wr_cycle[23296] = 1'b0;  addr_rom[23296]='h00002c00;  wr_data_rom[23296]='h00000000;
    rd_cycle[23297] = 1'b1;  wr_cycle[23297] = 1'b0;  addr_rom[23297]='h00002c04;  wr_data_rom[23297]='h00000000;
    rd_cycle[23298] = 1'b1;  wr_cycle[23298] = 1'b0;  addr_rom[23298]='h00002c08;  wr_data_rom[23298]='h00000000;
    rd_cycle[23299] = 1'b1;  wr_cycle[23299] = 1'b0;  addr_rom[23299]='h00002c0c;  wr_data_rom[23299]='h00000000;
    rd_cycle[23300] = 1'b1;  wr_cycle[23300] = 1'b0;  addr_rom[23300]='h00002c10;  wr_data_rom[23300]='h00000000;
    rd_cycle[23301] = 1'b1;  wr_cycle[23301] = 1'b0;  addr_rom[23301]='h00002c14;  wr_data_rom[23301]='h00000000;
    rd_cycle[23302] = 1'b1;  wr_cycle[23302] = 1'b0;  addr_rom[23302]='h00002c18;  wr_data_rom[23302]='h00000000;
    rd_cycle[23303] = 1'b1;  wr_cycle[23303] = 1'b0;  addr_rom[23303]='h00002c1c;  wr_data_rom[23303]='h00000000;
    rd_cycle[23304] = 1'b1;  wr_cycle[23304] = 1'b0;  addr_rom[23304]='h00002c20;  wr_data_rom[23304]='h00000000;
    rd_cycle[23305] = 1'b1;  wr_cycle[23305] = 1'b0;  addr_rom[23305]='h00002c24;  wr_data_rom[23305]='h00000000;
    rd_cycle[23306] = 1'b1;  wr_cycle[23306] = 1'b0;  addr_rom[23306]='h00002c28;  wr_data_rom[23306]='h00000000;
    rd_cycle[23307] = 1'b1;  wr_cycle[23307] = 1'b0;  addr_rom[23307]='h00002c2c;  wr_data_rom[23307]='h00000000;
    rd_cycle[23308] = 1'b1;  wr_cycle[23308] = 1'b0;  addr_rom[23308]='h00002c30;  wr_data_rom[23308]='h00000000;
    rd_cycle[23309] = 1'b1;  wr_cycle[23309] = 1'b0;  addr_rom[23309]='h00002c34;  wr_data_rom[23309]='h00000000;
    rd_cycle[23310] = 1'b1;  wr_cycle[23310] = 1'b0;  addr_rom[23310]='h00002c38;  wr_data_rom[23310]='h00000000;
    rd_cycle[23311] = 1'b1;  wr_cycle[23311] = 1'b0;  addr_rom[23311]='h00002c3c;  wr_data_rom[23311]='h00000000;
    rd_cycle[23312] = 1'b1;  wr_cycle[23312] = 1'b0;  addr_rom[23312]='h00002c40;  wr_data_rom[23312]='h00000000;
    rd_cycle[23313] = 1'b1;  wr_cycle[23313] = 1'b0;  addr_rom[23313]='h00002c44;  wr_data_rom[23313]='h00000000;
    rd_cycle[23314] = 1'b1;  wr_cycle[23314] = 1'b0;  addr_rom[23314]='h00002c48;  wr_data_rom[23314]='h00000000;
    rd_cycle[23315] = 1'b1;  wr_cycle[23315] = 1'b0;  addr_rom[23315]='h00002c4c;  wr_data_rom[23315]='h00000000;
    rd_cycle[23316] = 1'b1;  wr_cycle[23316] = 1'b0;  addr_rom[23316]='h00002c50;  wr_data_rom[23316]='h00000000;
    rd_cycle[23317] = 1'b1;  wr_cycle[23317] = 1'b0;  addr_rom[23317]='h00002c54;  wr_data_rom[23317]='h00000000;
    rd_cycle[23318] = 1'b1;  wr_cycle[23318] = 1'b0;  addr_rom[23318]='h00002c58;  wr_data_rom[23318]='h00000000;
    rd_cycle[23319] = 1'b1;  wr_cycle[23319] = 1'b0;  addr_rom[23319]='h00002c5c;  wr_data_rom[23319]='h00000000;
    rd_cycle[23320] = 1'b1;  wr_cycle[23320] = 1'b0;  addr_rom[23320]='h00002c60;  wr_data_rom[23320]='h00000000;
    rd_cycle[23321] = 1'b1;  wr_cycle[23321] = 1'b0;  addr_rom[23321]='h00002c64;  wr_data_rom[23321]='h00000000;
    rd_cycle[23322] = 1'b1;  wr_cycle[23322] = 1'b0;  addr_rom[23322]='h00002c68;  wr_data_rom[23322]='h00000000;
    rd_cycle[23323] = 1'b1;  wr_cycle[23323] = 1'b0;  addr_rom[23323]='h00002c6c;  wr_data_rom[23323]='h00000000;
    rd_cycle[23324] = 1'b1;  wr_cycle[23324] = 1'b0;  addr_rom[23324]='h00002c70;  wr_data_rom[23324]='h00000000;
    rd_cycle[23325] = 1'b1;  wr_cycle[23325] = 1'b0;  addr_rom[23325]='h00002c74;  wr_data_rom[23325]='h00000000;
    rd_cycle[23326] = 1'b1;  wr_cycle[23326] = 1'b0;  addr_rom[23326]='h00002c78;  wr_data_rom[23326]='h00000000;
    rd_cycle[23327] = 1'b1;  wr_cycle[23327] = 1'b0;  addr_rom[23327]='h00002c7c;  wr_data_rom[23327]='h00000000;
    rd_cycle[23328] = 1'b1;  wr_cycle[23328] = 1'b0;  addr_rom[23328]='h00002c80;  wr_data_rom[23328]='h00000000;
    rd_cycle[23329] = 1'b1;  wr_cycle[23329] = 1'b0;  addr_rom[23329]='h00002c84;  wr_data_rom[23329]='h00000000;
    rd_cycle[23330] = 1'b1;  wr_cycle[23330] = 1'b0;  addr_rom[23330]='h00002c88;  wr_data_rom[23330]='h00000000;
    rd_cycle[23331] = 1'b1;  wr_cycle[23331] = 1'b0;  addr_rom[23331]='h00002c8c;  wr_data_rom[23331]='h00000000;
    rd_cycle[23332] = 1'b1;  wr_cycle[23332] = 1'b0;  addr_rom[23332]='h00002c90;  wr_data_rom[23332]='h00000000;
    rd_cycle[23333] = 1'b1;  wr_cycle[23333] = 1'b0;  addr_rom[23333]='h00002c94;  wr_data_rom[23333]='h00000000;
    rd_cycle[23334] = 1'b1;  wr_cycle[23334] = 1'b0;  addr_rom[23334]='h00002c98;  wr_data_rom[23334]='h00000000;
    rd_cycle[23335] = 1'b1;  wr_cycle[23335] = 1'b0;  addr_rom[23335]='h00002c9c;  wr_data_rom[23335]='h00000000;
    rd_cycle[23336] = 1'b1;  wr_cycle[23336] = 1'b0;  addr_rom[23336]='h00002ca0;  wr_data_rom[23336]='h00000000;
    rd_cycle[23337] = 1'b1;  wr_cycle[23337] = 1'b0;  addr_rom[23337]='h00002ca4;  wr_data_rom[23337]='h00000000;
    rd_cycle[23338] = 1'b1;  wr_cycle[23338] = 1'b0;  addr_rom[23338]='h00002ca8;  wr_data_rom[23338]='h00000000;
    rd_cycle[23339] = 1'b1;  wr_cycle[23339] = 1'b0;  addr_rom[23339]='h00002cac;  wr_data_rom[23339]='h00000000;
    rd_cycle[23340] = 1'b1;  wr_cycle[23340] = 1'b0;  addr_rom[23340]='h00002cb0;  wr_data_rom[23340]='h00000000;
    rd_cycle[23341] = 1'b1;  wr_cycle[23341] = 1'b0;  addr_rom[23341]='h00002cb4;  wr_data_rom[23341]='h00000000;
    rd_cycle[23342] = 1'b1;  wr_cycle[23342] = 1'b0;  addr_rom[23342]='h00002cb8;  wr_data_rom[23342]='h00000000;
    rd_cycle[23343] = 1'b1;  wr_cycle[23343] = 1'b0;  addr_rom[23343]='h00002cbc;  wr_data_rom[23343]='h00000000;
    rd_cycle[23344] = 1'b1;  wr_cycle[23344] = 1'b0;  addr_rom[23344]='h00002cc0;  wr_data_rom[23344]='h00000000;
    rd_cycle[23345] = 1'b1;  wr_cycle[23345] = 1'b0;  addr_rom[23345]='h00002cc4;  wr_data_rom[23345]='h00000000;
    rd_cycle[23346] = 1'b1;  wr_cycle[23346] = 1'b0;  addr_rom[23346]='h00002cc8;  wr_data_rom[23346]='h00000000;
    rd_cycle[23347] = 1'b1;  wr_cycle[23347] = 1'b0;  addr_rom[23347]='h00002ccc;  wr_data_rom[23347]='h00000000;
    rd_cycle[23348] = 1'b1;  wr_cycle[23348] = 1'b0;  addr_rom[23348]='h00002cd0;  wr_data_rom[23348]='h00000000;
    rd_cycle[23349] = 1'b1;  wr_cycle[23349] = 1'b0;  addr_rom[23349]='h00002cd4;  wr_data_rom[23349]='h00000000;
    rd_cycle[23350] = 1'b1;  wr_cycle[23350] = 1'b0;  addr_rom[23350]='h00002cd8;  wr_data_rom[23350]='h00000000;
    rd_cycle[23351] = 1'b1;  wr_cycle[23351] = 1'b0;  addr_rom[23351]='h00002cdc;  wr_data_rom[23351]='h00000000;
    rd_cycle[23352] = 1'b1;  wr_cycle[23352] = 1'b0;  addr_rom[23352]='h00002ce0;  wr_data_rom[23352]='h00000000;
    rd_cycle[23353] = 1'b1;  wr_cycle[23353] = 1'b0;  addr_rom[23353]='h00002ce4;  wr_data_rom[23353]='h00000000;
    rd_cycle[23354] = 1'b1;  wr_cycle[23354] = 1'b0;  addr_rom[23354]='h00002ce8;  wr_data_rom[23354]='h00000000;
    rd_cycle[23355] = 1'b1;  wr_cycle[23355] = 1'b0;  addr_rom[23355]='h00002cec;  wr_data_rom[23355]='h00000000;
    rd_cycle[23356] = 1'b1;  wr_cycle[23356] = 1'b0;  addr_rom[23356]='h00002cf0;  wr_data_rom[23356]='h00000000;
    rd_cycle[23357] = 1'b1;  wr_cycle[23357] = 1'b0;  addr_rom[23357]='h00002cf4;  wr_data_rom[23357]='h00000000;
    rd_cycle[23358] = 1'b1;  wr_cycle[23358] = 1'b0;  addr_rom[23358]='h00002cf8;  wr_data_rom[23358]='h00000000;
    rd_cycle[23359] = 1'b1;  wr_cycle[23359] = 1'b0;  addr_rom[23359]='h00002cfc;  wr_data_rom[23359]='h00000000;
    rd_cycle[23360] = 1'b1;  wr_cycle[23360] = 1'b0;  addr_rom[23360]='h00002d00;  wr_data_rom[23360]='h00000000;
    rd_cycle[23361] = 1'b1;  wr_cycle[23361] = 1'b0;  addr_rom[23361]='h00002d04;  wr_data_rom[23361]='h00000000;
    rd_cycle[23362] = 1'b1;  wr_cycle[23362] = 1'b0;  addr_rom[23362]='h00002d08;  wr_data_rom[23362]='h00000000;
    rd_cycle[23363] = 1'b1;  wr_cycle[23363] = 1'b0;  addr_rom[23363]='h00002d0c;  wr_data_rom[23363]='h00000000;
    rd_cycle[23364] = 1'b1;  wr_cycle[23364] = 1'b0;  addr_rom[23364]='h00002d10;  wr_data_rom[23364]='h00000000;
    rd_cycle[23365] = 1'b1;  wr_cycle[23365] = 1'b0;  addr_rom[23365]='h00002d14;  wr_data_rom[23365]='h00000000;
    rd_cycle[23366] = 1'b1;  wr_cycle[23366] = 1'b0;  addr_rom[23366]='h00002d18;  wr_data_rom[23366]='h00000000;
    rd_cycle[23367] = 1'b1;  wr_cycle[23367] = 1'b0;  addr_rom[23367]='h00002d1c;  wr_data_rom[23367]='h00000000;
    rd_cycle[23368] = 1'b1;  wr_cycle[23368] = 1'b0;  addr_rom[23368]='h00002d20;  wr_data_rom[23368]='h00000000;
    rd_cycle[23369] = 1'b1;  wr_cycle[23369] = 1'b0;  addr_rom[23369]='h00002d24;  wr_data_rom[23369]='h00000000;
    rd_cycle[23370] = 1'b1;  wr_cycle[23370] = 1'b0;  addr_rom[23370]='h00002d28;  wr_data_rom[23370]='h00000000;
    rd_cycle[23371] = 1'b1;  wr_cycle[23371] = 1'b0;  addr_rom[23371]='h00002d2c;  wr_data_rom[23371]='h00000000;
    rd_cycle[23372] = 1'b1;  wr_cycle[23372] = 1'b0;  addr_rom[23372]='h00002d30;  wr_data_rom[23372]='h00000000;
    rd_cycle[23373] = 1'b1;  wr_cycle[23373] = 1'b0;  addr_rom[23373]='h00002d34;  wr_data_rom[23373]='h00000000;
    rd_cycle[23374] = 1'b1;  wr_cycle[23374] = 1'b0;  addr_rom[23374]='h00002d38;  wr_data_rom[23374]='h00000000;
    rd_cycle[23375] = 1'b1;  wr_cycle[23375] = 1'b0;  addr_rom[23375]='h00002d3c;  wr_data_rom[23375]='h00000000;
    rd_cycle[23376] = 1'b1;  wr_cycle[23376] = 1'b0;  addr_rom[23376]='h00002d40;  wr_data_rom[23376]='h00000000;
    rd_cycle[23377] = 1'b1;  wr_cycle[23377] = 1'b0;  addr_rom[23377]='h00002d44;  wr_data_rom[23377]='h00000000;
    rd_cycle[23378] = 1'b1;  wr_cycle[23378] = 1'b0;  addr_rom[23378]='h00002d48;  wr_data_rom[23378]='h00000000;
    rd_cycle[23379] = 1'b1;  wr_cycle[23379] = 1'b0;  addr_rom[23379]='h00002d4c;  wr_data_rom[23379]='h00000000;
    rd_cycle[23380] = 1'b1;  wr_cycle[23380] = 1'b0;  addr_rom[23380]='h00002d50;  wr_data_rom[23380]='h00000000;
    rd_cycle[23381] = 1'b1;  wr_cycle[23381] = 1'b0;  addr_rom[23381]='h00002d54;  wr_data_rom[23381]='h00000000;
    rd_cycle[23382] = 1'b1;  wr_cycle[23382] = 1'b0;  addr_rom[23382]='h00002d58;  wr_data_rom[23382]='h00000000;
    rd_cycle[23383] = 1'b1;  wr_cycle[23383] = 1'b0;  addr_rom[23383]='h00002d5c;  wr_data_rom[23383]='h00000000;
    rd_cycle[23384] = 1'b1;  wr_cycle[23384] = 1'b0;  addr_rom[23384]='h00002d60;  wr_data_rom[23384]='h00000000;
    rd_cycle[23385] = 1'b1;  wr_cycle[23385] = 1'b0;  addr_rom[23385]='h00002d64;  wr_data_rom[23385]='h00000000;
    rd_cycle[23386] = 1'b1;  wr_cycle[23386] = 1'b0;  addr_rom[23386]='h00002d68;  wr_data_rom[23386]='h00000000;
    rd_cycle[23387] = 1'b1;  wr_cycle[23387] = 1'b0;  addr_rom[23387]='h00002d6c;  wr_data_rom[23387]='h00000000;
    rd_cycle[23388] = 1'b1;  wr_cycle[23388] = 1'b0;  addr_rom[23388]='h00002d70;  wr_data_rom[23388]='h00000000;
    rd_cycle[23389] = 1'b1;  wr_cycle[23389] = 1'b0;  addr_rom[23389]='h00002d74;  wr_data_rom[23389]='h00000000;
    rd_cycle[23390] = 1'b1;  wr_cycle[23390] = 1'b0;  addr_rom[23390]='h00002d78;  wr_data_rom[23390]='h00000000;
    rd_cycle[23391] = 1'b1;  wr_cycle[23391] = 1'b0;  addr_rom[23391]='h00002d7c;  wr_data_rom[23391]='h00000000;
    rd_cycle[23392] = 1'b1;  wr_cycle[23392] = 1'b0;  addr_rom[23392]='h00002d80;  wr_data_rom[23392]='h00000000;
    rd_cycle[23393] = 1'b1;  wr_cycle[23393] = 1'b0;  addr_rom[23393]='h00002d84;  wr_data_rom[23393]='h00000000;
    rd_cycle[23394] = 1'b1;  wr_cycle[23394] = 1'b0;  addr_rom[23394]='h00002d88;  wr_data_rom[23394]='h00000000;
    rd_cycle[23395] = 1'b1;  wr_cycle[23395] = 1'b0;  addr_rom[23395]='h00002d8c;  wr_data_rom[23395]='h00000000;
    rd_cycle[23396] = 1'b1;  wr_cycle[23396] = 1'b0;  addr_rom[23396]='h00002d90;  wr_data_rom[23396]='h00000000;
    rd_cycle[23397] = 1'b1;  wr_cycle[23397] = 1'b0;  addr_rom[23397]='h00002d94;  wr_data_rom[23397]='h00000000;
    rd_cycle[23398] = 1'b1;  wr_cycle[23398] = 1'b0;  addr_rom[23398]='h00002d98;  wr_data_rom[23398]='h00000000;
    rd_cycle[23399] = 1'b1;  wr_cycle[23399] = 1'b0;  addr_rom[23399]='h00002d9c;  wr_data_rom[23399]='h00000000;
    rd_cycle[23400] = 1'b1;  wr_cycle[23400] = 1'b0;  addr_rom[23400]='h00002da0;  wr_data_rom[23400]='h00000000;
    rd_cycle[23401] = 1'b1;  wr_cycle[23401] = 1'b0;  addr_rom[23401]='h00002da4;  wr_data_rom[23401]='h00000000;
    rd_cycle[23402] = 1'b1;  wr_cycle[23402] = 1'b0;  addr_rom[23402]='h00002da8;  wr_data_rom[23402]='h00000000;
    rd_cycle[23403] = 1'b1;  wr_cycle[23403] = 1'b0;  addr_rom[23403]='h00002dac;  wr_data_rom[23403]='h00000000;
    rd_cycle[23404] = 1'b1;  wr_cycle[23404] = 1'b0;  addr_rom[23404]='h00002db0;  wr_data_rom[23404]='h00000000;
    rd_cycle[23405] = 1'b1;  wr_cycle[23405] = 1'b0;  addr_rom[23405]='h00002db4;  wr_data_rom[23405]='h00000000;
    rd_cycle[23406] = 1'b1;  wr_cycle[23406] = 1'b0;  addr_rom[23406]='h00002db8;  wr_data_rom[23406]='h00000000;
    rd_cycle[23407] = 1'b1;  wr_cycle[23407] = 1'b0;  addr_rom[23407]='h00002dbc;  wr_data_rom[23407]='h00000000;
    rd_cycle[23408] = 1'b1;  wr_cycle[23408] = 1'b0;  addr_rom[23408]='h00002dc0;  wr_data_rom[23408]='h00000000;
    rd_cycle[23409] = 1'b1;  wr_cycle[23409] = 1'b0;  addr_rom[23409]='h00002dc4;  wr_data_rom[23409]='h00000000;
    rd_cycle[23410] = 1'b1;  wr_cycle[23410] = 1'b0;  addr_rom[23410]='h00002dc8;  wr_data_rom[23410]='h00000000;
    rd_cycle[23411] = 1'b1;  wr_cycle[23411] = 1'b0;  addr_rom[23411]='h00002dcc;  wr_data_rom[23411]='h00000000;
    rd_cycle[23412] = 1'b1;  wr_cycle[23412] = 1'b0;  addr_rom[23412]='h00002dd0;  wr_data_rom[23412]='h00000000;
    rd_cycle[23413] = 1'b1;  wr_cycle[23413] = 1'b0;  addr_rom[23413]='h00002dd4;  wr_data_rom[23413]='h00000000;
    rd_cycle[23414] = 1'b1;  wr_cycle[23414] = 1'b0;  addr_rom[23414]='h00002dd8;  wr_data_rom[23414]='h00000000;
    rd_cycle[23415] = 1'b1;  wr_cycle[23415] = 1'b0;  addr_rom[23415]='h00002ddc;  wr_data_rom[23415]='h00000000;
    rd_cycle[23416] = 1'b1;  wr_cycle[23416] = 1'b0;  addr_rom[23416]='h00002de0;  wr_data_rom[23416]='h00000000;
    rd_cycle[23417] = 1'b1;  wr_cycle[23417] = 1'b0;  addr_rom[23417]='h00002de4;  wr_data_rom[23417]='h00000000;
    rd_cycle[23418] = 1'b1;  wr_cycle[23418] = 1'b0;  addr_rom[23418]='h00002de8;  wr_data_rom[23418]='h00000000;
    rd_cycle[23419] = 1'b1;  wr_cycle[23419] = 1'b0;  addr_rom[23419]='h00002dec;  wr_data_rom[23419]='h00000000;
    rd_cycle[23420] = 1'b1;  wr_cycle[23420] = 1'b0;  addr_rom[23420]='h00002df0;  wr_data_rom[23420]='h00000000;
    rd_cycle[23421] = 1'b1;  wr_cycle[23421] = 1'b0;  addr_rom[23421]='h00002df4;  wr_data_rom[23421]='h00000000;
    rd_cycle[23422] = 1'b1;  wr_cycle[23422] = 1'b0;  addr_rom[23422]='h00002df8;  wr_data_rom[23422]='h00000000;
    rd_cycle[23423] = 1'b1;  wr_cycle[23423] = 1'b0;  addr_rom[23423]='h00002dfc;  wr_data_rom[23423]='h00000000;
    rd_cycle[23424] = 1'b1;  wr_cycle[23424] = 1'b0;  addr_rom[23424]='h00002e00;  wr_data_rom[23424]='h00000000;
    rd_cycle[23425] = 1'b1;  wr_cycle[23425] = 1'b0;  addr_rom[23425]='h00002e04;  wr_data_rom[23425]='h00000000;
    rd_cycle[23426] = 1'b1;  wr_cycle[23426] = 1'b0;  addr_rom[23426]='h00002e08;  wr_data_rom[23426]='h00000000;
    rd_cycle[23427] = 1'b1;  wr_cycle[23427] = 1'b0;  addr_rom[23427]='h00002e0c;  wr_data_rom[23427]='h00000000;
    rd_cycle[23428] = 1'b1;  wr_cycle[23428] = 1'b0;  addr_rom[23428]='h00002e10;  wr_data_rom[23428]='h00000000;
    rd_cycle[23429] = 1'b1;  wr_cycle[23429] = 1'b0;  addr_rom[23429]='h00002e14;  wr_data_rom[23429]='h00000000;
    rd_cycle[23430] = 1'b1;  wr_cycle[23430] = 1'b0;  addr_rom[23430]='h00002e18;  wr_data_rom[23430]='h00000000;
    rd_cycle[23431] = 1'b1;  wr_cycle[23431] = 1'b0;  addr_rom[23431]='h00002e1c;  wr_data_rom[23431]='h00000000;
    rd_cycle[23432] = 1'b1;  wr_cycle[23432] = 1'b0;  addr_rom[23432]='h00002e20;  wr_data_rom[23432]='h00000000;
    rd_cycle[23433] = 1'b1;  wr_cycle[23433] = 1'b0;  addr_rom[23433]='h00002e24;  wr_data_rom[23433]='h00000000;
    rd_cycle[23434] = 1'b1;  wr_cycle[23434] = 1'b0;  addr_rom[23434]='h00002e28;  wr_data_rom[23434]='h00000000;
    rd_cycle[23435] = 1'b1;  wr_cycle[23435] = 1'b0;  addr_rom[23435]='h00002e2c;  wr_data_rom[23435]='h00000000;
    rd_cycle[23436] = 1'b1;  wr_cycle[23436] = 1'b0;  addr_rom[23436]='h00002e30;  wr_data_rom[23436]='h00000000;
    rd_cycle[23437] = 1'b1;  wr_cycle[23437] = 1'b0;  addr_rom[23437]='h00002e34;  wr_data_rom[23437]='h00000000;
    rd_cycle[23438] = 1'b1;  wr_cycle[23438] = 1'b0;  addr_rom[23438]='h00002e38;  wr_data_rom[23438]='h00000000;
    rd_cycle[23439] = 1'b1;  wr_cycle[23439] = 1'b0;  addr_rom[23439]='h00002e3c;  wr_data_rom[23439]='h00000000;
    rd_cycle[23440] = 1'b1;  wr_cycle[23440] = 1'b0;  addr_rom[23440]='h00002e40;  wr_data_rom[23440]='h00000000;
    rd_cycle[23441] = 1'b1;  wr_cycle[23441] = 1'b0;  addr_rom[23441]='h00002e44;  wr_data_rom[23441]='h00000000;
    rd_cycle[23442] = 1'b1;  wr_cycle[23442] = 1'b0;  addr_rom[23442]='h00002e48;  wr_data_rom[23442]='h00000000;
    rd_cycle[23443] = 1'b1;  wr_cycle[23443] = 1'b0;  addr_rom[23443]='h00002e4c;  wr_data_rom[23443]='h00000000;
    rd_cycle[23444] = 1'b1;  wr_cycle[23444] = 1'b0;  addr_rom[23444]='h00002e50;  wr_data_rom[23444]='h00000000;
    rd_cycle[23445] = 1'b1;  wr_cycle[23445] = 1'b0;  addr_rom[23445]='h00002e54;  wr_data_rom[23445]='h00000000;
    rd_cycle[23446] = 1'b1;  wr_cycle[23446] = 1'b0;  addr_rom[23446]='h00002e58;  wr_data_rom[23446]='h00000000;
    rd_cycle[23447] = 1'b1;  wr_cycle[23447] = 1'b0;  addr_rom[23447]='h00002e5c;  wr_data_rom[23447]='h00000000;
    rd_cycle[23448] = 1'b1;  wr_cycle[23448] = 1'b0;  addr_rom[23448]='h00002e60;  wr_data_rom[23448]='h00000000;
    rd_cycle[23449] = 1'b1;  wr_cycle[23449] = 1'b0;  addr_rom[23449]='h00002e64;  wr_data_rom[23449]='h00000000;
    rd_cycle[23450] = 1'b1;  wr_cycle[23450] = 1'b0;  addr_rom[23450]='h00002e68;  wr_data_rom[23450]='h00000000;
    rd_cycle[23451] = 1'b1;  wr_cycle[23451] = 1'b0;  addr_rom[23451]='h00002e6c;  wr_data_rom[23451]='h00000000;
    rd_cycle[23452] = 1'b1;  wr_cycle[23452] = 1'b0;  addr_rom[23452]='h00002e70;  wr_data_rom[23452]='h00000000;
    rd_cycle[23453] = 1'b1;  wr_cycle[23453] = 1'b0;  addr_rom[23453]='h00002e74;  wr_data_rom[23453]='h00000000;
    rd_cycle[23454] = 1'b1;  wr_cycle[23454] = 1'b0;  addr_rom[23454]='h00002e78;  wr_data_rom[23454]='h00000000;
    rd_cycle[23455] = 1'b1;  wr_cycle[23455] = 1'b0;  addr_rom[23455]='h00002e7c;  wr_data_rom[23455]='h00000000;
    rd_cycle[23456] = 1'b1;  wr_cycle[23456] = 1'b0;  addr_rom[23456]='h00002e80;  wr_data_rom[23456]='h00000000;
    rd_cycle[23457] = 1'b1;  wr_cycle[23457] = 1'b0;  addr_rom[23457]='h00002e84;  wr_data_rom[23457]='h00000000;
    rd_cycle[23458] = 1'b1;  wr_cycle[23458] = 1'b0;  addr_rom[23458]='h00002e88;  wr_data_rom[23458]='h00000000;
    rd_cycle[23459] = 1'b1;  wr_cycle[23459] = 1'b0;  addr_rom[23459]='h00002e8c;  wr_data_rom[23459]='h00000000;
    rd_cycle[23460] = 1'b1;  wr_cycle[23460] = 1'b0;  addr_rom[23460]='h00002e90;  wr_data_rom[23460]='h00000000;
    rd_cycle[23461] = 1'b1;  wr_cycle[23461] = 1'b0;  addr_rom[23461]='h00002e94;  wr_data_rom[23461]='h00000000;
    rd_cycle[23462] = 1'b1;  wr_cycle[23462] = 1'b0;  addr_rom[23462]='h00002e98;  wr_data_rom[23462]='h00000000;
    rd_cycle[23463] = 1'b1;  wr_cycle[23463] = 1'b0;  addr_rom[23463]='h00002e9c;  wr_data_rom[23463]='h00000000;
    rd_cycle[23464] = 1'b1;  wr_cycle[23464] = 1'b0;  addr_rom[23464]='h00002ea0;  wr_data_rom[23464]='h00000000;
    rd_cycle[23465] = 1'b1;  wr_cycle[23465] = 1'b0;  addr_rom[23465]='h00002ea4;  wr_data_rom[23465]='h00000000;
    rd_cycle[23466] = 1'b1;  wr_cycle[23466] = 1'b0;  addr_rom[23466]='h00002ea8;  wr_data_rom[23466]='h00000000;
    rd_cycle[23467] = 1'b1;  wr_cycle[23467] = 1'b0;  addr_rom[23467]='h00002eac;  wr_data_rom[23467]='h00000000;
    rd_cycle[23468] = 1'b1;  wr_cycle[23468] = 1'b0;  addr_rom[23468]='h00002eb0;  wr_data_rom[23468]='h00000000;
    rd_cycle[23469] = 1'b1;  wr_cycle[23469] = 1'b0;  addr_rom[23469]='h00002eb4;  wr_data_rom[23469]='h00000000;
    rd_cycle[23470] = 1'b1;  wr_cycle[23470] = 1'b0;  addr_rom[23470]='h00002eb8;  wr_data_rom[23470]='h00000000;
    rd_cycle[23471] = 1'b1;  wr_cycle[23471] = 1'b0;  addr_rom[23471]='h00002ebc;  wr_data_rom[23471]='h00000000;
    rd_cycle[23472] = 1'b1;  wr_cycle[23472] = 1'b0;  addr_rom[23472]='h00002ec0;  wr_data_rom[23472]='h00000000;
    rd_cycle[23473] = 1'b1;  wr_cycle[23473] = 1'b0;  addr_rom[23473]='h00002ec4;  wr_data_rom[23473]='h00000000;
    rd_cycle[23474] = 1'b1;  wr_cycle[23474] = 1'b0;  addr_rom[23474]='h00002ec8;  wr_data_rom[23474]='h00000000;
    rd_cycle[23475] = 1'b1;  wr_cycle[23475] = 1'b0;  addr_rom[23475]='h00002ecc;  wr_data_rom[23475]='h00000000;
    rd_cycle[23476] = 1'b1;  wr_cycle[23476] = 1'b0;  addr_rom[23476]='h00002ed0;  wr_data_rom[23476]='h00000000;
    rd_cycle[23477] = 1'b1;  wr_cycle[23477] = 1'b0;  addr_rom[23477]='h00002ed4;  wr_data_rom[23477]='h00000000;
    rd_cycle[23478] = 1'b1;  wr_cycle[23478] = 1'b0;  addr_rom[23478]='h00002ed8;  wr_data_rom[23478]='h00000000;
    rd_cycle[23479] = 1'b1;  wr_cycle[23479] = 1'b0;  addr_rom[23479]='h00002edc;  wr_data_rom[23479]='h00000000;
    rd_cycle[23480] = 1'b1;  wr_cycle[23480] = 1'b0;  addr_rom[23480]='h00002ee0;  wr_data_rom[23480]='h00000000;
    rd_cycle[23481] = 1'b1;  wr_cycle[23481] = 1'b0;  addr_rom[23481]='h00002ee4;  wr_data_rom[23481]='h00000000;
    rd_cycle[23482] = 1'b1;  wr_cycle[23482] = 1'b0;  addr_rom[23482]='h00002ee8;  wr_data_rom[23482]='h00000000;
    rd_cycle[23483] = 1'b1;  wr_cycle[23483] = 1'b0;  addr_rom[23483]='h00002eec;  wr_data_rom[23483]='h00000000;
    rd_cycle[23484] = 1'b1;  wr_cycle[23484] = 1'b0;  addr_rom[23484]='h00002ef0;  wr_data_rom[23484]='h00000000;
    rd_cycle[23485] = 1'b1;  wr_cycle[23485] = 1'b0;  addr_rom[23485]='h00002ef4;  wr_data_rom[23485]='h00000000;
    rd_cycle[23486] = 1'b1;  wr_cycle[23486] = 1'b0;  addr_rom[23486]='h00002ef8;  wr_data_rom[23486]='h00000000;
    rd_cycle[23487] = 1'b1;  wr_cycle[23487] = 1'b0;  addr_rom[23487]='h00002efc;  wr_data_rom[23487]='h00000000;
    rd_cycle[23488] = 1'b1;  wr_cycle[23488] = 1'b0;  addr_rom[23488]='h00002f00;  wr_data_rom[23488]='h00000000;
    rd_cycle[23489] = 1'b1;  wr_cycle[23489] = 1'b0;  addr_rom[23489]='h00002f04;  wr_data_rom[23489]='h00000000;
    rd_cycle[23490] = 1'b1;  wr_cycle[23490] = 1'b0;  addr_rom[23490]='h00002f08;  wr_data_rom[23490]='h00000000;
    rd_cycle[23491] = 1'b1;  wr_cycle[23491] = 1'b0;  addr_rom[23491]='h00002f0c;  wr_data_rom[23491]='h00000000;
    rd_cycle[23492] = 1'b1;  wr_cycle[23492] = 1'b0;  addr_rom[23492]='h00002f10;  wr_data_rom[23492]='h00000000;
    rd_cycle[23493] = 1'b1;  wr_cycle[23493] = 1'b0;  addr_rom[23493]='h00002f14;  wr_data_rom[23493]='h00000000;
    rd_cycle[23494] = 1'b1;  wr_cycle[23494] = 1'b0;  addr_rom[23494]='h00002f18;  wr_data_rom[23494]='h00000000;
    rd_cycle[23495] = 1'b1;  wr_cycle[23495] = 1'b0;  addr_rom[23495]='h00002f1c;  wr_data_rom[23495]='h00000000;
    rd_cycle[23496] = 1'b1;  wr_cycle[23496] = 1'b0;  addr_rom[23496]='h00002f20;  wr_data_rom[23496]='h00000000;
    rd_cycle[23497] = 1'b1;  wr_cycle[23497] = 1'b0;  addr_rom[23497]='h00002f24;  wr_data_rom[23497]='h00000000;
    rd_cycle[23498] = 1'b1;  wr_cycle[23498] = 1'b0;  addr_rom[23498]='h00002f28;  wr_data_rom[23498]='h00000000;
    rd_cycle[23499] = 1'b1;  wr_cycle[23499] = 1'b0;  addr_rom[23499]='h00002f2c;  wr_data_rom[23499]='h00000000;
    rd_cycle[23500] = 1'b1;  wr_cycle[23500] = 1'b0;  addr_rom[23500]='h00002f30;  wr_data_rom[23500]='h00000000;
    rd_cycle[23501] = 1'b1;  wr_cycle[23501] = 1'b0;  addr_rom[23501]='h00002f34;  wr_data_rom[23501]='h00000000;
    rd_cycle[23502] = 1'b1;  wr_cycle[23502] = 1'b0;  addr_rom[23502]='h00002f38;  wr_data_rom[23502]='h00000000;
    rd_cycle[23503] = 1'b1;  wr_cycle[23503] = 1'b0;  addr_rom[23503]='h00002f3c;  wr_data_rom[23503]='h00000000;
    rd_cycle[23504] = 1'b1;  wr_cycle[23504] = 1'b0;  addr_rom[23504]='h00002f40;  wr_data_rom[23504]='h00000000;
    rd_cycle[23505] = 1'b1;  wr_cycle[23505] = 1'b0;  addr_rom[23505]='h00002f44;  wr_data_rom[23505]='h00000000;
    rd_cycle[23506] = 1'b1;  wr_cycle[23506] = 1'b0;  addr_rom[23506]='h00002f48;  wr_data_rom[23506]='h00000000;
    rd_cycle[23507] = 1'b1;  wr_cycle[23507] = 1'b0;  addr_rom[23507]='h00002f4c;  wr_data_rom[23507]='h00000000;
    rd_cycle[23508] = 1'b1;  wr_cycle[23508] = 1'b0;  addr_rom[23508]='h00002f50;  wr_data_rom[23508]='h00000000;
    rd_cycle[23509] = 1'b1;  wr_cycle[23509] = 1'b0;  addr_rom[23509]='h00002f54;  wr_data_rom[23509]='h00000000;
    rd_cycle[23510] = 1'b1;  wr_cycle[23510] = 1'b0;  addr_rom[23510]='h00002f58;  wr_data_rom[23510]='h00000000;
    rd_cycle[23511] = 1'b1;  wr_cycle[23511] = 1'b0;  addr_rom[23511]='h00002f5c;  wr_data_rom[23511]='h00000000;
    rd_cycle[23512] = 1'b1;  wr_cycle[23512] = 1'b0;  addr_rom[23512]='h00002f60;  wr_data_rom[23512]='h00000000;
    rd_cycle[23513] = 1'b1;  wr_cycle[23513] = 1'b0;  addr_rom[23513]='h00002f64;  wr_data_rom[23513]='h00000000;
    rd_cycle[23514] = 1'b1;  wr_cycle[23514] = 1'b0;  addr_rom[23514]='h00002f68;  wr_data_rom[23514]='h00000000;
    rd_cycle[23515] = 1'b1;  wr_cycle[23515] = 1'b0;  addr_rom[23515]='h00002f6c;  wr_data_rom[23515]='h00000000;
    rd_cycle[23516] = 1'b1;  wr_cycle[23516] = 1'b0;  addr_rom[23516]='h00002f70;  wr_data_rom[23516]='h00000000;
    rd_cycle[23517] = 1'b1;  wr_cycle[23517] = 1'b0;  addr_rom[23517]='h00002f74;  wr_data_rom[23517]='h00000000;
    rd_cycle[23518] = 1'b1;  wr_cycle[23518] = 1'b0;  addr_rom[23518]='h00002f78;  wr_data_rom[23518]='h00000000;
    rd_cycle[23519] = 1'b1;  wr_cycle[23519] = 1'b0;  addr_rom[23519]='h00002f7c;  wr_data_rom[23519]='h00000000;
    rd_cycle[23520] = 1'b1;  wr_cycle[23520] = 1'b0;  addr_rom[23520]='h00002f80;  wr_data_rom[23520]='h00000000;
    rd_cycle[23521] = 1'b1;  wr_cycle[23521] = 1'b0;  addr_rom[23521]='h00002f84;  wr_data_rom[23521]='h00000000;
    rd_cycle[23522] = 1'b1;  wr_cycle[23522] = 1'b0;  addr_rom[23522]='h00002f88;  wr_data_rom[23522]='h00000000;
    rd_cycle[23523] = 1'b1;  wr_cycle[23523] = 1'b0;  addr_rom[23523]='h00002f8c;  wr_data_rom[23523]='h00000000;
    rd_cycle[23524] = 1'b1;  wr_cycle[23524] = 1'b0;  addr_rom[23524]='h00002f90;  wr_data_rom[23524]='h00000000;
    rd_cycle[23525] = 1'b1;  wr_cycle[23525] = 1'b0;  addr_rom[23525]='h00002f94;  wr_data_rom[23525]='h00000000;
    rd_cycle[23526] = 1'b1;  wr_cycle[23526] = 1'b0;  addr_rom[23526]='h00002f98;  wr_data_rom[23526]='h00000000;
    rd_cycle[23527] = 1'b1;  wr_cycle[23527] = 1'b0;  addr_rom[23527]='h00002f9c;  wr_data_rom[23527]='h00000000;
    rd_cycle[23528] = 1'b1;  wr_cycle[23528] = 1'b0;  addr_rom[23528]='h00002fa0;  wr_data_rom[23528]='h00000000;
    rd_cycle[23529] = 1'b1;  wr_cycle[23529] = 1'b0;  addr_rom[23529]='h00002fa4;  wr_data_rom[23529]='h00000000;
    rd_cycle[23530] = 1'b1;  wr_cycle[23530] = 1'b0;  addr_rom[23530]='h00002fa8;  wr_data_rom[23530]='h00000000;
    rd_cycle[23531] = 1'b1;  wr_cycle[23531] = 1'b0;  addr_rom[23531]='h00002fac;  wr_data_rom[23531]='h00000000;
    rd_cycle[23532] = 1'b1;  wr_cycle[23532] = 1'b0;  addr_rom[23532]='h00002fb0;  wr_data_rom[23532]='h00000000;
    rd_cycle[23533] = 1'b1;  wr_cycle[23533] = 1'b0;  addr_rom[23533]='h00002fb4;  wr_data_rom[23533]='h00000000;
    rd_cycle[23534] = 1'b1;  wr_cycle[23534] = 1'b0;  addr_rom[23534]='h00002fb8;  wr_data_rom[23534]='h00000000;
    rd_cycle[23535] = 1'b1;  wr_cycle[23535] = 1'b0;  addr_rom[23535]='h00002fbc;  wr_data_rom[23535]='h00000000;
    rd_cycle[23536] = 1'b1;  wr_cycle[23536] = 1'b0;  addr_rom[23536]='h00002fc0;  wr_data_rom[23536]='h00000000;
    rd_cycle[23537] = 1'b1;  wr_cycle[23537] = 1'b0;  addr_rom[23537]='h00002fc4;  wr_data_rom[23537]='h00000000;
    rd_cycle[23538] = 1'b1;  wr_cycle[23538] = 1'b0;  addr_rom[23538]='h00002fc8;  wr_data_rom[23538]='h00000000;
    rd_cycle[23539] = 1'b1;  wr_cycle[23539] = 1'b0;  addr_rom[23539]='h00002fcc;  wr_data_rom[23539]='h00000000;
    rd_cycle[23540] = 1'b1;  wr_cycle[23540] = 1'b0;  addr_rom[23540]='h00002fd0;  wr_data_rom[23540]='h00000000;
    rd_cycle[23541] = 1'b1;  wr_cycle[23541] = 1'b0;  addr_rom[23541]='h00002fd4;  wr_data_rom[23541]='h00000000;
    rd_cycle[23542] = 1'b1;  wr_cycle[23542] = 1'b0;  addr_rom[23542]='h00002fd8;  wr_data_rom[23542]='h00000000;
    rd_cycle[23543] = 1'b1;  wr_cycle[23543] = 1'b0;  addr_rom[23543]='h00002fdc;  wr_data_rom[23543]='h00000000;
    rd_cycle[23544] = 1'b1;  wr_cycle[23544] = 1'b0;  addr_rom[23544]='h00002fe0;  wr_data_rom[23544]='h00000000;
    rd_cycle[23545] = 1'b1;  wr_cycle[23545] = 1'b0;  addr_rom[23545]='h00002fe4;  wr_data_rom[23545]='h00000000;
    rd_cycle[23546] = 1'b1;  wr_cycle[23546] = 1'b0;  addr_rom[23546]='h00002fe8;  wr_data_rom[23546]='h00000000;
    rd_cycle[23547] = 1'b1;  wr_cycle[23547] = 1'b0;  addr_rom[23547]='h00002fec;  wr_data_rom[23547]='h00000000;
    rd_cycle[23548] = 1'b1;  wr_cycle[23548] = 1'b0;  addr_rom[23548]='h00002ff0;  wr_data_rom[23548]='h00000000;
    rd_cycle[23549] = 1'b1;  wr_cycle[23549] = 1'b0;  addr_rom[23549]='h00002ff4;  wr_data_rom[23549]='h00000000;
    rd_cycle[23550] = 1'b1;  wr_cycle[23550] = 1'b0;  addr_rom[23550]='h00002ff8;  wr_data_rom[23550]='h00000000;
    rd_cycle[23551] = 1'b1;  wr_cycle[23551] = 1'b0;  addr_rom[23551]='h00002ffc;  wr_data_rom[23551]='h00000000;
    rd_cycle[23552] = 1'b1;  wr_cycle[23552] = 1'b0;  addr_rom[23552]='h00003000;  wr_data_rom[23552]='h00000000;
    rd_cycle[23553] = 1'b1;  wr_cycle[23553] = 1'b0;  addr_rom[23553]='h00003004;  wr_data_rom[23553]='h00000000;
    rd_cycle[23554] = 1'b1;  wr_cycle[23554] = 1'b0;  addr_rom[23554]='h00003008;  wr_data_rom[23554]='h00000000;
    rd_cycle[23555] = 1'b1;  wr_cycle[23555] = 1'b0;  addr_rom[23555]='h0000300c;  wr_data_rom[23555]='h00000000;
    rd_cycle[23556] = 1'b1;  wr_cycle[23556] = 1'b0;  addr_rom[23556]='h00003010;  wr_data_rom[23556]='h00000000;
    rd_cycle[23557] = 1'b1;  wr_cycle[23557] = 1'b0;  addr_rom[23557]='h00003014;  wr_data_rom[23557]='h00000000;
    rd_cycle[23558] = 1'b1;  wr_cycle[23558] = 1'b0;  addr_rom[23558]='h00003018;  wr_data_rom[23558]='h00000000;
    rd_cycle[23559] = 1'b1;  wr_cycle[23559] = 1'b0;  addr_rom[23559]='h0000301c;  wr_data_rom[23559]='h00000000;
    rd_cycle[23560] = 1'b1;  wr_cycle[23560] = 1'b0;  addr_rom[23560]='h00003020;  wr_data_rom[23560]='h00000000;
    rd_cycle[23561] = 1'b1;  wr_cycle[23561] = 1'b0;  addr_rom[23561]='h00003024;  wr_data_rom[23561]='h00000000;
    rd_cycle[23562] = 1'b1;  wr_cycle[23562] = 1'b0;  addr_rom[23562]='h00003028;  wr_data_rom[23562]='h00000000;
    rd_cycle[23563] = 1'b1;  wr_cycle[23563] = 1'b0;  addr_rom[23563]='h0000302c;  wr_data_rom[23563]='h00000000;
    rd_cycle[23564] = 1'b1;  wr_cycle[23564] = 1'b0;  addr_rom[23564]='h00003030;  wr_data_rom[23564]='h00000000;
    rd_cycle[23565] = 1'b1;  wr_cycle[23565] = 1'b0;  addr_rom[23565]='h00003034;  wr_data_rom[23565]='h00000000;
    rd_cycle[23566] = 1'b1;  wr_cycle[23566] = 1'b0;  addr_rom[23566]='h00003038;  wr_data_rom[23566]='h00000000;
    rd_cycle[23567] = 1'b1;  wr_cycle[23567] = 1'b0;  addr_rom[23567]='h0000303c;  wr_data_rom[23567]='h00000000;
    rd_cycle[23568] = 1'b1;  wr_cycle[23568] = 1'b0;  addr_rom[23568]='h00003040;  wr_data_rom[23568]='h00000000;
    rd_cycle[23569] = 1'b1;  wr_cycle[23569] = 1'b0;  addr_rom[23569]='h00003044;  wr_data_rom[23569]='h00000000;
    rd_cycle[23570] = 1'b1;  wr_cycle[23570] = 1'b0;  addr_rom[23570]='h00003048;  wr_data_rom[23570]='h00000000;
    rd_cycle[23571] = 1'b1;  wr_cycle[23571] = 1'b0;  addr_rom[23571]='h0000304c;  wr_data_rom[23571]='h00000000;
    rd_cycle[23572] = 1'b1;  wr_cycle[23572] = 1'b0;  addr_rom[23572]='h00003050;  wr_data_rom[23572]='h00000000;
    rd_cycle[23573] = 1'b1;  wr_cycle[23573] = 1'b0;  addr_rom[23573]='h00003054;  wr_data_rom[23573]='h00000000;
    rd_cycle[23574] = 1'b1;  wr_cycle[23574] = 1'b0;  addr_rom[23574]='h00003058;  wr_data_rom[23574]='h00000000;
    rd_cycle[23575] = 1'b1;  wr_cycle[23575] = 1'b0;  addr_rom[23575]='h0000305c;  wr_data_rom[23575]='h00000000;
    rd_cycle[23576] = 1'b1;  wr_cycle[23576] = 1'b0;  addr_rom[23576]='h00003060;  wr_data_rom[23576]='h00000000;
    rd_cycle[23577] = 1'b1;  wr_cycle[23577] = 1'b0;  addr_rom[23577]='h00003064;  wr_data_rom[23577]='h00000000;
    rd_cycle[23578] = 1'b1;  wr_cycle[23578] = 1'b0;  addr_rom[23578]='h00003068;  wr_data_rom[23578]='h00000000;
    rd_cycle[23579] = 1'b1;  wr_cycle[23579] = 1'b0;  addr_rom[23579]='h0000306c;  wr_data_rom[23579]='h00000000;
    rd_cycle[23580] = 1'b1;  wr_cycle[23580] = 1'b0;  addr_rom[23580]='h00003070;  wr_data_rom[23580]='h00000000;
    rd_cycle[23581] = 1'b1;  wr_cycle[23581] = 1'b0;  addr_rom[23581]='h00003074;  wr_data_rom[23581]='h00000000;
    rd_cycle[23582] = 1'b1;  wr_cycle[23582] = 1'b0;  addr_rom[23582]='h00003078;  wr_data_rom[23582]='h00000000;
    rd_cycle[23583] = 1'b1;  wr_cycle[23583] = 1'b0;  addr_rom[23583]='h0000307c;  wr_data_rom[23583]='h00000000;
    rd_cycle[23584] = 1'b1;  wr_cycle[23584] = 1'b0;  addr_rom[23584]='h00003080;  wr_data_rom[23584]='h00000000;
    rd_cycle[23585] = 1'b1;  wr_cycle[23585] = 1'b0;  addr_rom[23585]='h00003084;  wr_data_rom[23585]='h00000000;
    rd_cycle[23586] = 1'b1;  wr_cycle[23586] = 1'b0;  addr_rom[23586]='h00003088;  wr_data_rom[23586]='h00000000;
    rd_cycle[23587] = 1'b1;  wr_cycle[23587] = 1'b0;  addr_rom[23587]='h0000308c;  wr_data_rom[23587]='h00000000;
    rd_cycle[23588] = 1'b1;  wr_cycle[23588] = 1'b0;  addr_rom[23588]='h00003090;  wr_data_rom[23588]='h00000000;
    rd_cycle[23589] = 1'b1;  wr_cycle[23589] = 1'b0;  addr_rom[23589]='h00003094;  wr_data_rom[23589]='h00000000;
    rd_cycle[23590] = 1'b1;  wr_cycle[23590] = 1'b0;  addr_rom[23590]='h00003098;  wr_data_rom[23590]='h00000000;
    rd_cycle[23591] = 1'b1;  wr_cycle[23591] = 1'b0;  addr_rom[23591]='h0000309c;  wr_data_rom[23591]='h00000000;
    rd_cycle[23592] = 1'b1;  wr_cycle[23592] = 1'b0;  addr_rom[23592]='h000030a0;  wr_data_rom[23592]='h00000000;
    rd_cycle[23593] = 1'b1;  wr_cycle[23593] = 1'b0;  addr_rom[23593]='h000030a4;  wr_data_rom[23593]='h00000000;
    rd_cycle[23594] = 1'b1;  wr_cycle[23594] = 1'b0;  addr_rom[23594]='h000030a8;  wr_data_rom[23594]='h00000000;
    rd_cycle[23595] = 1'b1;  wr_cycle[23595] = 1'b0;  addr_rom[23595]='h000030ac;  wr_data_rom[23595]='h00000000;
    rd_cycle[23596] = 1'b1;  wr_cycle[23596] = 1'b0;  addr_rom[23596]='h000030b0;  wr_data_rom[23596]='h00000000;
    rd_cycle[23597] = 1'b1;  wr_cycle[23597] = 1'b0;  addr_rom[23597]='h000030b4;  wr_data_rom[23597]='h00000000;
    rd_cycle[23598] = 1'b1;  wr_cycle[23598] = 1'b0;  addr_rom[23598]='h000030b8;  wr_data_rom[23598]='h00000000;
    rd_cycle[23599] = 1'b1;  wr_cycle[23599] = 1'b0;  addr_rom[23599]='h000030bc;  wr_data_rom[23599]='h00000000;
    rd_cycle[23600] = 1'b1;  wr_cycle[23600] = 1'b0;  addr_rom[23600]='h000030c0;  wr_data_rom[23600]='h00000000;
    rd_cycle[23601] = 1'b1;  wr_cycle[23601] = 1'b0;  addr_rom[23601]='h000030c4;  wr_data_rom[23601]='h00000000;
    rd_cycle[23602] = 1'b1;  wr_cycle[23602] = 1'b0;  addr_rom[23602]='h000030c8;  wr_data_rom[23602]='h00000000;
    rd_cycle[23603] = 1'b1;  wr_cycle[23603] = 1'b0;  addr_rom[23603]='h000030cc;  wr_data_rom[23603]='h00000000;
    rd_cycle[23604] = 1'b1;  wr_cycle[23604] = 1'b0;  addr_rom[23604]='h000030d0;  wr_data_rom[23604]='h00000000;
    rd_cycle[23605] = 1'b1;  wr_cycle[23605] = 1'b0;  addr_rom[23605]='h000030d4;  wr_data_rom[23605]='h00000000;
    rd_cycle[23606] = 1'b1;  wr_cycle[23606] = 1'b0;  addr_rom[23606]='h000030d8;  wr_data_rom[23606]='h00000000;
    rd_cycle[23607] = 1'b1;  wr_cycle[23607] = 1'b0;  addr_rom[23607]='h000030dc;  wr_data_rom[23607]='h00000000;
    rd_cycle[23608] = 1'b1;  wr_cycle[23608] = 1'b0;  addr_rom[23608]='h000030e0;  wr_data_rom[23608]='h00000000;
    rd_cycle[23609] = 1'b1;  wr_cycle[23609] = 1'b0;  addr_rom[23609]='h000030e4;  wr_data_rom[23609]='h00000000;
    rd_cycle[23610] = 1'b1;  wr_cycle[23610] = 1'b0;  addr_rom[23610]='h000030e8;  wr_data_rom[23610]='h00000000;
    rd_cycle[23611] = 1'b1;  wr_cycle[23611] = 1'b0;  addr_rom[23611]='h000030ec;  wr_data_rom[23611]='h00000000;
    rd_cycle[23612] = 1'b1;  wr_cycle[23612] = 1'b0;  addr_rom[23612]='h000030f0;  wr_data_rom[23612]='h00000000;
    rd_cycle[23613] = 1'b1;  wr_cycle[23613] = 1'b0;  addr_rom[23613]='h000030f4;  wr_data_rom[23613]='h00000000;
    rd_cycle[23614] = 1'b1;  wr_cycle[23614] = 1'b0;  addr_rom[23614]='h000030f8;  wr_data_rom[23614]='h00000000;
    rd_cycle[23615] = 1'b1;  wr_cycle[23615] = 1'b0;  addr_rom[23615]='h000030fc;  wr_data_rom[23615]='h00000000;
    rd_cycle[23616] = 1'b1;  wr_cycle[23616] = 1'b0;  addr_rom[23616]='h00003100;  wr_data_rom[23616]='h00000000;
    rd_cycle[23617] = 1'b1;  wr_cycle[23617] = 1'b0;  addr_rom[23617]='h00003104;  wr_data_rom[23617]='h00000000;
    rd_cycle[23618] = 1'b1;  wr_cycle[23618] = 1'b0;  addr_rom[23618]='h00003108;  wr_data_rom[23618]='h00000000;
    rd_cycle[23619] = 1'b1;  wr_cycle[23619] = 1'b0;  addr_rom[23619]='h0000310c;  wr_data_rom[23619]='h00000000;
    rd_cycle[23620] = 1'b1;  wr_cycle[23620] = 1'b0;  addr_rom[23620]='h00003110;  wr_data_rom[23620]='h00000000;
    rd_cycle[23621] = 1'b1;  wr_cycle[23621] = 1'b0;  addr_rom[23621]='h00003114;  wr_data_rom[23621]='h00000000;
    rd_cycle[23622] = 1'b1;  wr_cycle[23622] = 1'b0;  addr_rom[23622]='h00003118;  wr_data_rom[23622]='h00000000;
    rd_cycle[23623] = 1'b1;  wr_cycle[23623] = 1'b0;  addr_rom[23623]='h0000311c;  wr_data_rom[23623]='h00000000;
    rd_cycle[23624] = 1'b1;  wr_cycle[23624] = 1'b0;  addr_rom[23624]='h00003120;  wr_data_rom[23624]='h00000000;
    rd_cycle[23625] = 1'b1;  wr_cycle[23625] = 1'b0;  addr_rom[23625]='h00003124;  wr_data_rom[23625]='h00000000;
    rd_cycle[23626] = 1'b1;  wr_cycle[23626] = 1'b0;  addr_rom[23626]='h00003128;  wr_data_rom[23626]='h00000000;
    rd_cycle[23627] = 1'b1;  wr_cycle[23627] = 1'b0;  addr_rom[23627]='h0000312c;  wr_data_rom[23627]='h00000000;
    rd_cycle[23628] = 1'b1;  wr_cycle[23628] = 1'b0;  addr_rom[23628]='h00003130;  wr_data_rom[23628]='h00000000;
    rd_cycle[23629] = 1'b1;  wr_cycle[23629] = 1'b0;  addr_rom[23629]='h00003134;  wr_data_rom[23629]='h00000000;
    rd_cycle[23630] = 1'b1;  wr_cycle[23630] = 1'b0;  addr_rom[23630]='h00003138;  wr_data_rom[23630]='h00000000;
    rd_cycle[23631] = 1'b1;  wr_cycle[23631] = 1'b0;  addr_rom[23631]='h0000313c;  wr_data_rom[23631]='h00000000;
    rd_cycle[23632] = 1'b1;  wr_cycle[23632] = 1'b0;  addr_rom[23632]='h00003140;  wr_data_rom[23632]='h00000000;
    rd_cycle[23633] = 1'b1;  wr_cycle[23633] = 1'b0;  addr_rom[23633]='h00003144;  wr_data_rom[23633]='h00000000;
    rd_cycle[23634] = 1'b1;  wr_cycle[23634] = 1'b0;  addr_rom[23634]='h00003148;  wr_data_rom[23634]='h00000000;
    rd_cycle[23635] = 1'b1;  wr_cycle[23635] = 1'b0;  addr_rom[23635]='h0000314c;  wr_data_rom[23635]='h00000000;
    rd_cycle[23636] = 1'b1;  wr_cycle[23636] = 1'b0;  addr_rom[23636]='h00003150;  wr_data_rom[23636]='h00000000;
    rd_cycle[23637] = 1'b1;  wr_cycle[23637] = 1'b0;  addr_rom[23637]='h00003154;  wr_data_rom[23637]='h00000000;
    rd_cycle[23638] = 1'b1;  wr_cycle[23638] = 1'b0;  addr_rom[23638]='h00003158;  wr_data_rom[23638]='h00000000;
    rd_cycle[23639] = 1'b1;  wr_cycle[23639] = 1'b0;  addr_rom[23639]='h0000315c;  wr_data_rom[23639]='h00000000;
    rd_cycle[23640] = 1'b1;  wr_cycle[23640] = 1'b0;  addr_rom[23640]='h00003160;  wr_data_rom[23640]='h00000000;
    rd_cycle[23641] = 1'b1;  wr_cycle[23641] = 1'b0;  addr_rom[23641]='h00003164;  wr_data_rom[23641]='h00000000;
    rd_cycle[23642] = 1'b1;  wr_cycle[23642] = 1'b0;  addr_rom[23642]='h00003168;  wr_data_rom[23642]='h00000000;
    rd_cycle[23643] = 1'b1;  wr_cycle[23643] = 1'b0;  addr_rom[23643]='h0000316c;  wr_data_rom[23643]='h00000000;
    rd_cycle[23644] = 1'b1;  wr_cycle[23644] = 1'b0;  addr_rom[23644]='h00003170;  wr_data_rom[23644]='h00000000;
    rd_cycle[23645] = 1'b1;  wr_cycle[23645] = 1'b0;  addr_rom[23645]='h00003174;  wr_data_rom[23645]='h00000000;
    rd_cycle[23646] = 1'b1;  wr_cycle[23646] = 1'b0;  addr_rom[23646]='h00003178;  wr_data_rom[23646]='h00000000;
    rd_cycle[23647] = 1'b1;  wr_cycle[23647] = 1'b0;  addr_rom[23647]='h0000317c;  wr_data_rom[23647]='h00000000;
    rd_cycle[23648] = 1'b1;  wr_cycle[23648] = 1'b0;  addr_rom[23648]='h00003180;  wr_data_rom[23648]='h00000000;
    rd_cycle[23649] = 1'b1;  wr_cycle[23649] = 1'b0;  addr_rom[23649]='h00003184;  wr_data_rom[23649]='h00000000;
    rd_cycle[23650] = 1'b1;  wr_cycle[23650] = 1'b0;  addr_rom[23650]='h00003188;  wr_data_rom[23650]='h00000000;
    rd_cycle[23651] = 1'b1;  wr_cycle[23651] = 1'b0;  addr_rom[23651]='h0000318c;  wr_data_rom[23651]='h00000000;
    rd_cycle[23652] = 1'b1;  wr_cycle[23652] = 1'b0;  addr_rom[23652]='h00003190;  wr_data_rom[23652]='h00000000;
    rd_cycle[23653] = 1'b1;  wr_cycle[23653] = 1'b0;  addr_rom[23653]='h00003194;  wr_data_rom[23653]='h00000000;
    rd_cycle[23654] = 1'b1;  wr_cycle[23654] = 1'b0;  addr_rom[23654]='h00003198;  wr_data_rom[23654]='h00000000;
    rd_cycle[23655] = 1'b1;  wr_cycle[23655] = 1'b0;  addr_rom[23655]='h0000319c;  wr_data_rom[23655]='h00000000;
    rd_cycle[23656] = 1'b1;  wr_cycle[23656] = 1'b0;  addr_rom[23656]='h000031a0;  wr_data_rom[23656]='h00000000;
    rd_cycle[23657] = 1'b1;  wr_cycle[23657] = 1'b0;  addr_rom[23657]='h000031a4;  wr_data_rom[23657]='h00000000;
    rd_cycle[23658] = 1'b1;  wr_cycle[23658] = 1'b0;  addr_rom[23658]='h000031a8;  wr_data_rom[23658]='h00000000;
    rd_cycle[23659] = 1'b1;  wr_cycle[23659] = 1'b0;  addr_rom[23659]='h000031ac;  wr_data_rom[23659]='h00000000;
    rd_cycle[23660] = 1'b1;  wr_cycle[23660] = 1'b0;  addr_rom[23660]='h000031b0;  wr_data_rom[23660]='h00000000;
    rd_cycle[23661] = 1'b1;  wr_cycle[23661] = 1'b0;  addr_rom[23661]='h000031b4;  wr_data_rom[23661]='h00000000;
    rd_cycle[23662] = 1'b1;  wr_cycle[23662] = 1'b0;  addr_rom[23662]='h000031b8;  wr_data_rom[23662]='h00000000;
    rd_cycle[23663] = 1'b1;  wr_cycle[23663] = 1'b0;  addr_rom[23663]='h000031bc;  wr_data_rom[23663]='h00000000;
    rd_cycle[23664] = 1'b1;  wr_cycle[23664] = 1'b0;  addr_rom[23664]='h000031c0;  wr_data_rom[23664]='h00000000;
    rd_cycle[23665] = 1'b1;  wr_cycle[23665] = 1'b0;  addr_rom[23665]='h000031c4;  wr_data_rom[23665]='h00000000;
    rd_cycle[23666] = 1'b1;  wr_cycle[23666] = 1'b0;  addr_rom[23666]='h000031c8;  wr_data_rom[23666]='h00000000;
    rd_cycle[23667] = 1'b1;  wr_cycle[23667] = 1'b0;  addr_rom[23667]='h000031cc;  wr_data_rom[23667]='h00000000;
    rd_cycle[23668] = 1'b1;  wr_cycle[23668] = 1'b0;  addr_rom[23668]='h000031d0;  wr_data_rom[23668]='h00000000;
    rd_cycle[23669] = 1'b1;  wr_cycle[23669] = 1'b0;  addr_rom[23669]='h000031d4;  wr_data_rom[23669]='h00000000;
    rd_cycle[23670] = 1'b1;  wr_cycle[23670] = 1'b0;  addr_rom[23670]='h000031d8;  wr_data_rom[23670]='h00000000;
    rd_cycle[23671] = 1'b1;  wr_cycle[23671] = 1'b0;  addr_rom[23671]='h000031dc;  wr_data_rom[23671]='h00000000;
    rd_cycle[23672] = 1'b1;  wr_cycle[23672] = 1'b0;  addr_rom[23672]='h000031e0;  wr_data_rom[23672]='h00000000;
    rd_cycle[23673] = 1'b1;  wr_cycle[23673] = 1'b0;  addr_rom[23673]='h000031e4;  wr_data_rom[23673]='h00000000;
    rd_cycle[23674] = 1'b1;  wr_cycle[23674] = 1'b0;  addr_rom[23674]='h000031e8;  wr_data_rom[23674]='h00000000;
    rd_cycle[23675] = 1'b1;  wr_cycle[23675] = 1'b0;  addr_rom[23675]='h000031ec;  wr_data_rom[23675]='h00000000;
    rd_cycle[23676] = 1'b1;  wr_cycle[23676] = 1'b0;  addr_rom[23676]='h000031f0;  wr_data_rom[23676]='h00000000;
    rd_cycle[23677] = 1'b1;  wr_cycle[23677] = 1'b0;  addr_rom[23677]='h000031f4;  wr_data_rom[23677]='h00000000;
    rd_cycle[23678] = 1'b1;  wr_cycle[23678] = 1'b0;  addr_rom[23678]='h000031f8;  wr_data_rom[23678]='h00000000;
    rd_cycle[23679] = 1'b1;  wr_cycle[23679] = 1'b0;  addr_rom[23679]='h000031fc;  wr_data_rom[23679]='h00000000;
    rd_cycle[23680] = 1'b1;  wr_cycle[23680] = 1'b0;  addr_rom[23680]='h00003200;  wr_data_rom[23680]='h00000000;
    rd_cycle[23681] = 1'b1;  wr_cycle[23681] = 1'b0;  addr_rom[23681]='h00003204;  wr_data_rom[23681]='h00000000;
    rd_cycle[23682] = 1'b1;  wr_cycle[23682] = 1'b0;  addr_rom[23682]='h00003208;  wr_data_rom[23682]='h00000000;
    rd_cycle[23683] = 1'b1;  wr_cycle[23683] = 1'b0;  addr_rom[23683]='h0000320c;  wr_data_rom[23683]='h00000000;
    rd_cycle[23684] = 1'b1;  wr_cycle[23684] = 1'b0;  addr_rom[23684]='h00003210;  wr_data_rom[23684]='h00000000;
    rd_cycle[23685] = 1'b1;  wr_cycle[23685] = 1'b0;  addr_rom[23685]='h00003214;  wr_data_rom[23685]='h00000000;
    rd_cycle[23686] = 1'b1;  wr_cycle[23686] = 1'b0;  addr_rom[23686]='h00003218;  wr_data_rom[23686]='h00000000;
    rd_cycle[23687] = 1'b1;  wr_cycle[23687] = 1'b0;  addr_rom[23687]='h0000321c;  wr_data_rom[23687]='h00000000;
    rd_cycle[23688] = 1'b1;  wr_cycle[23688] = 1'b0;  addr_rom[23688]='h00003220;  wr_data_rom[23688]='h00000000;
    rd_cycle[23689] = 1'b1;  wr_cycle[23689] = 1'b0;  addr_rom[23689]='h00003224;  wr_data_rom[23689]='h00000000;
    rd_cycle[23690] = 1'b1;  wr_cycle[23690] = 1'b0;  addr_rom[23690]='h00003228;  wr_data_rom[23690]='h00000000;
    rd_cycle[23691] = 1'b1;  wr_cycle[23691] = 1'b0;  addr_rom[23691]='h0000322c;  wr_data_rom[23691]='h00000000;
    rd_cycle[23692] = 1'b1;  wr_cycle[23692] = 1'b0;  addr_rom[23692]='h00003230;  wr_data_rom[23692]='h00000000;
    rd_cycle[23693] = 1'b1;  wr_cycle[23693] = 1'b0;  addr_rom[23693]='h00003234;  wr_data_rom[23693]='h00000000;
    rd_cycle[23694] = 1'b1;  wr_cycle[23694] = 1'b0;  addr_rom[23694]='h00003238;  wr_data_rom[23694]='h00000000;
    rd_cycle[23695] = 1'b1;  wr_cycle[23695] = 1'b0;  addr_rom[23695]='h0000323c;  wr_data_rom[23695]='h00000000;
    rd_cycle[23696] = 1'b1;  wr_cycle[23696] = 1'b0;  addr_rom[23696]='h00003240;  wr_data_rom[23696]='h00000000;
    rd_cycle[23697] = 1'b1;  wr_cycle[23697] = 1'b0;  addr_rom[23697]='h00003244;  wr_data_rom[23697]='h00000000;
    rd_cycle[23698] = 1'b1;  wr_cycle[23698] = 1'b0;  addr_rom[23698]='h00003248;  wr_data_rom[23698]='h00000000;
    rd_cycle[23699] = 1'b1;  wr_cycle[23699] = 1'b0;  addr_rom[23699]='h0000324c;  wr_data_rom[23699]='h00000000;
    rd_cycle[23700] = 1'b1;  wr_cycle[23700] = 1'b0;  addr_rom[23700]='h00003250;  wr_data_rom[23700]='h00000000;
    rd_cycle[23701] = 1'b1;  wr_cycle[23701] = 1'b0;  addr_rom[23701]='h00003254;  wr_data_rom[23701]='h00000000;
    rd_cycle[23702] = 1'b1;  wr_cycle[23702] = 1'b0;  addr_rom[23702]='h00003258;  wr_data_rom[23702]='h00000000;
    rd_cycle[23703] = 1'b1;  wr_cycle[23703] = 1'b0;  addr_rom[23703]='h0000325c;  wr_data_rom[23703]='h00000000;
    rd_cycle[23704] = 1'b1;  wr_cycle[23704] = 1'b0;  addr_rom[23704]='h00003260;  wr_data_rom[23704]='h00000000;
    rd_cycle[23705] = 1'b1;  wr_cycle[23705] = 1'b0;  addr_rom[23705]='h00003264;  wr_data_rom[23705]='h00000000;
    rd_cycle[23706] = 1'b1;  wr_cycle[23706] = 1'b0;  addr_rom[23706]='h00003268;  wr_data_rom[23706]='h00000000;
    rd_cycle[23707] = 1'b1;  wr_cycle[23707] = 1'b0;  addr_rom[23707]='h0000326c;  wr_data_rom[23707]='h00000000;
    rd_cycle[23708] = 1'b1;  wr_cycle[23708] = 1'b0;  addr_rom[23708]='h00003270;  wr_data_rom[23708]='h00000000;
    rd_cycle[23709] = 1'b1;  wr_cycle[23709] = 1'b0;  addr_rom[23709]='h00003274;  wr_data_rom[23709]='h00000000;
    rd_cycle[23710] = 1'b1;  wr_cycle[23710] = 1'b0;  addr_rom[23710]='h00003278;  wr_data_rom[23710]='h00000000;
    rd_cycle[23711] = 1'b1;  wr_cycle[23711] = 1'b0;  addr_rom[23711]='h0000327c;  wr_data_rom[23711]='h00000000;
    rd_cycle[23712] = 1'b1;  wr_cycle[23712] = 1'b0;  addr_rom[23712]='h00003280;  wr_data_rom[23712]='h00000000;
    rd_cycle[23713] = 1'b1;  wr_cycle[23713] = 1'b0;  addr_rom[23713]='h00003284;  wr_data_rom[23713]='h00000000;
    rd_cycle[23714] = 1'b1;  wr_cycle[23714] = 1'b0;  addr_rom[23714]='h00003288;  wr_data_rom[23714]='h00000000;
    rd_cycle[23715] = 1'b1;  wr_cycle[23715] = 1'b0;  addr_rom[23715]='h0000328c;  wr_data_rom[23715]='h00000000;
    rd_cycle[23716] = 1'b1;  wr_cycle[23716] = 1'b0;  addr_rom[23716]='h00003290;  wr_data_rom[23716]='h00000000;
    rd_cycle[23717] = 1'b1;  wr_cycle[23717] = 1'b0;  addr_rom[23717]='h00003294;  wr_data_rom[23717]='h00000000;
    rd_cycle[23718] = 1'b1;  wr_cycle[23718] = 1'b0;  addr_rom[23718]='h00003298;  wr_data_rom[23718]='h00000000;
    rd_cycle[23719] = 1'b1;  wr_cycle[23719] = 1'b0;  addr_rom[23719]='h0000329c;  wr_data_rom[23719]='h00000000;
    rd_cycle[23720] = 1'b1;  wr_cycle[23720] = 1'b0;  addr_rom[23720]='h000032a0;  wr_data_rom[23720]='h00000000;
    rd_cycle[23721] = 1'b1;  wr_cycle[23721] = 1'b0;  addr_rom[23721]='h000032a4;  wr_data_rom[23721]='h00000000;
    rd_cycle[23722] = 1'b1;  wr_cycle[23722] = 1'b0;  addr_rom[23722]='h000032a8;  wr_data_rom[23722]='h00000000;
    rd_cycle[23723] = 1'b1;  wr_cycle[23723] = 1'b0;  addr_rom[23723]='h000032ac;  wr_data_rom[23723]='h00000000;
    rd_cycle[23724] = 1'b1;  wr_cycle[23724] = 1'b0;  addr_rom[23724]='h000032b0;  wr_data_rom[23724]='h00000000;
    rd_cycle[23725] = 1'b1;  wr_cycle[23725] = 1'b0;  addr_rom[23725]='h000032b4;  wr_data_rom[23725]='h00000000;
    rd_cycle[23726] = 1'b1;  wr_cycle[23726] = 1'b0;  addr_rom[23726]='h000032b8;  wr_data_rom[23726]='h00000000;
    rd_cycle[23727] = 1'b1;  wr_cycle[23727] = 1'b0;  addr_rom[23727]='h000032bc;  wr_data_rom[23727]='h00000000;
    rd_cycle[23728] = 1'b1;  wr_cycle[23728] = 1'b0;  addr_rom[23728]='h000032c0;  wr_data_rom[23728]='h00000000;
    rd_cycle[23729] = 1'b1;  wr_cycle[23729] = 1'b0;  addr_rom[23729]='h000032c4;  wr_data_rom[23729]='h00000000;
    rd_cycle[23730] = 1'b1;  wr_cycle[23730] = 1'b0;  addr_rom[23730]='h000032c8;  wr_data_rom[23730]='h00000000;
    rd_cycle[23731] = 1'b1;  wr_cycle[23731] = 1'b0;  addr_rom[23731]='h000032cc;  wr_data_rom[23731]='h00000000;
    rd_cycle[23732] = 1'b1;  wr_cycle[23732] = 1'b0;  addr_rom[23732]='h000032d0;  wr_data_rom[23732]='h00000000;
    rd_cycle[23733] = 1'b1;  wr_cycle[23733] = 1'b0;  addr_rom[23733]='h000032d4;  wr_data_rom[23733]='h00000000;
    rd_cycle[23734] = 1'b1;  wr_cycle[23734] = 1'b0;  addr_rom[23734]='h000032d8;  wr_data_rom[23734]='h00000000;
    rd_cycle[23735] = 1'b1;  wr_cycle[23735] = 1'b0;  addr_rom[23735]='h000032dc;  wr_data_rom[23735]='h00000000;
    rd_cycle[23736] = 1'b1;  wr_cycle[23736] = 1'b0;  addr_rom[23736]='h000032e0;  wr_data_rom[23736]='h00000000;
    rd_cycle[23737] = 1'b1;  wr_cycle[23737] = 1'b0;  addr_rom[23737]='h000032e4;  wr_data_rom[23737]='h00000000;
    rd_cycle[23738] = 1'b1;  wr_cycle[23738] = 1'b0;  addr_rom[23738]='h000032e8;  wr_data_rom[23738]='h00000000;
    rd_cycle[23739] = 1'b1;  wr_cycle[23739] = 1'b0;  addr_rom[23739]='h000032ec;  wr_data_rom[23739]='h00000000;
    rd_cycle[23740] = 1'b1;  wr_cycle[23740] = 1'b0;  addr_rom[23740]='h000032f0;  wr_data_rom[23740]='h00000000;
    rd_cycle[23741] = 1'b1;  wr_cycle[23741] = 1'b0;  addr_rom[23741]='h000032f4;  wr_data_rom[23741]='h00000000;
    rd_cycle[23742] = 1'b1;  wr_cycle[23742] = 1'b0;  addr_rom[23742]='h000032f8;  wr_data_rom[23742]='h00000000;
    rd_cycle[23743] = 1'b1;  wr_cycle[23743] = 1'b0;  addr_rom[23743]='h000032fc;  wr_data_rom[23743]='h00000000;
    rd_cycle[23744] = 1'b1;  wr_cycle[23744] = 1'b0;  addr_rom[23744]='h00003300;  wr_data_rom[23744]='h00000000;
    rd_cycle[23745] = 1'b1;  wr_cycle[23745] = 1'b0;  addr_rom[23745]='h00003304;  wr_data_rom[23745]='h00000000;
    rd_cycle[23746] = 1'b1;  wr_cycle[23746] = 1'b0;  addr_rom[23746]='h00003308;  wr_data_rom[23746]='h00000000;
    rd_cycle[23747] = 1'b1;  wr_cycle[23747] = 1'b0;  addr_rom[23747]='h0000330c;  wr_data_rom[23747]='h00000000;
    rd_cycle[23748] = 1'b1;  wr_cycle[23748] = 1'b0;  addr_rom[23748]='h00003310;  wr_data_rom[23748]='h00000000;
    rd_cycle[23749] = 1'b1;  wr_cycle[23749] = 1'b0;  addr_rom[23749]='h00003314;  wr_data_rom[23749]='h00000000;
    rd_cycle[23750] = 1'b1;  wr_cycle[23750] = 1'b0;  addr_rom[23750]='h00003318;  wr_data_rom[23750]='h00000000;
    rd_cycle[23751] = 1'b1;  wr_cycle[23751] = 1'b0;  addr_rom[23751]='h0000331c;  wr_data_rom[23751]='h00000000;
    rd_cycle[23752] = 1'b1;  wr_cycle[23752] = 1'b0;  addr_rom[23752]='h00003320;  wr_data_rom[23752]='h00000000;
    rd_cycle[23753] = 1'b1;  wr_cycle[23753] = 1'b0;  addr_rom[23753]='h00003324;  wr_data_rom[23753]='h00000000;
    rd_cycle[23754] = 1'b1;  wr_cycle[23754] = 1'b0;  addr_rom[23754]='h00003328;  wr_data_rom[23754]='h00000000;
    rd_cycle[23755] = 1'b1;  wr_cycle[23755] = 1'b0;  addr_rom[23755]='h0000332c;  wr_data_rom[23755]='h00000000;
    rd_cycle[23756] = 1'b1;  wr_cycle[23756] = 1'b0;  addr_rom[23756]='h00003330;  wr_data_rom[23756]='h00000000;
    rd_cycle[23757] = 1'b1;  wr_cycle[23757] = 1'b0;  addr_rom[23757]='h00003334;  wr_data_rom[23757]='h00000000;
    rd_cycle[23758] = 1'b1;  wr_cycle[23758] = 1'b0;  addr_rom[23758]='h00003338;  wr_data_rom[23758]='h00000000;
    rd_cycle[23759] = 1'b1;  wr_cycle[23759] = 1'b0;  addr_rom[23759]='h0000333c;  wr_data_rom[23759]='h00000000;
    rd_cycle[23760] = 1'b1;  wr_cycle[23760] = 1'b0;  addr_rom[23760]='h00003340;  wr_data_rom[23760]='h00000000;
    rd_cycle[23761] = 1'b1;  wr_cycle[23761] = 1'b0;  addr_rom[23761]='h00003344;  wr_data_rom[23761]='h00000000;
    rd_cycle[23762] = 1'b1;  wr_cycle[23762] = 1'b0;  addr_rom[23762]='h00003348;  wr_data_rom[23762]='h00000000;
    rd_cycle[23763] = 1'b1;  wr_cycle[23763] = 1'b0;  addr_rom[23763]='h0000334c;  wr_data_rom[23763]='h00000000;
    rd_cycle[23764] = 1'b1;  wr_cycle[23764] = 1'b0;  addr_rom[23764]='h00003350;  wr_data_rom[23764]='h00000000;
    rd_cycle[23765] = 1'b1;  wr_cycle[23765] = 1'b0;  addr_rom[23765]='h00003354;  wr_data_rom[23765]='h00000000;
    rd_cycle[23766] = 1'b1;  wr_cycle[23766] = 1'b0;  addr_rom[23766]='h00003358;  wr_data_rom[23766]='h00000000;
    rd_cycle[23767] = 1'b1;  wr_cycle[23767] = 1'b0;  addr_rom[23767]='h0000335c;  wr_data_rom[23767]='h00000000;
    rd_cycle[23768] = 1'b1;  wr_cycle[23768] = 1'b0;  addr_rom[23768]='h00003360;  wr_data_rom[23768]='h00000000;
    rd_cycle[23769] = 1'b1;  wr_cycle[23769] = 1'b0;  addr_rom[23769]='h00003364;  wr_data_rom[23769]='h00000000;
    rd_cycle[23770] = 1'b1;  wr_cycle[23770] = 1'b0;  addr_rom[23770]='h00003368;  wr_data_rom[23770]='h00000000;
    rd_cycle[23771] = 1'b1;  wr_cycle[23771] = 1'b0;  addr_rom[23771]='h0000336c;  wr_data_rom[23771]='h00000000;
    rd_cycle[23772] = 1'b1;  wr_cycle[23772] = 1'b0;  addr_rom[23772]='h00003370;  wr_data_rom[23772]='h00000000;
    rd_cycle[23773] = 1'b1;  wr_cycle[23773] = 1'b0;  addr_rom[23773]='h00003374;  wr_data_rom[23773]='h00000000;
    rd_cycle[23774] = 1'b1;  wr_cycle[23774] = 1'b0;  addr_rom[23774]='h00003378;  wr_data_rom[23774]='h00000000;
    rd_cycle[23775] = 1'b1;  wr_cycle[23775] = 1'b0;  addr_rom[23775]='h0000337c;  wr_data_rom[23775]='h00000000;
    rd_cycle[23776] = 1'b1;  wr_cycle[23776] = 1'b0;  addr_rom[23776]='h00003380;  wr_data_rom[23776]='h00000000;
    rd_cycle[23777] = 1'b1;  wr_cycle[23777] = 1'b0;  addr_rom[23777]='h00003384;  wr_data_rom[23777]='h00000000;
    rd_cycle[23778] = 1'b1;  wr_cycle[23778] = 1'b0;  addr_rom[23778]='h00003388;  wr_data_rom[23778]='h00000000;
    rd_cycle[23779] = 1'b1;  wr_cycle[23779] = 1'b0;  addr_rom[23779]='h0000338c;  wr_data_rom[23779]='h00000000;
    rd_cycle[23780] = 1'b1;  wr_cycle[23780] = 1'b0;  addr_rom[23780]='h00003390;  wr_data_rom[23780]='h00000000;
    rd_cycle[23781] = 1'b1;  wr_cycle[23781] = 1'b0;  addr_rom[23781]='h00003394;  wr_data_rom[23781]='h00000000;
    rd_cycle[23782] = 1'b1;  wr_cycle[23782] = 1'b0;  addr_rom[23782]='h00003398;  wr_data_rom[23782]='h00000000;
    rd_cycle[23783] = 1'b1;  wr_cycle[23783] = 1'b0;  addr_rom[23783]='h0000339c;  wr_data_rom[23783]='h00000000;
    rd_cycle[23784] = 1'b1;  wr_cycle[23784] = 1'b0;  addr_rom[23784]='h000033a0;  wr_data_rom[23784]='h00000000;
    rd_cycle[23785] = 1'b1;  wr_cycle[23785] = 1'b0;  addr_rom[23785]='h000033a4;  wr_data_rom[23785]='h00000000;
    rd_cycle[23786] = 1'b1;  wr_cycle[23786] = 1'b0;  addr_rom[23786]='h000033a8;  wr_data_rom[23786]='h00000000;
    rd_cycle[23787] = 1'b1;  wr_cycle[23787] = 1'b0;  addr_rom[23787]='h000033ac;  wr_data_rom[23787]='h00000000;
    rd_cycle[23788] = 1'b1;  wr_cycle[23788] = 1'b0;  addr_rom[23788]='h000033b0;  wr_data_rom[23788]='h00000000;
    rd_cycle[23789] = 1'b1;  wr_cycle[23789] = 1'b0;  addr_rom[23789]='h000033b4;  wr_data_rom[23789]='h00000000;
    rd_cycle[23790] = 1'b1;  wr_cycle[23790] = 1'b0;  addr_rom[23790]='h000033b8;  wr_data_rom[23790]='h00000000;
    rd_cycle[23791] = 1'b1;  wr_cycle[23791] = 1'b0;  addr_rom[23791]='h000033bc;  wr_data_rom[23791]='h00000000;
    rd_cycle[23792] = 1'b1;  wr_cycle[23792] = 1'b0;  addr_rom[23792]='h000033c0;  wr_data_rom[23792]='h00000000;
    rd_cycle[23793] = 1'b1;  wr_cycle[23793] = 1'b0;  addr_rom[23793]='h000033c4;  wr_data_rom[23793]='h00000000;
    rd_cycle[23794] = 1'b1;  wr_cycle[23794] = 1'b0;  addr_rom[23794]='h000033c8;  wr_data_rom[23794]='h00000000;
    rd_cycle[23795] = 1'b1;  wr_cycle[23795] = 1'b0;  addr_rom[23795]='h000033cc;  wr_data_rom[23795]='h00000000;
    rd_cycle[23796] = 1'b1;  wr_cycle[23796] = 1'b0;  addr_rom[23796]='h000033d0;  wr_data_rom[23796]='h00000000;
    rd_cycle[23797] = 1'b1;  wr_cycle[23797] = 1'b0;  addr_rom[23797]='h000033d4;  wr_data_rom[23797]='h00000000;
    rd_cycle[23798] = 1'b1;  wr_cycle[23798] = 1'b0;  addr_rom[23798]='h000033d8;  wr_data_rom[23798]='h00000000;
    rd_cycle[23799] = 1'b1;  wr_cycle[23799] = 1'b0;  addr_rom[23799]='h000033dc;  wr_data_rom[23799]='h00000000;
    rd_cycle[23800] = 1'b1;  wr_cycle[23800] = 1'b0;  addr_rom[23800]='h000033e0;  wr_data_rom[23800]='h00000000;
    rd_cycle[23801] = 1'b1;  wr_cycle[23801] = 1'b0;  addr_rom[23801]='h000033e4;  wr_data_rom[23801]='h00000000;
    rd_cycle[23802] = 1'b1;  wr_cycle[23802] = 1'b0;  addr_rom[23802]='h000033e8;  wr_data_rom[23802]='h00000000;
    rd_cycle[23803] = 1'b1;  wr_cycle[23803] = 1'b0;  addr_rom[23803]='h000033ec;  wr_data_rom[23803]='h00000000;
    rd_cycle[23804] = 1'b1;  wr_cycle[23804] = 1'b0;  addr_rom[23804]='h000033f0;  wr_data_rom[23804]='h00000000;
    rd_cycle[23805] = 1'b1;  wr_cycle[23805] = 1'b0;  addr_rom[23805]='h000033f4;  wr_data_rom[23805]='h00000000;
    rd_cycle[23806] = 1'b1;  wr_cycle[23806] = 1'b0;  addr_rom[23806]='h000033f8;  wr_data_rom[23806]='h00000000;
    rd_cycle[23807] = 1'b1;  wr_cycle[23807] = 1'b0;  addr_rom[23807]='h000033fc;  wr_data_rom[23807]='h00000000;
    rd_cycle[23808] = 1'b1;  wr_cycle[23808] = 1'b0;  addr_rom[23808]='h00003400;  wr_data_rom[23808]='h00000000;
    rd_cycle[23809] = 1'b1;  wr_cycle[23809] = 1'b0;  addr_rom[23809]='h00003404;  wr_data_rom[23809]='h00000000;
    rd_cycle[23810] = 1'b1;  wr_cycle[23810] = 1'b0;  addr_rom[23810]='h00003408;  wr_data_rom[23810]='h00000000;
    rd_cycle[23811] = 1'b1;  wr_cycle[23811] = 1'b0;  addr_rom[23811]='h0000340c;  wr_data_rom[23811]='h00000000;
    rd_cycle[23812] = 1'b1;  wr_cycle[23812] = 1'b0;  addr_rom[23812]='h00003410;  wr_data_rom[23812]='h00000000;
    rd_cycle[23813] = 1'b1;  wr_cycle[23813] = 1'b0;  addr_rom[23813]='h00003414;  wr_data_rom[23813]='h00000000;
    rd_cycle[23814] = 1'b1;  wr_cycle[23814] = 1'b0;  addr_rom[23814]='h00003418;  wr_data_rom[23814]='h00000000;
    rd_cycle[23815] = 1'b1;  wr_cycle[23815] = 1'b0;  addr_rom[23815]='h0000341c;  wr_data_rom[23815]='h00000000;
    rd_cycle[23816] = 1'b1;  wr_cycle[23816] = 1'b0;  addr_rom[23816]='h00003420;  wr_data_rom[23816]='h00000000;
    rd_cycle[23817] = 1'b1;  wr_cycle[23817] = 1'b0;  addr_rom[23817]='h00003424;  wr_data_rom[23817]='h00000000;
    rd_cycle[23818] = 1'b1;  wr_cycle[23818] = 1'b0;  addr_rom[23818]='h00003428;  wr_data_rom[23818]='h00000000;
    rd_cycle[23819] = 1'b1;  wr_cycle[23819] = 1'b0;  addr_rom[23819]='h0000342c;  wr_data_rom[23819]='h00000000;
    rd_cycle[23820] = 1'b1;  wr_cycle[23820] = 1'b0;  addr_rom[23820]='h00003430;  wr_data_rom[23820]='h00000000;
    rd_cycle[23821] = 1'b1;  wr_cycle[23821] = 1'b0;  addr_rom[23821]='h00003434;  wr_data_rom[23821]='h00000000;
    rd_cycle[23822] = 1'b1;  wr_cycle[23822] = 1'b0;  addr_rom[23822]='h00003438;  wr_data_rom[23822]='h00000000;
    rd_cycle[23823] = 1'b1;  wr_cycle[23823] = 1'b0;  addr_rom[23823]='h0000343c;  wr_data_rom[23823]='h00000000;
    rd_cycle[23824] = 1'b1;  wr_cycle[23824] = 1'b0;  addr_rom[23824]='h00003440;  wr_data_rom[23824]='h00000000;
    rd_cycle[23825] = 1'b1;  wr_cycle[23825] = 1'b0;  addr_rom[23825]='h00003444;  wr_data_rom[23825]='h00000000;
    rd_cycle[23826] = 1'b1;  wr_cycle[23826] = 1'b0;  addr_rom[23826]='h00003448;  wr_data_rom[23826]='h00000000;
    rd_cycle[23827] = 1'b1;  wr_cycle[23827] = 1'b0;  addr_rom[23827]='h0000344c;  wr_data_rom[23827]='h00000000;
    rd_cycle[23828] = 1'b1;  wr_cycle[23828] = 1'b0;  addr_rom[23828]='h00003450;  wr_data_rom[23828]='h00000000;
    rd_cycle[23829] = 1'b1;  wr_cycle[23829] = 1'b0;  addr_rom[23829]='h00003454;  wr_data_rom[23829]='h00000000;
    rd_cycle[23830] = 1'b1;  wr_cycle[23830] = 1'b0;  addr_rom[23830]='h00003458;  wr_data_rom[23830]='h00000000;
    rd_cycle[23831] = 1'b1;  wr_cycle[23831] = 1'b0;  addr_rom[23831]='h0000345c;  wr_data_rom[23831]='h00000000;
    rd_cycle[23832] = 1'b1;  wr_cycle[23832] = 1'b0;  addr_rom[23832]='h00003460;  wr_data_rom[23832]='h00000000;
    rd_cycle[23833] = 1'b1;  wr_cycle[23833] = 1'b0;  addr_rom[23833]='h00003464;  wr_data_rom[23833]='h00000000;
    rd_cycle[23834] = 1'b1;  wr_cycle[23834] = 1'b0;  addr_rom[23834]='h00003468;  wr_data_rom[23834]='h00000000;
    rd_cycle[23835] = 1'b1;  wr_cycle[23835] = 1'b0;  addr_rom[23835]='h0000346c;  wr_data_rom[23835]='h00000000;
    rd_cycle[23836] = 1'b1;  wr_cycle[23836] = 1'b0;  addr_rom[23836]='h00003470;  wr_data_rom[23836]='h00000000;
    rd_cycle[23837] = 1'b1;  wr_cycle[23837] = 1'b0;  addr_rom[23837]='h00003474;  wr_data_rom[23837]='h00000000;
    rd_cycle[23838] = 1'b1;  wr_cycle[23838] = 1'b0;  addr_rom[23838]='h00003478;  wr_data_rom[23838]='h00000000;
    rd_cycle[23839] = 1'b1;  wr_cycle[23839] = 1'b0;  addr_rom[23839]='h0000347c;  wr_data_rom[23839]='h00000000;
    rd_cycle[23840] = 1'b1;  wr_cycle[23840] = 1'b0;  addr_rom[23840]='h00003480;  wr_data_rom[23840]='h00000000;
    rd_cycle[23841] = 1'b1;  wr_cycle[23841] = 1'b0;  addr_rom[23841]='h00003484;  wr_data_rom[23841]='h00000000;
    rd_cycle[23842] = 1'b1;  wr_cycle[23842] = 1'b0;  addr_rom[23842]='h00003488;  wr_data_rom[23842]='h00000000;
    rd_cycle[23843] = 1'b1;  wr_cycle[23843] = 1'b0;  addr_rom[23843]='h0000348c;  wr_data_rom[23843]='h00000000;
    rd_cycle[23844] = 1'b1;  wr_cycle[23844] = 1'b0;  addr_rom[23844]='h00003490;  wr_data_rom[23844]='h00000000;
    rd_cycle[23845] = 1'b1;  wr_cycle[23845] = 1'b0;  addr_rom[23845]='h00003494;  wr_data_rom[23845]='h00000000;
    rd_cycle[23846] = 1'b1;  wr_cycle[23846] = 1'b0;  addr_rom[23846]='h00003498;  wr_data_rom[23846]='h00000000;
    rd_cycle[23847] = 1'b1;  wr_cycle[23847] = 1'b0;  addr_rom[23847]='h0000349c;  wr_data_rom[23847]='h00000000;
    rd_cycle[23848] = 1'b1;  wr_cycle[23848] = 1'b0;  addr_rom[23848]='h000034a0;  wr_data_rom[23848]='h00000000;
    rd_cycle[23849] = 1'b1;  wr_cycle[23849] = 1'b0;  addr_rom[23849]='h000034a4;  wr_data_rom[23849]='h00000000;
    rd_cycle[23850] = 1'b1;  wr_cycle[23850] = 1'b0;  addr_rom[23850]='h000034a8;  wr_data_rom[23850]='h00000000;
    rd_cycle[23851] = 1'b1;  wr_cycle[23851] = 1'b0;  addr_rom[23851]='h000034ac;  wr_data_rom[23851]='h00000000;
    rd_cycle[23852] = 1'b1;  wr_cycle[23852] = 1'b0;  addr_rom[23852]='h000034b0;  wr_data_rom[23852]='h00000000;
    rd_cycle[23853] = 1'b1;  wr_cycle[23853] = 1'b0;  addr_rom[23853]='h000034b4;  wr_data_rom[23853]='h00000000;
    rd_cycle[23854] = 1'b1;  wr_cycle[23854] = 1'b0;  addr_rom[23854]='h000034b8;  wr_data_rom[23854]='h00000000;
    rd_cycle[23855] = 1'b1;  wr_cycle[23855] = 1'b0;  addr_rom[23855]='h000034bc;  wr_data_rom[23855]='h00000000;
    rd_cycle[23856] = 1'b1;  wr_cycle[23856] = 1'b0;  addr_rom[23856]='h000034c0;  wr_data_rom[23856]='h00000000;
    rd_cycle[23857] = 1'b1;  wr_cycle[23857] = 1'b0;  addr_rom[23857]='h000034c4;  wr_data_rom[23857]='h00000000;
    rd_cycle[23858] = 1'b1;  wr_cycle[23858] = 1'b0;  addr_rom[23858]='h000034c8;  wr_data_rom[23858]='h00000000;
    rd_cycle[23859] = 1'b1;  wr_cycle[23859] = 1'b0;  addr_rom[23859]='h000034cc;  wr_data_rom[23859]='h00000000;
    rd_cycle[23860] = 1'b1;  wr_cycle[23860] = 1'b0;  addr_rom[23860]='h000034d0;  wr_data_rom[23860]='h00000000;
    rd_cycle[23861] = 1'b1;  wr_cycle[23861] = 1'b0;  addr_rom[23861]='h000034d4;  wr_data_rom[23861]='h00000000;
    rd_cycle[23862] = 1'b1;  wr_cycle[23862] = 1'b0;  addr_rom[23862]='h000034d8;  wr_data_rom[23862]='h00000000;
    rd_cycle[23863] = 1'b1;  wr_cycle[23863] = 1'b0;  addr_rom[23863]='h000034dc;  wr_data_rom[23863]='h00000000;
    rd_cycle[23864] = 1'b1;  wr_cycle[23864] = 1'b0;  addr_rom[23864]='h000034e0;  wr_data_rom[23864]='h00000000;
    rd_cycle[23865] = 1'b1;  wr_cycle[23865] = 1'b0;  addr_rom[23865]='h000034e4;  wr_data_rom[23865]='h00000000;
    rd_cycle[23866] = 1'b1;  wr_cycle[23866] = 1'b0;  addr_rom[23866]='h000034e8;  wr_data_rom[23866]='h00000000;
    rd_cycle[23867] = 1'b1;  wr_cycle[23867] = 1'b0;  addr_rom[23867]='h000034ec;  wr_data_rom[23867]='h00000000;
    rd_cycle[23868] = 1'b1;  wr_cycle[23868] = 1'b0;  addr_rom[23868]='h000034f0;  wr_data_rom[23868]='h00000000;
    rd_cycle[23869] = 1'b1;  wr_cycle[23869] = 1'b0;  addr_rom[23869]='h000034f4;  wr_data_rom[23869]='h00000000;
    rd_cycle[23870] = 1'b1;  wr_cycle[23870] = 1'b0;  addr_rom[23870]='h000034f8;  wr_data_rom[23870]='h00000000;
    rd_cycle[23871] = 1'b1;  wr_cycle[23871] = 1'b0;  addr_rom[23871]='h000034fc;  wr_data_rom[23871]='h00000000;
    rd_cycle[23872] = 1'b1;  wr_cycle[23872] = 1'b0;  addr_rom[23872]='h00003500;  wr_data_rom[23872]='h00000000;
    rd_cycle[23873] = 1'b1;  wr_cycle[23873] = 1'b0;  addr_rom[23873]='h00003504;  wr_data_rom[23873]='h00000000;
    rd_cycle[23874] = 1'b1;  wr_cycle[23874] = 1'b0;  addr_rom[23874]='h00003508;  wr_data_rom[23874]='h00000000;
    rd_cycle[23875] = 1'b1;  wr_cycle[23875] = 1'b0;  addr_rom[23875]='h0000350c;  wr_data_rom[23875]='h00000000;
    rd_cycle[23876] = 1'b1;  wr_cycle[23876] = 1'b0;  addr_rom[23876]='h00003510;  wr_data_rom[23876]='h00000000;
    rd_cycle[23877] = 1'b1;  wr_cycle[23877] = 1'b0;  addr_rom[23877]='h00003514;  wr_data_rom[23877]='h00000000;
    rd_cycle[23878] = 1'b1;  wr_cycle[23878] = 1'b0;  addr_rom[23878]='h00003518;  wr_data_rom[23878]='h00000000;
    rd_cycle[23879] = 1'b1;  wr_cycle[23879] = 1'b0;  addr_rom[23879]='h0000351c;  wr_data_rom[23879]='h00000000;
    rd_cycle[23880] = 1'b1;  wr_cycle[23880] = 1'b0;  addr_rom[23880]='h00003520;  wr_data_rom[23880]='h00000000;
    rd_cycle[23881] = 1'b1;  wr_cycle[23881] = 1'b0;  addr_rom[23881]='h00003524;  wr_data_rom[23881]='h00000000;
    rd_cycle[23882] = 1'b1;  wr_cycle[23882] = 1'b0;  addr_rom[23882]='h00003528;  wr_data_rom[23882]='h00000000;
    rd_cycle[23883] = 1'b1;  wr_cycle[23883] = 1'b0;  addr_rom[23883]='h0000352c;  wr_data_rom[23883]='h00000000;
    rd_cycle[23884] = 1'b1;  wr_cycle[23884] = 1'b0;  addr_rom[23884]='h00003530;  wr_data_rom[23884]='h00000000;
    rd_cycle[23885] = 1'b1;  wr_cycle[23885] = 1'b0;  addr_rom[23885]='h00003534;  wr_data_rom[23885]='h00000000;
    rd_cycle[23886] = 1'b1;  wr_cycle[23886] = 1'b0;  addr_rom[23886]='h00003538;  wr_data_rom[23886]='h00000000;
    rd_cycle[23887] = 1'b1;  wr_cycle[23887] = 1'b0;  addr_rom[23887]='h0000353c;  wr_data_rom[23887]='h00000000;
    rd_cycle[23888] = 1'b1;  wr_cycle[23888] = 1'b0;  addr_rom[23888]='h00003540;  wr_data_rom[23888]='h00000000;
    rd_cycle[23889] = 1'b1;  wr_cycle[23889] = 1'b0;  addr_rom[23889]='h00003544;  wr_data_rom[23889]='h00000000;
    rd_cycle[23890] = 1'b1;  wr_cycle[23890] = 1'b0;  addr_rom[23890]='h00003548;  wr_data_rom[23890]='h00000000;
    rd_cycle[23891] = 1'b1;  wr_cycle[23891] = 1'b0;  addr_rom[23891]='h0000354c;  wr_data_rom[23891]='h00000000;
    rd_cycle[23892] = 1'b1;  wr_cycle[23892] = 1'b0;  addr_rom[23892]='h00003550;  wr_data_rom[23892]='h00000000;
    rd_cycle[23893] = 1'b1;  wr_cycle[23893] = 1'b0;  addr_rom[23893]='h00003554;  wr_data_rom[23893]='h00000000;
    rd_cycle[23894] = 1'b1;  wr_cycle[23894] = 1'b0;  addr_rom[23894]='h00003558;  wr_data_rom[23894]='h00000000;
    rd_cycle[23895] = 1'b1;  wr_cycle[23895] = 1'b0;  addr_rom[23895]='h0000355c;  wr_data_rom[23895]='h00000000;
    rd_cycle[23896] = 1'b1;  wr_cycle[23896] = 1'b0;  addr_rom[23896]='h00003560;  wr_data_rom[23896]='h00000000;
    rd_cycle[23897] = 1'b1;  wr_cycle[23897] = 1'b0;  addr_rom[23897]='h00003564;  wr_data_rom[23897]='h00000000;
    rd_cycle[23898] = 1'b1;  wr_cycle[23898] = 1'b0;  addr_rom[23898]='h00003568;  wr_data_rom[23898]='h00000000;
    rd_cycle[23899] = 1'b1;  wr_cycle[23899] = 1'b0;  addr_rom[23899]='h0000356c;  wr_data_rom[23899]='h00000000;
    rd_cycle[23900] = 1'b1;  wr_cycle[23900] = 1'b0;  addr_rom[23900]='h00003570;  wr_data_rom[23900]='h00000000;
    rd_cycle[23901] = 1'b1;  wr_cycle[23901] = 1'b0;  addr_rom[23901]='h00003574;  wr_data_rom[23901]='h00000000;
    rd_cycle[23902] = 1'b1;  wr_cycle[23902] = 1'b0;  addr_rom[23902]='h00003578;  wr_data_rom[23902]='h00000000;
    rd_cycle[23903] = 1'b1;  wr_cycle[23903] = 1'b0;  addr_rom[23903]='h0000357c;  wr_data_rom[23903]='h00000000;
    rd_cycle[23904] = 1'b1;  wr_cycle[23904] = 1'b0;  addr_rom[23904]='h00003580;  wr_data_rom[23904]='h00000000;
    rd_cycle[23905] = 1'b1;  wr_cycle[23905] = 1'b0;  addr_rom[23905]='h00003584;  wr_data_rom[23905]='h00000000;
    rd_cycle[23906] = 1'b1;  wr_cycle[23906] = 1'b0;  addr_rom[23906]='h00003588;  wr_data_rom[23906]='h00000000;
    rd_cycle[23907] = 1'b1;  wr_cycle[23907] = 1'b0;  addr_rom[23907]='h0000358c;  wr_data_rom[23907]='h00000000;
    rd_cycle[23908] = 1'b1;  wr_cycle[23908] = 1'b0;  addr_rom[23908]='h00003590;  wr_data_rom[23908]='h00000000;
    rd_cycle[23909] = 1'b1;  wr_cycle[23909] = 1'b0;  addr_rom[23909]='h00003594;  wr_data_rom[23909]='h00000000;
    rd_cycle[23910] = 1'b1;  wr_cycle[23910] = 1'b0;  addr_rom[23910]='h00003598;  wr_data_rom[23910]='h00000000;
    rd_cycle[23911] = 1'b1;  wr_cycle[23911] = 1'b0;  addr_rom[23911]='h0000359c;  wr_data_rom[23911]='h00000000;
    rd_cycle[23912] = 1'b1;  wr_cycle[23912] = 1'b0;  addr_rom[23912]='h000035a0;  wr_data_rom[23912]='h00000000;
    rd_cycle[23913] = 1'b1;  wr_cycle[23913] = 1'b0;  addr_rom[23913]='h000035a4;  wr_data_rom[23913]='h00000000;
    rd_cycle[23914] = 1'b1;  wr_cycle[23914] = 1'b0;  addr_rom[23914]='h000035a8;  wr_data_rom[23914]='h00000000;
    rd_cycle[23915] = 1'b1;  wr_cycle[23915] = 1'b0;  addr_rom[23915]='h000035ac;  wr_data_rom[23915]='h00000000;
    rd_cycle[23916] = 1'b1;  wr_cycle[23916] = 1'b0;  addr_rom[23916]='h000035b0;  wr_data_rom[23916]='h00000000;
    rd_cycle[23917] = 1'b1;  wr_cycle[23917] = 1'b0;  addr_rom[23917]='h000035b4;  wr_data_rom[23917]='h00000000;
    rd_cycle[23918] = 1'b1;  wr_cycle[23918] = 1'b0;  addr_rom[23918]='h000035b8;  wr_data_rom[23918]='h00000000;
    rd_cycle[23919] = 1'b1;  wr_cycle[23919] = 1'b0;  addr_rom[23919]='h000035bc;  wr_data_rom[23919]='h00000000;
    rd_cycle[23920] = 1'b1;  wr_cycle[23920] = 1'b0;  addr_rom[23920]='h000035c0;  wr_data_rom[23920]='h00000000;
    rd_cycle[23921] = 1'b1;  wr_cycle[23921] = 1'b0;  addr_rom[23921]='h000035c4;  wr_data_rom[23921]='h00000000;
    rd_cycle[23922] = 1'b1;  wr_cycle[23922] = 1'b0;  addr_rom[23922]='h000035c8;  wr_data_rom[23922]='h00000000;
    rd_cycle[23923] = 1'b1;  wr_cycle[23923] = 1'b0;  addr_rom[23923]='h000035cc;  wr_data_rom[23923]='h00000000;
    rd_cycle[23924] = 1'b1;  wr_cycle[23924] = 1'b0;  addr_rom[23924]='h000035d0;  wr_data_rom[23924]='h00000000;
    rd_cycle[23925] = 1'b1;  wr_cycle[23925] = 1'b0;  addr_rom[23925]='h000035d4;  wr_data_rom[23925]='h00000000;
    rd_cycle[23926] = 1'b1;  wr_cycle[23926] = 1'b0;  addr_rom[23926]='h000035d8;  wr_data_rom[23926]='h00000000;
    rd_cycle[23927] = 1'b1;  wr_cycle[23927] = 1'b0;  addr_rom[23927]='h000035dc;  wr_data_rom[23927]='h00000000;
    rd_cycle[23928] = 1'b1;  wr_cycle[23928] = 1'b0;  addr_rom[23928]='h000035e0;  wr_data_rom[23928]='h00000000;
    rd_cycle[23929] = 1'b1;  wr_cycle[23929] = 1'b0;  addr_rom[23929]='h000035e4;  wr_data_rom[23929]='h00000000;
    rd_cycle[23930] = 1'b1;  wr_cycle[23930] = 1'b0;  addr_rom[23930]='h000035e8;  wr_data_rom[23930]='h00000000;
    rd_cycle[23931] = 1'b1;  wr_cycle[23931] = 1'b0;  addr_rom[23931]='h000035ec;  wr_data_rom[23931]='h00000000;
    rd_cycle[23932] = 1'b1;  wr_cycle[23932] = 1'b0;  addr_rom[23932]='h000035f0;  wr_data_rom[23932]='h00000000;
    rd_cycle[23933] = 1'b1;  wr_cycle[23933] = 1'b0;  addr_rom[23933]='h000035f4;  wr_data_rom[23933]='h00000000;
    rd_cycle[23934] = 1'b1;  wr_cycle[23934] = 1'b0;  addr_rom[23934]='h000035f8;  wr_data_rom[23934]='h00000000;
    rd_cycle[23935] = 1'b1;  wr_cycle[23935] = 1'b0;  addr_rom[23935]='h000035fc;  wr_data_rom[23935]='h00000000;
    rd_cycle[23936] = 1'b1;  wr_cycle[23936] = 1'b0;  addr_rom[23936]='h00003600;  wr_data_rom[23936]='h00000000;
    rd_cycle[23937] = 1'b1;  wr_cycle[23937] = 1'b0;  addr_rom[23937]='h00003604;  wr_data_rom[23937]='h00000000;
    rd_cycle[23938] = 1'b1;  wr_cycle[23938] = 1'b0;  addr_rom[23938]='h00003608;  wr_data_rom[23938]='h00000000;
    rd_cycle[23939] = 1'b1;  wr_cycle[23939] = 1'b0;  addr_rom[23939]='h0000360c;  wr_data_rom[23939]='h00000000;
    rd_cycle[23940] = 1'b1;  wr_cycle[23940] = 1'b0;  addr_rom[23940]='h00003610;  wr_data_rom[23940]='h00000000;
    rd_cycle[23941] = 1'b1;  wr_cycle[23941] = 1'b0;  addr_rom[23941]='h00003614;  wr_data_rom[23941]='h00000000;
    rd_cycle[23942] = 1'b1;  wr_cycle[23942] = 1'b0;  addr_rom[23942]='h00003618;  wr_data_rom[23942]='h00000000;
    rd_cycle[23943] = 1'b1;  wr_cycle[23943] = 1'b0;  addr_rom[23943]='h0000361c;  wr_data_rom[23943]='h00000000;
    rd_cycle[23944] = 1'b1;  wr_cycle[23944] = 1'b0;  addr_rom[23944]='h00003620;  wr_data_rom[23944]='h00000000;
    rd_cycle[23945] = 1'b1;  wr_cycle[23945] = 1'b0;  addr_rom[23945]='h00003624;  wr_data_rom[23945]='h00000000;
    rd_cycle[23946] = 1'b1;  wr_cycle[23946] = 1'b0;  addr_rom[23946]='h00003628;  wr_data_rom[23946]='h00000000;
    rd_cycle[23947] = 1'b1;  wr_cycle[23947] = 1'b0;  addr_rom[23947]='h0000362c;  wr_data_rom[23947]='h00000000;
    rd_cycle[23948] = 1'b1;  wr_cycle[23948] = 1'b0;  addr_rom[23948]='h00003630;  wr_data_rom[23948]='h00000000;
    rd_cycle[23949] = 1'b1;  wr_cycle[23949] = 1'b0;  addr_rom[23949]='h00003634;  wr_data_rom[23949]='h00000000;
    rd_cycle[23950] = 1'b1;  wr_cycle[23950] = 1'b0;  addr_rom[23950]='h00003638;  wr_data_rom[23950]='h00000000;
    rd_cycle[23951] = 1'b1;  wr_cycle[23951] = 1'b0;  addr_rom[23951]='h0000363c;  wr_data_rom[23951]='h00000000;
    rd_cycle[23952] = 1'b1;  wr_cycle[23952] = 1'b0;  addr_rom[23952]='h00003640;  wr_data_rom[23952]='h00000000;
    rd_cycle[23953] = 1'b1;  wr_cycle[23953] = 1'b0;  addr_rom[23953]='h00003644;  wr_data_rom[23953]='h00000000;
    rd_cycle[23954] = 1'b1;  wr_cycle[23954] = 1'b0;  addr_rom[23954]='h00003648;  wr_data_rom[23954]='h00000000;
    rd_cycle[23955] = 1'b1;  wr_cycle[23955] = 1'b0;  addr_rom[23955]='h0000364c;  wr_data_rom[23955]='h00000000;
    rd_cycle[23956] = 1'b1;  wr_cycle[23956] = 1'b0;  addr_rom[23956]='h00003650;  wr_data_rom[23956]='h00000000;
    rd_cycle[23957] = 1'b1;  wr_cycle[23957] = 1'b0;  addr_rom[23957]='h00003654;  wr_data_rom[23957]='h00000000;
    rd_cycle[23958] = 1'b1;  wr_cycle[23958] = 1'b0;  addr_rom[23958]='h00003658;  wr_data_rom[23958]='h00000000;
    rd_cycle[23959] = 1'b1;  wr_cycle[23959] = 1'b0;  addr_rom[23959]='h0000365c;  wr_data_rom[23959]='h00000000;
    rd_cycle[23960] = 1'b1;  wr_cycle[23960] = 1'b0;  addr_rom[23960]='h00003660;  wr_data_rom[23960]='h00000000;
    rd_cycle[23961] = 1'b1;  wr_cycle[23961] = 1'b0;  addr_rom[23961]='h00003664;  wr_data_rom[23961]='h00000000;
    rd_cycle[23962] = 1'b1;  wr_cycle[23962] = 1'b0;  addr_rom[23962]='h00003668;  wr_data_rom[23962]='h00000000;
    rd_cycle[23963] = 1'b1;  wr_cycle[23963] = 1'b0;  addr_rom[23963]='h0000366c;  wr_data_rom[23963]='h00000000;
    rd_cycle[23964] = 1'b1;  wr_cycle[23964] = 1'b0;  addr_rom[23964]='h00003670;  wr_data_rom[23964]='h00000000;
    rd_cycle[23965] = 1'b1;  wr_cycle[23965] = 1'b0;  addr_rom[23965]='h00003674;  wr_data_rom[23965]='h00000000;
    rd_cycle[23966] = 1'b1;  wr_cycle[23966] = 1'b0;  addr_rom[23966]='h00003678;  wr_data_rom[23966]='h00000000;
    rd_cycle[23967] = 1'b1;  wr_cycle[23967] = 1'b0;  addr_rom[23967]='h0000367c;  wr_data_rom[23967]='h00000000;
    rd_cycle[23968] = 1'b1;  wr_cycle[23968] = 1'b0;  addr_rom[23968]='h00003680;  wr_data_rom[23968]='h00000000;
    rd_cycle[23969] = 1'b1;  wr_cycle[23969] = 1'b0;  addr_rom[23969]='h00003684;  wr_data_rom[23969]='h00000000;
    rd_cycle[23970] = 1'b1;  wr_cycle[23970] = 1'b0;  addr_rom[23970]='h00003688;  wr_data_rom[23970]='h00000000;
    rd_cycle[23971] = 1'b1;  wr_cycle[23971] = 1'b0;  addr_rom[23971]='h0000368c;  wr_data_rom[23971]='h00000000;
    rd_cycle[23972] = 1'b1;  wr_cycle[23972] = 1'b0;  addr_rom[23972]='h00003690;  wr_data_rom[23972]='h00000000;
    rd_cycle[23973] = 1'b1;  wr_cycle[23973] = 1'b0;  addr_rom[23973]='h00003694;  wr_data_rom[23973]='h00000000;
    rd_cycle[23974] = 1'b1;  wr_cycle[23974] = 1'b0;  addr_rom[23974]='h00003698;  wr_data_rom[23974]='h00000000;
    rd_cycle[23975] = 1'b1;  wr_cycle[23975] = 1'b0;  addr_rom[23975]='h0000369c;  wr_data_rom[23975]='h00000000;
    rd_cycle[23976] = 1'b1;  wr_cycle[23976] = 1'b0;  addr_rom[23976]='h000036a0;  wr_data_rom[23976]='h00000000;
    rd_cycle[23977] = 1'b1;  wr_cycle[23977] = 1'b0;  addr_rom[23977]='h000036a4;  wr_data_rom[23977]='h00000000;
    rd_cycle[23978] = 1'b1;  wr_cycle[23978] = 1'b0;  addr_rom[23978]='h000036a8;  wr_data_rom[23978]='h00000000;
    rd_cycle[23979] = 1'b1;  wr_cycle[23979] = 1'b0;  addr_rom[23979]='h000036ac;  wr_data_rom[23979]='h00000000;
    rd_cycle[23980] = 1'b1;  wr_cycle[23980] = 1'b0;  addr_rom[23980]='h000036b0;  wr_data_rom[23980]='h00000000;
    rd_cycle[23981] = 1'b1;  wr_cycle[23981] = 1'b0;  addr_rom[23981]='h000036b4;  wr_data_rom[23981]='h00000000;
    rd_cycle[23982] = 1'b1;  wr_cycle[23982] = 1'b0;  addr_rom[23982]='h000036b8;  wr_data_rom[23982]='h00000000;
    rd_cycle[23983] = 1'b1;  wr_cycle[23983] = 1'b0;  addr_rom[23983]='h000036bc;  wr_data_rom[23983]='h00000000;
    rd_cycle[23984] = 1'b1;  wr_cycle[23984] = 1'b0;  addr_rom[23984]='h000036c0;  wr_data_rom[23984]='h00000000;
    rd_cycle[23985] = 1'b1;  wr_cycle[23985] = 1'b0;  addr_rom[23985]='h000036c4;  wr_data_rom[23985]='h00000000;
    rd_cycle[23986] = 1'b1;  wr_cycle[23986] = 1'b0;  addr_rom[23986]='h000036c8;  wr_data_rom[23986]='h00000000;
    rd_cycle[23987] = 1'b1;  wr_cycle[23987] = 1'b0;  addr_rom[23987]='h000036cc;  wr_data_rom[23987]='h00000000;
    rd_cycle[23988] = 1'b1;  wr_cycle[23988] = 1'b0;  addr_rom[23988]='h000036d0;  wr_data_rom[23988]='h00000000;
    rd_cycle[23989] = 1'b1;  wr_cycle[23989] = 1'b0;  addr_rom[23989]='h000036d4;  wr_data_rom[23989]='h00000000;
    rd_cycle[23990] = 1'b1;  wr_cycle[23990] = 1'b0;  addr_rom[23990]='h000036d8;  wr_data_rom[23990]='h00000000;
    rd_cycle[23991] = 1'b1;  wr_cycle[23991] = 1'b0;  addr_rom[23991]='h000036dc;  wr_data_rom[23991]='h00000000;
    rd_cycle[23992] = 1'b1;  wr_cycle[23992] = 1'b0;  addr_rom[23992]='h000036e0;  wr_data_rom[23992]='h00000000;
    rd_cycle[23993] = 1'b1;  wr_cycle[23993] = 1'b0;  addr_rom[23993]='h000036e4;  wr_data_rom[23993]='h00000000;
    rd_cycle[23994] = 1'b1;  wr_cycle[23994] = 1'b0;  addr_rom[23994]='h000036e8;  wr_data_rom[23994]='h00000000;
    rd_cycle[23995] = 1'b1;  wr_cycle[23995] = 1'b0;  addr_rom[23995]='h000036ec;  wr_data_rom[23995]='h00000000;
    rd_cycle[23996] = 1'b1;  wr_cycle[23996] = 1'b0;  addr_rom[23996]='h000036f0;  wr_data_rom[23996]='h00000000;
    rd_cycle[23997] = 1'b1;  wr_cycle[23997] = 1'b0;  addr_rom[23997]='h000036f4;  wr_data_rom[23997]='h00000000;
    rd_cycle[23998] = 1'b1;  wr_cycle[23998] = 1'b0;  addr_rom[23998]='h000036f8;  wr_data_rom[23998]='h00000000;
    rd_cycle[23999] = 1'b1;  wr_cycle[23999] = 1'b0;  addr_rom[23999]='h000036fc;  wr_data_rom[23999]='h00000000;
    rd_cycle[24000] = 1'b1;  wr_cycle[24000] = 1'b0;  addr_rom[24000]='h00003700;  wr_data_rom[24000]='h00000000;
    rd_cycle[24001] = 1'b1;  wr_cycle[24001] = 1'b0;  addr_rom[24001]='h00003704;  wr_data_rom[24001]='h00000000;
    rd_cycle[24002] = 1'b1;  wr_cycle[24002] = 1'b0;  addr_rom[24002]='h00003708;  wr_data_rom[24002]='h00000000;
    rd_cycle[24003] = 1'b1;  wr_cycle[24003] = 1'b0;  addr_rom[24003]='h0000370c;  wr_data_rom[24003]='h00000000;
    rd_cycle[24004] = 1'b1;  wr_cycle[24004] = 1'b0;  addr_rom[24004]='h00003710;  wr_data_rom[24004]='h00000000;
    rd_cycle[24005] = 1'b1;  wr_cycle[24005] = 1'b0;  addr_rom[24005]='h00003714;  wr_data_rom[24005]='h00000000;
    rd_cycle[24006] = 1'b1;  wr_cycle[24006] = 1'b0;  addr_rom[24006]='h00003718;  wr_data_rom[24006]='h00000000;
    rd_cycle[24007] = 1'b1;  wr_cycle[24007] = 1'b0;  addr_rom[24007]='h0000371c;  wr_data_rom[24007]='h00000000;
    rd_cycle[24008] = 1'b1;  wr_cycle[24008] = 1'b0;  addr_rom[24008]='h00003720;  wr_data_rom[24008]='h00000000;
    rd_cycle[24009] = 1'b1;  wr_cycle[24009] = 1'b0;  addr_rom[24009]='h00003724;  wr_data_rom[24009]='h00000000;
    rd_cycle[24010] = 1'b1;  wr_cycle[24010] = 1'b0;  addr_rom[24010]='h00003728;  wr_data_rom[24010]='h00000000;
    rd_cycle[24011] = 1'b1;  wr_cycle[24011] = 1'b0;  addr_rom[24011]='h0000372c;  wr_data_rom[24011]='h00000000;
    rd_cycle[24012] = 1'b1;  wr_cycle[24012] = 1'b0;  addr_rom[24012]='h00003730;  wr_data_rom[24012]='h00000000;
    rd_cycle[24013] = 1'b1;  wr_cycle[24013] = 1'b0;  addr_rom[24013]='h00003734;  wr_data_rom[24013]='h00000000;
    rd_cycle[24014] = 1'b1;  wr_cycle[24014] = 1'b0;  addr_rom[24014]='h00003738;  wr_data_rom[24014]='h00000000;
    rd_cycle[24015] = 1'b1;  wr_cycle[24015] = 1'b0;  addr_rom[24015]='h0000373c;  wr_data_rom[24015]='h00000000;
    rd_cycle[24016] = 1'b1;  wr_cycle[24016] = 1'b0;  addr_rom[24016]='h00003740;  wr_data_rom[24016]='h00000000;
    rd_cycle[24017] = 1'b1;  wr_cycle[24017] = 1'b0;  addr_rom[24017]='h00003744;  wr_data_rom[24017]='h00000000;
    rd_cycle[24018] = 1'b1;  wr_cycle[24018] = 1'b0;  addr_rom[24018]='h00003748;  wr_data_rom[24018]='h00000000;
    rd_cycle[24019] = 1'b1;  wr_cycle[24019] = 1'b0;  addr_rom[24019]='h0000374c;  wr_data_rom[24019]='h00000000;
    rd_cycle[24020] = 1'b1;  wr_cycle[24020] = 1'b0;  addr_rom[24020]='h00003750;  wr_data_rom[24020]='h00000000;
    rd_cycle[24021] = 1'b1;  wr_cycle[24021] = 1'b0;  addr_rom[24021]='h00003754;  wr_data_rom[24021]='h00000000;
    rd_cycle[24022] = 1'b1;  wr_cycle[24022] = 1'b0;  addr_rom[24022]='h00003758;  wr_data_rom[24022]='h00000000;
    rd_cycle[24023] = 1'b1;  wr_cycle[24023] = 1'b0;  addr_rom[24023]='h0000375c;  wr_data_rom[24023]='h00000000;
    rd_cycle[24024] = 1'b1;  wr_cycle[24024] = 1'b0;  addr_rom[24024]='h00003760;  wr_data_rom[24024]='h00000000;
    rd_cycle[24025] = 1'b1;  wr_cycle[24025] = 1'b0;  addr_rom[24025]='h00003764;  wr_data_rom[24025]='h00000000;
    rd_cycle[24026] = 1'b1;  wr_cycle[24026] = 1'b0;  addr_rom[24026]='h00003768;  wr_data_rom[24026]='h00000000;
    rd_cycle[24027] = 1'b1;  wr_cycle[24027] = 1'b0;  addr_rom[24027]='h0000376c;  wr_data_rom[24027]='h00000000;
    rd_cycle[24028] = 1'b1;  wr_cycle[24028] = 1'b0;  addr_rom[24028]='h00003770;  wr_data_rom[24028]='h00000000;
    rd_cycle[24029] = 1'b1;  wr_cycle[24029] = 1'b0;  addr_rom[24029]='h00003774;  wr_data_rom[24029]='h00000000;
    rd_cycle[24030] = 1'b1;  wr_cycle[24030] = 1'b0;  addr_rom[24030]='h00003778;  wr_data_rom[24030]='h00000000;
    rd_cycle[24031] = 1'b1;  wr_cycle[24031] = 1'b0;  addr_rom[24031]='h0000377c;  wr_data_rom[24031]='h00000000;
    rd_cycle[24032] = 1'b1;  wr_cycle[24032] = 1'b0;  addr_rom[24032]='h00003780;  wr_data_rom[24032]='h00000000;
    rd_cycle[24033] = 1'b1;  wr_cycle[24033] = 1'b0;  addr_rom[24033]='h00003784;  wr_data_rom[24033]='h00000000;
    rd_cycle[24034] = 1'b1;  wr_cycle[24034] = 1'b0;  addr_rom[24034]='h00003788;  wr_data_rom[24034]='h00000000;
    rd_cycle[24035] = 1'b1;  wr_cycle[24035] = 1'b0;  addr_rom[24035]='h0000378c;  wr_data_rom[24035]='h00000000;
    rd_cycle[24036] = 1'b1;  wr_cycle[24036] = 1'b0;  addr_rom[24036]='h00003790;  wr_data_rom[24036]='h00000000;
    rd_cycle[24037] = 1'b1;  wr_cycle[24037] = 1'b0;  addr_rom[24037]='h00003794;  wr_data_rom[24037]='h00000000;
    rd_cycle[24038] = 1'b1;  wr_cycle[24038] = 1'b0;  addr_rom[24038]='h00003798;  wr_data_rom[24038]='h00000000;
    rd_cycle[24039] = 1'b1;  wr_cycle[24039] = 1'b0;  addr_rom[24039]='h0000379c;  wr_data_rom[24039]='h00000000;
    rd_cycle[24040] = 1'b1;  wr_cycle[24040] = 1'b0;  addr_rom[24040]='h000037a0;  wr_data_rom[24040]='h00000000;
    rd_cycle[24041] = 1'b1;  wr_cycle[24041] = 1'b0;  addr_rom[24041]='h000037a4;  wr_data_rom[24041]='h00000000;
    rd_cycle[24042] = 1'b1;  wr_cycle[24042] = 1'b0;  addr_rom[24042]='h000037a8;  wr_data_rom[24042]='h00000000;
    rd_cycle[24043] = 1'b1;  wr_cycle[24043] = 1'b0;  addr_rom[24043]='h000037ac;  wr_data_rom[24043]='h00000000;
    rd_cycle[24044] = 1'b1;  wr_cycle[24044] = 1'b0;  addr_rom[24044]='h000037b0;  wr_data_rom[24044]='h00000000;
    rd_cycle[24045] = 1'b1;  wr_cycle[24045] = 1'b0;  addr_rom[24045]='h000037b4;  wr_data_rom[24045]='h00000000;
    rd_cycle[24046] = 1'b1;  wr_cycle[24046] = 1'b0;  addr_rom[24046]='h000037b8;  wr_data_rom[24046]='h00000000;
    rd_cycle[24047] = 1'b1;  wr_cycle[24047] = 1'b0;  addr_rom[24047]='h000037bc;  wr_data_rom[24047]='h00000000;
    rd_cycle[24048] = 1'b1;  wr_cycle[24048] = 1'b0;  addr_rom[24048]='h000037c0;  wr_data_rom[24048]='h00000000;
    rd_cycle[24049] = 1'b1;  wr_cycle[24049] = 1'b0;  addr_rom[24049]='h000037c4;  wr_data_rom[24049]='h00000000;
    rd_cycle[24050] = 1'b1;  wr_cycle[24050] = 1'b0;  addr_rom[24050]='h000037c8;  wr_data_rom[24050]='h00000000;
    rd_cycle[24051] = 1'b1;  wr_cycle[24051] = 1'b0;  addr_rom[24051]='h000037cc;  wr_data_rom[24051]='h00000000;
    rd_cycle[24052] = 1'b1;  wr_cycle[24052] = 1'b0;  addr_rom[24052]='h000037d0;  wr_data_rom[24052]='h00000000;
    rd_cycle[24053] = 1'b1;  wr_cycle[24053] = 1'b0;  addr_rom[24053]='h000037d4;  wr_data_rom[24053]='h00000000;
    rd_cycle[24054] = 1'b1;  wr_cycle[24054] = 1'b0;  addr_rom[24054]='h000037d8;  wr_data_rom[24054]='h00000000;
    rd_cycle[24055] = 1'b1;  wr_cycle[24055] = 1'b0;  addr_rom[24055]='h000037dc;  wr_data_rom[24055]='h00000000;
    rd_cycle[24056] = 1'b1;  wr_cycle[24056] = 1'b0;  addr_rom[24056]='h000037e0;  wr_data_rom[24056]='h00000000;
    rd_cycle[24057] = 1'b1;  wr_cycle[24057] = 1'b0;  addr_rom[24057]='h000037e4;  wr_data_rom[24057]='h00000000;
    rd_cycle[24058] = 1'b1;  wr_cycle[24058] = 1'b0;  addr_rom[24058]='h000037e8;  wr_data_rom[24058]='h00000000;
    rd_cycle[24059] = 1'b1;  wr_cycle[24059] = 1'b0;  addr_rom[24059]='h000037ec;  wr_data_rom[24059]='h00000000;
    rd_cycle[24060] = 1'b1;  wr_cycle[24060] = 1'b0;  addr_rom[24060]='h000037f0;  wr_data_rom[24060]='h00000000;
    rd_cycle[24061] = 1'b1;  wr_cycle[24061] = 1'b0;  addr_rom[24061]='h000037f4;  wr_data_rom[24061]='h00000000;
    rd_cycle[24062] = 1'b1;  wr_cycle[24062] = 1'b0;  addr_rom[24062]='h000037f8;  wr_data_rom[24062]='h00000000;
    rd_cycle[24063] = 1'b1;  wr_cycle[24063] = 1'b0;  addr_rom[24063]='h000037fc;  wr_data_rom[24063]='h00000000;
    rd_cycle[24064] = 1'b1;  wr_cycle[24064] = 1'b0;  addr_rom[24064]='h00003800;  wr_data_rom[24064]='h00000000;
    rd_cycle[24065] = 1'b1;  wr_cycle[24065] = 1'b0;  addr_rom[24065]='h00003804;  wr_data_rom[24065]='h00000000;
    rd_cycle[24066] = 1'b1;  wr_cycle[24066] = 1'b0;  addr_rom[24066]='h00003808;  wr_data_rom[24066]='h00000000;
    rd_cycle[24067] = 1'b1;  wr_cycle[24067] = 1'b0;  addr_rom[24067]='h0000380c;  wr_data_rom[24067]='h00000000;
    rd_cycle[24068] = 1'b1;  wr_cycle[24068] = 1'b0;  addr_rom[24068]='h00003810;  wr_data_rom[24068]='h00000000;
    rd_cycle[24069] = 1'b1;  wr_cycle[24069] = 1'b0;  addr_rom[24069]='h00003814;  wr_data_rom[24069]='h00000000;
    rd_cycle[24070] = 1'b1;  wr_cycle[24070] = 1'b0;  addr_rom[24070]='h00003818;  wr_data_rom[24070]='h00000000;
    rd_cycle[24071] = 1'b1;  wr_cycle[24071] = 1'b0;  addr_rom[24071]='h0000381c;  wr_data_rom[24071]='h00000000;
    rd_cycle[24072] = 1'b1;  wr_cycle[24072] = 1'b0;  addr_rom[24072]='h00003820;  wr_data_rom[24072]='h00000000;
    rd_cycle[24073] = 1'b1;  wr_cycle[24073] = 1'b0;  addr_rom[24073]='h00003824;  wr_data_rom[24073]='h00000000;
    rd_cycle[24074] = 1'b1;  wr_cycle[24074] = 1'b0;  addr_rom[24074]='h00003828;  wr_data_rom[24074]='h00000000;
    rd_cycle[24075] = 1'b1;  wr_cycle[24075] = 1'b0;  addr_rom[24075]='h0000382c;  wr_data_rom[24075]='h00000000;
    rd_cycle[24076] = 1'b1;  wr_cycle[24076] = 1'b0;  addr_rom[24076]='h00003830;  wr_data_rom[24076]='h00000000;
    rd_cycle[24077] = 1'b1;  wr_cycle[24077] = 1'b0;  addr_rom[24077]='h00003834;  wr_data_rom[24077]='h00000000;
    rd_cycle[24078] = 1'b1;  wr_cycle[24078] = 1'b0;  addr_rom[24078]='h00003838;  wr_data_rom[24078]='h00000000;
    rd_cycle[24079] = 1'b1;  wr_cycle[24079] = 1'b0;  addr_rom[24079]='h0000383c;  wr_data_rom[24079]='h00000000;
    rd_cycle[24080] = 1'b1;  wr_cycle[24080] = 1'b0;  addr_rom[24080]='h00003840;  wr_data_rom[24080]='h00000000;
    rd_cycle[24081] = 1'b1;  wr_cycle[24081] = 1'b0;  addr_rom[24081]='h00003844;  wr_data_rom[24081]='h00000000;
    rd_cycle[24082] = 1'b1;  wr_cycle[24082] = 1'b0;  addr_rom[24082]='h00003848;  wr_data_rom[24082]='h00000000;
    rd_cycle[24083] = 1'b1;  wr_cycle[24083] = 1'b0;  addr_rom[24083]='h0000384c;  wr_data_rom[24083]='h00000000;
    rd_cycle[24084] = 1'b1;  wr_cycle[24084] = 1'b0;  addr_rom[24084]='h00003850;  wr_data_rom[24084]='h00000000;
    rd_cycle[24085] = 1'b1;  wr_cycle[24085] = 1'b0;  addr_rom[24085]='h00003854;  wr_data_rom[24085]='h00000000;
    rd_cycle[24086] = 1'b1;  wr_cycle[24086] = 1'b0;  addr_rom[24086]='h00003858;  wr_data_rom[24086]='h00000000;
    rd_cycle[24087] = 1'b1;  wr_cycle[24087] = 1'b0;  addr_rom[24087]='h0000385c;  wr_data_rom[24087]='h00000000;
    rd_cycle[24088] = 1'b1;  wr_cycle[24088] = 1'b0;  addr_rom[24088]='h00003860;  wr_data_rom[24088]='h00000000;
    rd_cycle[24089] = 1'b1;  wr_cycle[24089] = 1'b0;  addr_rom[24089]='h00003864;  wr_data_rom[24089]='h00000000;
    rd_cycle[24090] = 1'b1;  wr_cycle[24090] = 1'b0;  addr_rom[24090]='h00003868;  wr_data_rom[24090]='h00000000;
    rd_cycle[24091] = 1'b1;  wr_cycle[24091] = 1'b0;  addr_rom[24091]='h0000386c;  wr_data_rom[24091]='h00000000;
    rd_cycle[24092] = 1'b1;  wr_cycle[24092] = 1'b0;  addr_rom[24092]='h00003870;  wr_data_rom[24092]='h00000000;
    rd_cycle[24093] = 1'b1;  wr_cycle[24093] = 1'b0;  addr_rom[24093]='h00003874;  wr_data_rom[24093]='h00000000;
    rd_cycle[24094] = 1'b1;  wr_cycle[24094] = 1'b0;  addr_rom[24094]='h00003878;  wr_data_rom[24094]='h00000000;
    rd_cycle[24095] = 1'b1;  wr_cycle[24095] = 1'b0;  addr_rom[24095]='h0000387c;  wr_data_rom[24095]='h00000000;
    rd_cycle[24096] = 1'b1;  wr_cycle[24096] = 1'b0;  addr_rom[24096]='h00003880;  wr_data_rom[24096]='h00000000;
    rd_cycle[24097] = 1'b1;  wr_cycle[24097] = 1'b0;  addr_rom[24097]='h00003884;  wr_data_rom[24097]='h00000000;
    rd_cycle[24098] = 1'b1;  wr_cycle[24098] = 1'b0;  addr_rom[24098]='h00003888;  wr_data_rom[24098]='h00000000;
    rd_cycle[24099] = 1'b1;  wr_cycle[24099] = 1'b0;  addr_rom[24099]='h0000388c;  wr_data_rom[24099]='h00000000;
    rd_cycle[24100] = 1'b1;  wr_cycle[24100] = 1'b0;  addr_rom[24100]='h00003890;  wr_data_rom[24100]='h00000000;
    rd_cycle[24101] = 1'b1;  wr_cycle[24101] = 1'b0;  addr_rom[24101]='h00003894;  wr_data_rom[24101]='h00000000;
    rd_cycle[24102] = 1'b1;  wr_cycle[24102] = 1'b0;  addr_rom[24102]='h00003898;  wr_data_rom[24102]='h00000000;
    rd_cycle[24103] = 1'b1;  wr_cycle[24103] = 1'b0;  addr_rom[24103]='h0000389c;  wr_data_rom[24103]='h00000000;
    rd_cycle[24104] = 1'b1;  wr_cycle[24104] = 1'b0;  addr_rom[24104]='h000038a0;  wr_data_rom[24104]='h00000000;
    rd_cycle[24105] = 1'b1;  wr_cycle[24105] = 1'b0;  addr_rom[24105]='h000038a4;  wr_data_rom[24105]='h00000000;
    rd_cycle[24106] = 1'b1;  wr_cycle[24106] = 1'b0;  addr_rom[24106]='h000038a8;  wr_data_rom[24106]='h00000000;
    rd_cycle[24107] = 1'b1;  wr_cycle[24107] = 1'b0;  addr_rom[24107]='h000038ac;  wr_data_rom[24107]='h00000000;
    rd_cycle[24108] = 1'b1;  wr_cycle[24108] = 1'b0;  addr_rom[24108]='h000038b0;  wr_data_rom[24108]='h00000000;
    rd_cycle[24109] = 1'b1;  wr_cycle[24109] = 1'b0;  addr_rom[24109]='h000038b4;  wr_data_rom[24109]='h00000000;
    rd_cycle[24110] = 1'b1;  wr_cycle[24110] = 1'b0;  addr_rom[24110]='h000038b8;  wr_data_rom[24110]='h00000000;
    rd_cycle[24111] = 1'b1;  wr_cycle[24111] = 1'b0;  addr_rom[24111]='h000038bc;  wr_data_rom[24111]='h00000000;
    rd_cycle[24112] = 1'b1;  wr_cycle[24112] = 1'b0;  addr_rom[24112]='h000038c0;  wr_data_rom[24112]='h00000000;
    rd_cycle[24113] = 1'b1;  wr_cycle[24113] = 1'b0;  addr_rom[24113]='h000038c4;  wr_data_rom[24113]='h00000000;
    rd_cycle[24114] = 1'b1;  wr_cycle[24114] = 1'b0;  addr_rom[24114]='h000038c8;  wr_data_rom[24114]='h00000000;
    rd_cycle[24115] = 1'b1;  wr_cycle[24115] = 1'b0;  addr_rom[24115]='h000038cc;  wr_data_rom[24115]='h00000000;
    rd_cycle[24116] = 1'b1;  wr_cycle[24116] = 1'b0;  addr_rom[24116]='h000038d0;  wr_data_rom[24116]='h00000000;
    rd_cycle[24117] = 1'b1;  wr_cycle[24117] = 1'b0;  addr_rom[24117]='h000038d4;  wr_data_rom[24117]='h00000000;
    rd_cycle[24118] = 1'b1;  wr_cycle[24118] = 1'b0;  addr_rom[24118]='h000038d8;  wr_data_rom[24118]='h00000000;
    rd_cycle[24119] = 1'b1;  wr_cycle[24119] = 1'b0;  addr_rom[24119]='h000038dc;  wr_data_rom[24119]='h00000000;
    rd_cycle[24120] = 1'b1;  wr_cycle[24120] = 1'b0;  addr_rom[24120]='h000038e0;  wr_data_rom[24120]='h00000000;
    rd_cycle[24121] = 1'b1;  wr_cycle[24121] = 1'b0;  addr_rom[24121]='h000038e4;  wr_data_rom[24121]='h00000000;
    rd_cycle[24122] = 1'b1;  wr_cycle[24122] = 1'b0;  addr_rom[24122]='h000038e8;  wr_data_rom[24122]='h00000000;
    rd_cycle[24123] = 1'b1;  wr_cycle[24123] = 1'b0;  addr_rom[24123]='h000038ec;  wr_data_rom[24123]='h00000000;
    rd_cycle[24124] = 1'b1;  wr_cycle[24124] = 1'b0;  addr_rom[24124]='h000038f0;  wr_data_rom[24124]='h00000000;
    rd_cycle[24125] = 1'b1;  wr_cycle[24125] = 1'b0;  addr_rom[24125]='h000038f4;  wr_data_rom[24125]='h00000000;
    rd_cycle[24126] = 1'b1;  wr_cycle[24126] = 1'b0;  addr_rom[24126]='h000038f8;  wr_data_rom[24126]='h00000000;
    rd_cycle[24127] = 1'b1;  wr_cycle[24127] = 1'b0;  addr_rom[24127]='h000038fc;  wr_data_rom[24127]='h00000000;
    rd_cycle[24128] = 1'b1;  wr_cycle[24128] = 1'b0;  addr_rom[24128]='h00003900;  wr_data_rom[24128]='h00000000;
    rd_cycle[24129] = 1'b1;  wr_cycle[24129] = 1'b0;  addr_rom[24129]='h00003904;  wr_data_rom[24129]='h00000000;
    rd_cycle[24130] = 1'b1;  wr_cycle[24130] = 1'b0;  addr_rom[24130]='h00003908;  wr_data_rom[24130]='h00000000;
    rd_cycle[24131] = 1'b1;  wr_cycle[24131] = 1'b0;  addr_rom[24131]='h0000390c;  wr_data_rom[24131]='h00000000;
    rd_cycle[24132] = 1'b1;  wr_cycle[24132] = 1'b0;  addr_rom[24132]='h00003910;  wr_data_rom[24132]='h00000000;
    rd_cycle[24133] = 1'b1;  wr_cycle[24133] = 1'b0;  addr_rom[24133]='h00003914;  wr_data_rom[24133]='h00000000;
    rd_cycle[24134] = 1'b1;  wr_cycle[24134] = 1'b0;  addr_rom[24134]='h00003918;  wr_data_rom[24134]='h00000000;
    rd_cycle[24135] = 1'b1;  wr_cycle[24135] = 1'b0;  addr_rom[24135]='h0000391c;  wr_data_rom[24135]='h00000000;
    rd_cycle[24136] = 1'b1;  wr_cycle[24136] = 1'b0;  addr_rom[24136]='h00003920;  wr_data_rom[24136]='h00000000;
    rd_cycle[24137] = 1'b1;  wr_cycle[24137] = 1'b0;  addr_rom[24137]='h00003924;  wr_data_rom[24137]='h00000000;
    rd_cycle[24138] = 1'b1;  wr_cycle[24138] = 1'b0;  addr_rom[24138]='h00003928;  wr_data_rom[24138]='h00000000;
    rd_cycle[24139] = 1'b1;  wr_cycle[24139] = 1'b0;  addr_rom[24139]='h0000392c;  wr_data_rom[24139]='h00000000;
    rd_cycle[24140] = 1'b1;  wr_cycle[24140] = 1'b0;  addr_rom[24140]='h00003930;  wr_data_rom[24140]='h00000000;
    rd_cycle[24141] = 1'b1;  wr_cycle[24141] = 1'b0;  addr_rom[24141]='h00003934;  wr_data_rom[24141]='h00000000;
    rd_cycle[24142] = 1'b1;  wr_cycle[24142] = 1'b0;  addr_rom[24142]='h00003938;  wr_data_rom[24142]='h00000000;
    rd_cycle[24143] = 1'b1;  wr_cycle[24143] = 1'b0;  addr_rom[24143]='h0000393c;  wr_data_rom[24143]='h00000000;
    rd_cycle[24144] = 1'b1;  wr_cycle[24144] = 1'b0;  addr_rom[24144]='h00003940;  wr_data_rom[24144]='h00000000;
    rd_cycle[24145] = 1'b1;  wr_cycle[24145] = 1'b0;  addr_rom[24145]='h00003944;  wr_data_rom[24145]='h00000000;
    rd_cycle[24146] = 1'b1;  wr_cycle[24146] = 1'b0;  addr_rom[24146]='h00003948;  wr_data_rom[24146]='h00000000;
    rd_cycle[24147] = 1'b1;  wr_cycle[24147] = 1'b0;  addr_rom[24147]='h0000394c;  wr_data_rom[24147]='h00000000;
    rd_cycle[24148] = 1'b1;  wr_cycle[24148] = 1'b0;  addr_rom[24148]='h00003950;  wr_data_rom[24148]='h00000000;
    rd_cycle[24149] = 1'b1;  wr_cycle[24149] = 1'b0;  addr_rom[24149]='h00003954;  wr_data_rom[24149]='h00000000;
    rd_cycle[24150] = 1'b1;  wr_cycle[24150] = 1'b0;  addr_rom[24150]='h00003958;  wr_data_rom[24150]='h00000000;
    rd_cycle[24151] = 1'b1;  wr_cycle[24151] = 1'b0;  addr_rom[24151]='h0000395c;  wr_data_rom[24151]='h00000000;
    rd_cycle[24152] = 1'b1;  wr_cycle[24152] = 1'b0;  addr_rom[24152]='h00003960;  wr_data_rom[24152]='h00000000;
    rd_cycle[24153] = 1'b1;  wr_cycle[24153] = 1'b0;  addr_rom[24153]='h00003964;  wr_data_rom[24153]='h00000000;
    rd_cycle[24154] = 1'b1;  wr_cycle[24154] = 1'b0;  addr_rom[24154]='h00003968;  wr_data_rom[24154]='h00000000;
    rd_cycle[24155] = 1'b1;  wr_cycle[24155] = 1'b0;  addr_rom[24155]='h0000396c;  wr_data_rom[24155]='h00000000;
    rd_cycle[24156] = 1'b1;  wr_cycle[24156] = 1'b0;  addr_rom[24156]='h00003970;  wr_data_rom[24156]='h00000000;
    rd_cycle[24157] = 1'b1;  wr_cycle[24157] = 1'b0;  addr_rom[24157]='h00003974;  wr_data_rom[24157]='h00000000;
    rd_cycle[24158] = 1'b1;  wr_cycle[24158] = 1'b0;  addr_rom[24158]='h00003978;  wr_data_rom[24158]='h00000000;
    rd_cycle[24159] = 1'b1;  wr_cycle[24159] = 1'b0;  addr_rom[24159]='h0000397c;  wr_data_rom[24159]='h00000000;
    rd_cycle[24160] = 1'b1;  wr_cycle[24160] = 1'b0;  addr_rom[24160]='h00003980;  wr_data_rom[24160]='h00000000;
    rd_cycle[24161] = 1'b1;  wr_cycle[24161] = 1'b0;  addr_rom[24161]='h00003984;  wr_data_rom[24161]='h00000000;
    rd_cycle[24162] = 1'b1;  wr_cycle[24162] = 1'b0;  addr_rom[24162]='h00003988;  wr_data_rom[24162]='h00000000;
    rd_cycle[24163] = 1'b1;  wr_cycle[24163] = 1'b0;  addr_rom[24163]='h0000398c;  wr_data_rom[24163]='h00000000;
    rd_cycle[24164] = 1'b1;  wr_cycle[24164] = 1'b0;  addr_rom[24164]='h00003990;  wr_data_rom[24164]='h00000000;
    rd_cycle[24165] = 1'b1;  wr_cycle[24165] = 1'b0;  addr_rom[24165]='h00003994;  wr_data_rom[24165]='h00000000;
    rd_cycle[24166] = 1'b1;  wr_cycle[24166] = 1'b0;  addr_rom[24166]='h00003998;  wr_data_rom[24166]='h00000000;
    rd_cycle[24167] = 1'b1;  wr_cycle[24167] = 1'b0;  addr_rom[24167]='h0000399c;  wr_data_rom[24167]='h00000000;
    rd_cycle[24168] = 1'b1;  wr_cycle[24168] = 1'b0;  addr_rom[24168]='h000039a0;  wr_data_rom[24168]='h00000000;
    rd_cycle[24169] = 1'b1;  wr_cycle[24169] = 1'b0;  addr_rom[24169]='h000039a4;  wr_data_rom[24169]='h00000000;
    rd_cycle[24170] = 1'b1;  wr_cycle[24170] = 1'b0;  addr_rom[24170]='h000039a8;  wr_data_rom[24170]='h00000000;
    rd_cycle[24171] = 1'b1;  wr_cycle[24171] = 1'b0;  addr_rom[24171]='h000039ac;  wr_data_rom[24171]='h00000000;
    rd_cycle[24172] = 1'b1;  wr_cycle[24172] = 1'b0;  addr_rom[24172]='h000039b0;  wr_data_rom[24172]='h00000000;
    rd_cycle[24173] = 1'b1;  wr_cycle[24173] = 1'b0;  addr_rom[24173]='h000039b4;  wr_data_rom[24173]='h00000000;
    rd_cycle[24174] = 1'b1;  wr_cycle[24174] = 1'b0;  addr_rom[24174]='h000039b8;  wr_data_rom[24174]='h00000000;
    rd_cycle[24175] = 1'b1;  wr_cycle[24175] = 1'b0;  addr_rom[24175]='h000039bc;  wr_data_rom[24175]='h00000000;
    rd_cycle[24176] = 1'b1;  wr_cycle[24176] = 1'b0;  addr_rom[24176]='h000039c0;  wr_data_rom[24176]='h00000000;
    rd_cycle[24177] = 1'b1;  wr_cycle[24177] = 1'b0;  addr_rom[24177]='h000039c4;  wr_data_rom[24177]='h00000000;
    rd_cycle[24178] = 1'b1;  wr_cycle[24178] = 1'b0;  addr_rom[24178]='h000039c8;  wr_data_rom[24178]='h00000000;
    rd_cycle[24179] = 1'b1;  wr_cycle[24179] = 1'b0;  addr_rom[24179]='h000039cc;  wr_data_rom[24179]='h00000000;
    rd_cycle[24180] = 1'b1;  wr_cycle[24180] = 1'b0;  addr_rom[24180]='h000039d0;  wr_data_rom[24180]='h00000000;
    rd_cycle[24181] = 1'b1;  wr_cycle[24181] = 1'b0;  addr_rom[24181]='h000039d4;  wr_data_rom[24181]='h00000000;
    rd_cycle[24182] = 1'b1;  wr_cycle[24182] = 1'b0;  addr_rom[24182]='h000039d8;  wr_data_rom[24182]='h00000000;
    rd_cycle[24183] = 1'b1;  wr_cycle[24183] = 1'b0;  addr_rom[24183]='h000039dc;  wr_data_rom[24183]='h00000000;
    rd_cycle[24184] = 1'b1;  wr_cycle[24184] = 1'b0;  addr_rom[24184]='h000039e0;  wr_data_rom[24184]='h00000000;
    rd_cycle[24185] = 1'b1;  wr_cycle[24185] = 1'b0;  addr_rom[24185]='h000039e4;  wr_data_rom[24185]='h00000000;
    rd_cycle[24186] = 1'b1;  wr_cycle[24186] = 1'b0;  addr_rom[24186]='h000039e8;  wr_data_rom[24186]='h00000000;
    rd_cycle[24187] = 1'b1;  wr_cycle[24187] = 1'b0;  addr_rom[24187]='h000039ec;  wr_data_rom[24187]='h00000000;
    rd_cycle[24188] = 1'b1;  wr_cycle[24188] = 1'b0;  addr_rom[24188]='h000039f0;  wr_data_rom[24188]='h00000000;
    rd_cycle[24189] = 1'b1;  wr_cycle[24189] = 1'b0;  addr_rom[24189]='h000039f4;  wr_data_rom[24189]='h00000000;
    rd_cycle[24190] = 1'b1;  wr_cycle[24190] = 1'b0;  addr_rom[24190]='h000039f8;  wr_data_rom[24190]='h00000000;
    rd_cycle[24191] = 1'b1;  wr_cycle[24191] = 1'b0;  addr_rom[24191]='h000039fc;  wr_data_rom[24191]='h00000000;
    rd_cycle[24192] = 1'b1;  wr_cycle[24192] = 1'b0;  addr_rom[24192]='h00003a00;  wr_data_rom[24192]='h00000000;
    rd_cycle[24193] = 1'b1;  wr_cycle[24193] = 1'b0;  addr_rom[24193]='h00003a04;  wr_data_rom[24193]='h00000000;
    rd_cycle[24194] = 1'b1;  wr_cycle[24194] = 1'b0;  addr_rom[24194]='h00003a08;  wr_data_rom[24194]='h00000000;
    rd_cycle[24195] = 1'b1;  wr_cycle[24195] = 1'b0;  addr_rom[24195]='h00003a0c;  wr_data_rom[24195]='h00000000;
    rd_cycle[24196] = 1'b1;  wr_cycle[24196] = 1'b0;  addr_rom[24196]='h00003a10;  wr_data_rom[24196]='h00000000;
    rd_cycle[24197] = 1'b1;  wr_cycle[24197] = 1'b0;  addr_rom[24197]='h00003a14;  wr_data_rom[24197]='h00000000;
    rd_cycle[24198] = 1'b1;  wr_cycle[24198] = 1'b0;  addr_rom[24198]='h00003a18;  wr_data_rom[24198]='h00000000;
    rd_cycle[24199] = 1'b1;  wr_cycle[24199] = 1'b0;  addr_rom[24199]='h00003a1c;  wr_data_rom[24199]='h00000000;
    rd_cycle[24200] = 1'b1;  wr_cycle[24200] = 1'b0;  addr_rom[24200]='h00003a20;  wr_data_rom[24200]='h00000000;
    rd_cycle[24201] = 1'b1;  wr_cycle[24201] = 1'b0;  addr_rom[24201]='h00003a24;  wr_data_rom[24201]='h00000000;
    rd_cycle[24202] = 1'b1;  wr_cycle[24202] = 1'b0;  addr_rom[24202]='h00003a28;  wr_data_rom[24202]='h00000000;
    rd_cycle[24203] = 1'b1;  wr_cycle[24203] = 1'b0;  addr_rom[24203]='h00003a2c;  wr_data_rom[24203]='h00000000;
    rd_cycle[24204] = 1'b1;  wr_cycle[24204] = 1'b0;  addr_rom[24204]='h00003a30;  wr_data_rom[24204]='h00000000;
    rd_cycle[24205] = 1'b1;  wr_cycle[24205] = 1'b0;  addr_rom[24205]='h00003a34;  wr_data_rom[24205]='h00000000;
    rd_cycle[24206] = 1'b1;  wr_cycle[24206] = 1'b0;  addr_rom[24206]='h00003a38;  wr_data_rom[24206]='h00000000;
    rd_cycle[24207] = 1'b1;  wr_cycle[24207] = 1'b0;  addr_rom[24207]='h00003a3c;  wr_data_rom[24207]='h00000000;
    rd_cycle[24208] = 1'b1;  wr_cycle[24208] = 1'b0;  addr_rom[24208]='h00003a40;  wr_data_rom[24208]='h00000000;
    rd_cycle[24209] = 1'b1;  wr_cycle[24209] = 1'b0;  addr_rom[24209]='h00003a44;  wr_data_rom[24209]='h00000000;
    rd_cycle[24210] = 1'b1;  wr_cycle[24210] = 1'b0;  addr_rom[24210]='h00003a48;  wr_data_rom[24210]='h00000000;
    rd_cycle[24211] = 1'b1;  wr_cycle[24211] = 1'b0;  addr_rom[24211]='h00003a4c;  wr_data_rom[24211]='h00000000;
    rd_cycle[24212] = 1'b1;  wr_cycle[24212] = 1'b0;  addr_rom[24212]='h00003a50;  wr_data_rom[24212]='h00000000;
    rd_cycle[24213] = 1'b1;  wr_cycle[24213] = 1'b0;  addr_rom[24213]='h00003a54;  wr_data_rom[24213]='h00000000;
    rd_cycle[24214] = 1'b1;  wr_cycle[24214] = 1'b0;  addr_rom[24214]='h00003a58;  wr_data_rom[24214]='h00000000;
    rd_cycle[24215] = 1'b1;  wr_cycle[24215] = 1'b0;  addr_rom[24215]='h00003a5c;  wr_data_rom[24215]='h00000000;
    rd_cycle[24216] = 1'b1;  wr_cycle[24216] = 1'b0;  addr_rom[24216]='h00003a60;  wr_data_rom[24216]='h00000000;
    rd_cycle[24217] = 1'b1;  wr_cycle[24217] = 1'b0;  addr_rom[24217]='h00003a64;  wr_data_rom[24217]='h00000000;
    rd_cycle[24218] = 1'b1;  wr_cycle[24218] = 1'b0;  addr_rom[24218]='h00003a68;  wr_data_rom[24218]='h00000000;
    rd_cycle[24219] = 1'b1;  wr_cycle[24219] = 1'b0;  addr_rom[24219]='h00003a6c;  wr_data_rom[24219]='h00000000;
    rd_cycle[24220] = 1'b1;  wr_cycle[24220] = 1'b0;  addr_rom[24220]='h00003a70;  wr_data_rom[24220]='h00000000;
    rd_cycle[24221] = 1'b1;  wr_cycle[24221] = 1'b0;  addr_rom[24221]='h00003a74;  wr_data_rom[24221]='h00000000;
    rd_cycle[24222] = 1'b1;  wr_cycle[24222] = 1'b0;  addr_rom[24222]='h00003a78;  wr_data_rom[24222]='h00000000;
    rd_cycle[24223] = 1'b1;  wr_cycle[24223] = 1'b0;  addr_rom[24223]='h00003a7c;  wr_data_rom[24223]='h00000000;
    rd_cycle[24224] = 1'b1;  wr_cycle[24224] = 1'b0;  addr_rom[24224]='h00003a80;  wr_data_rom[24224]='h00000000;
    rd_cycle[24225] = 1'b1;  wr_cycle[24225] = 1'b0;  addr_rom[24225]='h00003a84;  wr_data_rom[24225]='h00000000;
    rd_cycle[24226] = 1'b1;  wr_cycle[24226] = 1'b0;  addr_rom[24226]='h00003a88;  wr_data_rom[24226]='h00000000;
    rd_cycle[24227] = 1'b1;  wr_cycle[24227] = 1'b0;  addr_rom[24227]='h00003a8c;  wr_data_rom[24227]='h00000000;
    rd_cycle[24228] = 1'b1;  wr_cycle[24228] = 1'b0;  addr_rom[24228]='h00003a90;  wr_data_rom[24228]='h00000000;
    rd_cycle[24229] = 1'b1;  wr_cycle[24229] = 1'b0;  addr_rom[24229]='h00003a94;  wr_data_rom[24229]='h00000000;
    rd_cycle[24230] = 1'b1;  wr_cycle[24230] = 1'b0;  addr_rom[24230]='h00003a98;  wr_data_rom[24230]='h00000000;
    rd_cycle[24231] = 1'b1;  wr_cycle[24231] = 1'b0;  addr_rom[24231]='h00003a9c;  wr_data_rom[24231]='h00000000;
    rd_cycle[24232] = 1'b1;  wr_cycle[24232] = 1'b0;  addr_rom[24232]='h00003aa0;  wr_data_rom[24232]='h00000000;
    rd_cycle[24233] = 1'b1;  wr_cycle[24233] = 1'b0;  addr_rom[24233]='h00003aa4;  wr_data_rom[24233]='h00000000;
    rd_cycle[24234] = 1'b1;  wr_cycle[24234] = 1'b0;  addr_rom[24234]='h00003aa8;  wr_data_rom[24234]='h00000000;
    rd_cycle[24235] = 1'b1;  wr_cycle[24235] = 1'b0;  addr_rom[24235]='h00003aac;  wr_data_rom[24235]='h00000000;
    rd_cycle[24236] = 1'b1;  wr_cycle[24236] = 1'b0;  addr_rom[24236]='h00003ab0;  wr_data_rom[24236]='h00000000;
    rd_cycle[24237] = 1'b1;  wr_cycle[24237] = 1'b0;  addr_rom[24237]='h00003ab4;  wr_data_rom[24237]='h00000000;
    rd_cycle[24238] = 1'b1;  wr_cycle[24238] = 1'b0;  addr_rom[24238]='h00003ab8;  wr_data_rom[24238]='h00000000;
    rd_cycle[24239] = 1'b1;  wr_cycle[24239] = 1'b0;  addr_rom[24239]='h00003abc;  wr_data_rom[24239]='h00000000;
    rd_cycle[24240] = 1'b1;  wr_cycle[24240] = 1'b0;  addr_rom[24240]='h00003ac0;  wr_data_rom[24240]='h00000000;
    rd_cycle[24241] = 1'b1;  wr_cycle[24241] = 1'b0;  addr_rom[24241]='h00003ac4;  wr_data_rom[24241]='h00000000;
    rd_cycle[24242] = 1'b1;  wr_cycle[24242] = 1'b0;  addr_rom[24242]='h00003ac8;  wr_data_rom[24242]='h00000000;
    rd_cycle[24243] = 1'b1;  wr_cycle[24243] = 1'b0;  addr_rom[24243]='h00003acc;  wr_data_rom[24243]='h00000000;
    rd_cycle[24244] = 1'b1;  wr_cycle[24244] = 1'b0;  addr_rom[24244]='h00003ad0;  wr_data_rom[24244]='h00000000;
    rd_cycle[24245] = 1'b1;  wr_cycle[24245] = 1'b0;  addr_rom[24245]='h00003ad4;  wr_data_rom[24245]='h00000000;
    rd_cycle[24246] = 1'b1;  wr_cycle[24246] = 1'b0;  addr_rom[24246]='h00003ad8;  wr_data_rom[24246]='h00000000;
    rd_cycle[24247] = 1'b1;  wr_cycle[24247] = 1'b0;  addr_rom[24247]='h00003adc;  wr_data_rom[24247]='h00000000;
    rd_cycle[24248] = 1'b1;  wr_cycle[24248] = 1'b0;  addr_rom[24248]='h00003ae0;  wr_data_rom[24248]='h00000000;
    rd_cycle[24249] = 1'b1;  wr_cycle[24249] = 1'b0;  addr_rom[24249]='h00003ae4;  wr_data_rom[24249]='h00000000;
    rd_cycle[24250] = 1'b1;  wr_cycle[24250] = 1'b0;  addr_rom[24250]='h00003ae8;  wr_data_rom[24250]='h00000000;
    rd_cycle[24251] = 1'b1;  wr_cycle[24251] = 1'b0;  addr_rom[24251]='h00003aec;  wr_data_rom[24251]='h00000000;
    rd_cycle[24252] = 1'b1;  wr_cycle[24252] = 1'b0;  addr_rom[24252]='h00003af0;  wr_data_rom[24252]='h00000000;
    rd_cycle[24253] = 1'b1;  wr_cycle[24253] = 1'b0;  addr_rom[24253]='h00003af4;  wr_data_rom[24253]='h00000000;
    rd_cycle[24254] = 1'b1;  wr_cycle[24254] = 1'b0;  addr_rom[24254]='h00003af8;  wr_data_rom[24254]='h00000000;
    rd_cycle[24255] = 1'b1;  wr_cycle[24255] = 1'b0;  addr_rom[24255]='h00003afc;  wr_data_rom[24255]='h00000000;
    rd_cycle[24256] = 1'b1;  wr_cycle[24256] = 1'b0;  addr_rom[24256]='h00003b00;  wr_data_rom[24256]='h00000000;
    rd_cycle[24257] = 1'b1;  wr_cycle[24257] = 1'b0;  addr_rom[24257]='h00003b04;  wr_data_rom[24257]='h00000000;
    rd_cycle[24258] = 1'b1;  wr_cycle[24258] = 1'b0;  addr_rom[24258]='h00003b08;  wr_data_rom[24258]='h00000000;
    rd_cycle[24259] = 1'b1;  wr_cycle[24259] = 1'b0;  addr_rom[24259]='h00003b0c;  wr_data_rom[24259]='h00000000;
    rd_cycle[24260] = 1'b1;  wr_cycle[24260] = 1'b0;  addr_rom[24260]='h00003b10;  wr_data_rom[24260]='h00000000;
    rd_cycle[24261] = 1'b1;  wr_cycle[24261] = 1'b0;  addr_rom[24261]='h00003b14;  wr_data_rom[24261]='h00000000;
    rd_cycle[24262] = 1'b1;  wr_cycle[24262] = 1'b0;  addr_rom[24262]='h00003b18;  wr_data_rom[24262]='h00000000;
    rd_cycle[24263] = 1'b1;  wr_cycle[24263] = 1'b0;  addr_rom[24263]='h00003b1c;  wr_data_rom[24263]='h00000000;
    rd_cycle[24264] = 1'b1;  wr_cycle[24264] = 1'b0;  addr_rom[24264]='h00003b20;  wr_data_rom[24264]='h00000000;
    rd_cycle[24265] = 1'b1;  wr_cycle[24265] = 1'b0;  addr_rom[24265]='h00003b24;  wr_data_rom[24265]='h00000000;
    rd_cycle[24266] = 1'b1;  wr_cycle[24266] = 1'b0;  addr_rom[24266]='h00003b28;  wr_data_rom[24266]='h00000000;
    rd_cycle[24267] = 1'b1;  wr_cycle[24267] = 1'b0;  addr_rom[24267]='h00003b2c;  wr_data_rom[24267]='h00000000;
    rd_cycle[24268] = 1'b1;  wr_cycle[24268] = 1'b0;  addr_rom[24268]='h00003b30;  wr_data_rom[24268]='h00000000;
    rd_cycle[24269] = 1'b1;  wr_cycle[24269] = 1'b0;  addr_rom[24269]='h00003b34;  wr_data_rom[24269]='h00000000;
    rd_cycle[24270] = 1'b1;  wr_cycle[24270] = 1'b0;  addr_rom[24270]='h00003b38;  wr_data_rom[24270]='h00000000;
    rd_cycle[24271] = 1'b1;  wr_cycle[24271] = 1'b0;  addr_rom[24271]='h00003b3c;  wr_data_rom[24271]='h00000000;
    rd_cycle[24272] = 1'b1;  wr_cycle[24272] = 1'b0;  addr_rom[24272]='h00003b40;  wr_data_rom[24272]='h00000000;
    rd_cycle[24273] = 1'b1;  wr_cycle[24273] = 1'b0;  addr_rom[24273]='h00003b44;  wr_data_rom[24273]='h00000000;
    rd_cycle[24274] = 1'b1;  wr_cycle[24274] = 1'b0;  addr_rom[24274]='h00003b48;  wr_data_rom[24274]='h00000000;
    rd_cycle[24275] = 1'b1;  wr_cycle[24275] = 1'b0;  addr_rom[24275]='h00003b4c;  wr_data_rom[24275]='h00000000;
    rd_cycle[24276] = 1'b1;  wr_cycle[24276] = 1'b0;  addr_rom[24276]='h00003b50;  wr_data_rom[24276]='h00000000;
    rd_cycle[24277] = 1'b1;  wr_cycle[24277] = 1'b0;  addr_rom[24277]='h00003b54;  wr_data_rom[24277]='h00000000;
    rd_cycle[24278] = 1'b1;  wr_cycle[24278] = 1'b0;  addr_rom[24278]='h00003b58;  wr_data_rom[24278]='h00000000;
    rd_cycle[24279] = 1'b1;  wr_cycle[24279] = 1'b0;  addr_rom[24279]='h00003b5c;  wr_data_rom[24279]='h00000000;
    rd_cycle[24280] = 1'b1;  wr_cycle[24280] = 1'b0;  addr_rom[24280]='h00003b60;  wr_data_rom[24280]='h00000000;
    rd_cycle[24281] = 1'b1;  wr_cycle[24281] = 1'b0;  addr_rom[24281]='h00003b64;  wr_data_rom[24281]='h00000000;
    rd_cycle[24282] = 1'b1;  wr_cycle[24282] = 1'b0;  addr_rom[24282]='h00003b68;  wr_data_rom[24282]='h00000000;
    rd_cycle[24283] = 1'b1;  wr_cycle[24283] = 1'b0;  addr_rom[24283]='h00003b6c;  wr_data_rom[24283]='h00000000;
    rd_cycle[24284] = 1'b1;  wr_cycle[24284] = 1'b0;  addr_rom[24284]='h00003b70;  wr_data_rom[24284]='h00000000;
    rd_cycle[24285] = 1'b1;  wr_cycle[24285] = 1'b0;  addr_rom[24285]='h00003b74;  wr_data_rom[24285]='h00000000;
    rd_cycle[24286] = 1'b1;  wr_cycle[24286] = 1'b0;  addr_rom[24286]='h00003b78;  wr_data_rom[24286]='h00000000;
    rd_cycle[24287] = 1'b1;  wr_cycle[24287] = 1'b0;  addr_rom[24287]='h00003b7c;  wr_data_rom[24287]='h00000000;
    rd_cycle[24288] = 1'b1;  wr_cycle[24288] = 1'b0;  addr_rom[24288]='h00003b80;  wr_data_rom[24288]='h00000000;
    rd_cycle[24289] = 1'b1;  wr_cycle[24289] = 1'b0;  addr_rom[24289]='h00003b84;  wr_data_rom[24289]='h00000000;
    rd_cycle[24290] = 1'b1;  wr_cycle[24290] = 1'b0;  addr_rom[24290]='h00003b88;  wr_data_rom[24290]='h00000000;
    rd_cycle[24291] = 1'b1;  wr_cycle[24291] = 1'b0;  addr_rom[24291]='h00003b8c;  wr_data_rom[24291]='h00000000;
    rd_cycle[24292] = 1'b1;  wr_cycle[24292] = 1'b0;  addr_rom[24292]='h00003b90;  wr_data_rom[24292]='h00000000;
    rd_cycle[24293] = 1'b1;  wr_cycle[24293] = 1'b0;  addr_rom[24293]='h00003b94;  wr_data_rom[24293]='h00000000;
    rd_cycle[24294] = 1'b1;  wr_cycle[24294] = 1'b0;  addr_rom[24294]='h00003b98;  wr_data_rom[24294]='h00000000;
    rd_cycle[24295] = 1'b1;  wr_cycle[24295] = 1'b0;  addr_rom[24295]='h00003b9c;  wr_data_rom[24295]='h00000000;
    rd_cycle[24296] = 1'b1;  wr_cycle[24296] = 1'b0;  addr_rom[24296]='h00003ba0;  wr_data_rom[24296]='h00000000;
    rd_cycle[24297] = 1'b1;  wr_cycle[24297] = 1'b0;  addr_rom[24297]='h00003ba4;  wr_data_rom[24297]='h00000000;
    rd_cycle[24298] = 1'b1;  wr_cycle[24298] = 1'b0;  addr_rom[24298]='h00003ba8;  wr_data_rom[24298]='h00000000;
    rd_cycle[24299] = 1'b1;  wr_cycle[24299] = 1'b0;  addr_rom[24299]='h00003bac;  wr_data_rom[24299]='h00000000;
    rd_cycle[24300] = 1'b1;  wr_cycle[24300] = 1'b0;  addr_rom[24300]='h00003bb0;  wr_data_rom[24300]='h00000000;
    rd_cycle[24301] = 1'b1;  wr_cycle[24301] = 1'b0;  addr_rom[24301]='h00003bb4;  wr_data_rom[24301]='h00000000;
    rd_cycle[24302] = 1'b1;  wr_cycle[24302] = 1'b0;  addr_rom[24302]='h00003bb8;  wr_data_rom[24302]='h00000000;
    rd_cycle[24303] = 1'b1;  wr_cycle[24303] = 1'b0;  addr_rom[24303]='h00003bbc;  wr_data_rom[24303]='h00000000;
    rd_cycle[24304] = 1'b1;  wr_cycle[24304] = 1'b0;  addr_rom[24304]='h00003bc0;  wr_data_rom[24304]='h00000000;
    rd_cycle[24305] = 1'b1;  wr_cycle[24305] = 1'b0;  addr_rom[24305]='h00003bc4;  wr_data_rom[24305]='h00000000;
    rd_cycle[24306] = 1'b1;  wr_cycle[24306] = 1'b0;  addr_rom[24306]='h00003bc8;  wr_data_rom[24306]='h00000000;
    rd_cycle[24307] = 1'b1;  wr_cycle[24307] = 1'b0;  addr_rom[24307]='h00003bcc;  wr_data_rom[24307]='h00000000;
    rd_cycle[24308] = 1'b1;  wr_cycle[24308] = 1'b0;  addr_rom[24308]='h00003bd0;  wr_data_rom[24308]='h00000000;
    rd_cycle[24309] = 1'b1;  wr_cycle[24309] = 1'b0;  addr_rom[24309]='h00003bd4;  wr_data_rom[24309]='h00000000;
    rd_cycle[24310] = 1'b1;  wr_cycle[24310] = 1'b0;  addr_rom[24310]='h00003bd8;  wr_data_rom[24310]='h00000000;
    rd_cycle[24311] = 1'b1;  wr_cycle[24311] = 1'b0;  addr_rom[24311]='h00003bdc;  wr_data_rom[24311]='h00000000;
    rd_cycle[24312] = 1'b1;  wr_cycle[24312] = 1'b0;  addr_rom[24312]='h00003be0;  wr_data_rom[24312]='h00000000;
    rd_cycle[24313] = 1'b1;  wr_cycle[24313] = 1'b0;  addr_rom[24313]='h00003be4;  wr_data_rom[24313]='h00000000;
    rd_cycle[24314] = 1'b1;  wr_cycle[24314] = 1'b0;  addr_rom[24314]='h00003be8;  wr_data_rom[24314]='h00000000;
    rd_cycle[24315] = 1'b1;  wr_cycle[24315] = 1'b0;  addr_rom[24315]='h00003bec;  wr_data_rom[24315]='h00000000;
    rd_cycle[24316] = 1'b1;  wr_cycle[24316] = 1'b0;  addr_rom[24316]='h00003bf0;  wr_data_rom[24316]='h00000000;
    rd_cycle[24317] = 1'b1;  wr_cycle[24317] = 1'b0;  addr_rom[24317]='h00003bf4;  wr_data_rom[24317]='h00000000;
    rd_cycle[24318] = 1'b1;  wr_cycle[24318] = 1'b0;  addr_rom[24318]='h00003bf8;  wr_data_rom[24318]='h00000000;
    rd_cycle[24319] = 1'b1;  wr_cycle[24319] = 1'b0;  addr_rom[24319]='h00003bfc;  wr_data_rom[24319]='h00000000;
    rd_cycle[24320] = 1'b1;  wr_cycle[24320] = 1'b0;  addr_rom[24320]='h00003c00;  wr_data_rom[24320]='h00000000;
    rd_cycle[24321] = 1'b1;  wr_cycle[24321] = 1'b0;  addr_rom[24321]='h00003c04;  wr_data_rom[24321]='h00000000;
    rd_cycle[24322] = 1'b1;  wr_cycle[24322] = 1'b0;  addr_rom[24322]='h00003c08;  wr_data_rom[24322]='h00000000;
    rd_cycle[24323] = 1'b1;  wr_cycle[24323] = 1'b0;  addr_rom[24323]='h00003c0c;  wr_data_rom[24323]='h00000000;
    rd_cycle[24324] = 1'b1;  wr_cycle[24324] = 1'b0;  addr_rom[24324]='h00003c10;  wr_data_rom[24324]='h00000000;
    rd_cycle[24325] = 1'b1;  wr_cycle[24325] = 1'b0;  addr_rom[24325]='h00003c14;  wr_data_rom[24325]='h00000000;
    rd_cycle[24326] = 1'b1;  wr_cycle[24326] = 1'b0;  addr_rom[24326]='h00003c18;  wr_data_rom[24326]='h00000000;
    rd_cycle[24327] = 1'b1;  wr_cycle[24327] = 1'b0;  addr_rom[24327]='h00003c1c;  wr_data_rom[24327]='h00000000;
    rd_cycle[24328] = 1'b1;  wr_cycle[24328] = 1'b0;  addr_rom[24328]='h00003c20;  wr_data_rom[24328]='h00000000;
    rd_cycle[24329] = 1'b1;  wr_cycle[24329] = 1'b0;  addr_rom[24329]='h00003c24;  wr_data_rom[24329]='h00000000;
    rd_cycle[24330] = 1'b1;  wr_cycle[24330] = 1'b0;  addr_rom[24330]='h00003c28;  wr_data_rom[24330]='h00000000;
    rd_cycle[24331] = 1'b1;  wr_cycle[24331] = 1'b0;  addr_rom[24331]='h00003c2c;  wr_data_rom[24331]='h00000000;
    rd_cycle[24332] = 1'b1;  wr_cycle[24332] = 1'b0;  addr_rom[24332]='h00003c30;  wr_data_rom[24332]='h00000000;
    rd_cycle[24333] = 1'b1;  wr_cycle[24333] = 1'b0;  addr_rom[24333]='h00003c34;  wr_data_rom[24333]='h00000000;
    rd_cycle[24334] = 1'b1;  wr_cycle[24334] = 1'b0;  addr_rom[24334]='h00003c38;  wr_data_rom[24334]='h00000000;
    rd_cycle[24335] = 1'b1;  wr_cycle[24335] = 1'b0;  addr_rom[24335]='h00003c3c;  wr_data_rom[24335]='h00000000;
    rd_cycle[24336] = 1'b1;  wr_cycle[24336] = 1'b0;  addr_rom[24336]='h00003c40;  wr_data_rom[24336]='h00000000;
    rd_cycle[24337] = 1'b1;  wr_cycle[24337] = 1'b0;  addr_rom[24337]='h00003c44;  wr_data_rom[24337]='h00000000;
    rd_cycle[24338] = 1'b1;  wr_cycle[24338] = 1'b0;  addr_rom[24338]='h00003c48;  wr_data_rom[24338]='h00000000;
    rd_cycle[24339] = 1'b1;  wr_cycle[24339] = 1'b0;  addr_rom[24339]='h00003c4c;  wr_data_rom[24339]='h00000000;
    rd_cycle[24340] = 1'b1;  wr_cycle[24340] = 1'b0;  addr_rom[24340]='h00003c50;  wr_data_rom[24340]='h00000000;
    rd_cycle[24341] = 1'b1;  wr_cycle[24341] = 1'b0;  addr_rom[24341]='h00003c54;  wr_data_rom[24341]='h00000000;
    rd_cycle[24342] = 1'b1;  wr_cycle[24342] = 1'b0;  addr_rom[24342]='h00003c58;  wr_data_rom[24342]='h00000000;
    rd_cycle[24343] = 1'b1;  wr_cycle[24343] = 1'b0;  addr_rom[24343]='h00003c5c;  wr_data_rom[24343]='h00000000;
    rd_cycle[24344] = 1'b1;  wr_cycle[24344] = 1'b0;  addr_rom[24344]='h00003c60;  wr_data_rom[24344]='h00000000;
    rd_cycle[24345] = 1'b1;  wr_cycle[24345] = 1'b0;  addr_rom[24345]='h00003c64;  wr_data_rom[24345]='h00000000;
    rd_cycle[24346] = 1'b1;  wr_cycle[24346] = 1'b0;  addr_rom[24346]='h00003c68;  wr_data_rom[24346]='h00000000;
    rd_cycle[24347] = 1'b1;  wr_cycle[24347] = 1'b0;  addr_rom[24347]='h00003c6c;  wr_data_rom[24347]='h00000000;
    rd_cycle[24348] = 1'b1;  wr_cycle[24348] = 1'b0;  addr_rom[24348]='h00003c70;  wr_data_rom[24348]='h00000000;
    rd_cycle[24349] = 1'b1;  wr_cycle[24349] = 1'b0;  addr_rom[24349]='h00003c74;  wr_data_rom[24349]='h00000000;
    rd_cycle[24350] = 1'b1;  wr_cycle[24350] = 1'b0;  addr_rom[24350]='h00003c78;  wr_data_rom[24350]='h00000000;
    rd_cycle[24351] = 1'b1;  wr_cycle[24351] = 1'b0;  addr_rom[24351]='h00003c7c;  wr_data_rom[24351]='h00000000;
    rd_cycle[24352] = 1'b1;  wr_cycle[24352] = 1'b0;  addr_rom[24352]='h00003c80;  wr_data_rom[24352]='h00000000;
    rd_cycle[24353] = 1'b1;  wr_cycle[24353] = 1'b0;  addr_rom[24353]='h00003c84;  wr_data_rom[24353]='h00000000;
    rd_cycle[24354] = 1'b1;  wr_cycle[24354] = 1'b0;  addr_rom[24354]='h00003c88;  wr_data_rom[24354]='h00000000;
    rd_cycle[24355] = 1'b1;  wr_cycle[24355] = 1'b0;  addr_rom[24355]='h00003c8c;  wr_data_rom[24355]='h00000000;
    rd_cycle[24356] = 1'b1;  wr_cycle[24356] = 1'b0;  addr_rom[24356]='h00003c90;  wr_data_rom[24356]='h00000000;
    rd_cycle[24357] = 1'b1;  wr_cycle[24357] = 1'b0;  addr_rom[24357]='h00003c94;  wr_data_rom[24357]='h00000000;
    rd_cycle[24358] = 1'b1;  wr_cycle[24358] = 1'b0;  addr_rom[24358]='h00003c98;  wr_data_rom[24358]='h00000000;
    rd_cycle[24359] = 1'b1;  wr_cycle[24359] = 1'b0;  addr_rom[24359]='h00003c9c;  wr_data_rom[24359]='h00000000;
    rd_cycle[24360] = 1'b1;  wr_cycle[24360] = 1'b0;  addr_rom[24360]='h00003ca0;  wr_data_rom[24360]='h00000000;
    rd_cycle[24361] = 1'b1;  wr_cycle[24361] = 1'b0;  addr_rom[24361]='h00003ca4;  wr_data_rom[24361]='h00000000;
    rd_cycle[24362] = 1'b1;  wr_cycle[24362] = 1'b0;  addr_rom[24362]='h00003ca8;  wr_data_rom[24362]='h00000000;
    rd_cycle[24363] = 1'b1;  wr_cycle[24363] = 1'b0;  addr_rom[24363]='h00003cac;  wr_data_rom[24363]='h00000000;
    rd_cycle[24364] = 1'b1;  wr_cycle[24364] = 1'b0;  addr_rom[24364]='h00003cb0;  wr_data_rom[24364]='h00000000;
    rd_cycle[24365] = 1'b1;  wr_cycle[24365] = 1'b0;  addr_rom[24365]='h00003cb4;  wr_data_rom[24365]='h00000000;
    rd_cycle[24366] = 1'b1;  wr_cycle[24366] = 1'b0;  addr_rom[24366]='h00003cb8;  wr_data_rom[24366]='h00000000;
    rd_cycle[24367] = 1'b1;  wr_cycle[24367] = 1'b0;  addr_rom[24367]='h00003cbc;  wr_data_rom[24367]='h00000000;
    rd_cycle[24368] = 1'b1;  wr_cycle[24368] = 1'b0;  addr_rom[24368]='h00003cc0;  wr_data_rom[24368]='h00000000;
    rd_cycle[24369] = 1'b1;  wr_cycle[24369] = 1'b0;  addr_rom[24369]='h00003cc4;  wr_data_rom[24369]='h00000000;
    rd_cycle[24370] = 1'b1;  wr_cycle[24370] = 1'b0;  addr_rom[24370]='h00003cc8;  wr_data_rom[24370]='h00000000;
    rd_cycle[24371] = 1'b1;  wr_cycle[24371] = 1'b0;  addr_rom[24371]='h00003ccc;  wr_data_rom[24371]='h00000000;
    rd_cycle[24372] = 1'b1;  wr_cycle[24372] = 1'b0;  addr_rom[24372]='h00003cd0;  wr_data_rom[24372]='h00000000;
    rd_cycle[24373] = 1'b1;  wr_cycle[24373] = 1'b0;  addr_rom[24373]='h00003cd4;  wr_data_rom[24373]='h00000000;
    rd_cycle[24374] = 1'b1;  wr_cycle[24374] = 1'b0;  addr_rom[24374]='h00003cd8;  wr_data_rom[24374]='h00000000;
    rd_cycle[24375] = 1'b1;  wr_cycle[24375] = 1'b0;  addr_rom[24375]='h00003cdc;  wr_data_rom[24375]='h00000000;
    rd_cycle[24376] = 1'b1;  wr_cycle[24376] = 1'b0;  addr_rom[24376]='h00003ce0;  wr_data_rom[24376]='h00000000;
    rd_cycle[24377] = 1'b1;  wr_cycle[24377] = 1'b0;  addr_rom[24377]='h00003ce4;  wr_data_rom[24377]='h00000000;
    rd_cycle[24378] = 1'b1;  wr_cycle[24378] = 1'b0;  addr_rom[24378]='h00003ce8;  wr_data_rom[24378]='h00000000;
    rd_cycle[24379] = 1'b1;  wr_cycle[24379] = 1'b0;  addr_rom[24379]='h00003cec;  wr_data_rom[24379]='h00000000;
    rd_cycle[24380] = 1'b1;  wr_cycle[24380] = 1'b0;  addr_rom[24380]='h00003cf0;  wr_data_rom[24380]='h00000000;
    rd_cycle[24381] = 1'b1;  wr_cycle[24381] = 1'b0;  addr_rom[24381]='h00003cf4;  wr_data_rom[24381]='h00000000;
    rd_cycle[24382] = 1'b1;  wr_cycle[24382] = 1'b0;  addr_rom[24382]='h00003cf8;  wr_data_rom[24382]='h00000000;
    rd_cycle[24383] = 1'b1;  wr_cycle[24383] = 1'b0;  addr_rom[24383]='h00003cfc;  wr_data_rom[24383]='h00000000;
    rd_cycle[24384] = 1'b1;  wr_cycle[24384] = 1'b0;  addr_rom[24384]='h00003d00;  wr_data_rom[24384]='h00000000;
    rd_cycle[24385] = 1'b1;  wr_cycle[24385] = 1'b0;  addr_rom[24385]='h00003d04;  wr_data_rom[24385]='h00000000;
    rd_cycle[24386] = 1'b1;  wr_cycle[24386] = 1'b0;  addr_rom[24386]='h00003d08;  wr_data_rom[24386]='h00000000;
    rd_cycle[24387] = 1'b1;  wr_cycle[24387] = 1'b0;  addr_rom[24387]='h00003d0c;  wr_data_rom[24387]='h00000000;
    rd_cycle[24388] = 1'b1;  wr_cycle[24388] = 1'b0;  addr_rom[24388]='h00003d10;  wr_data_rom[24388]='h00000000;
    rd_cycle[24389] = 1'b1;  wr_cycle[24389] = 1'b0;  addr_rom[24389]='h00003d14;  wr_data_rom[24389]='h00000000;
    rd_cycle[24390] = 1'b1;  wr_cycle[24390] = 1'b0;  addr_rom[24390]='h00003d18;  wr_data_rom[24390]='h00000000;
    rd_cycle[24391] = 1'b1;  wr_cycle[24391] = 1'b0;  addr_rom[24391]='h00003d1c;  wr_data_rom[24391]='h00000000;
    rd_cycle[24392] = 1'b1;  wr_cycle[24392] = 1'b0;  addr_rom[24392]='h00003d20;  wr_data_rom[24392]='h00000000;
    rd_cycle[24393] = 1'b1;  wr_cycle[24393] = 1'b0;  addr_rom[24393]='h00003d24;  wr_data_rom[24393]='h00000000;
    rd_cycle[24394] = 1'b1;  wr_cycle[24394] = 1'b0;  addr_rom[24394]='h00003d28;  wr_data_rom[24394]='h00000000;
    rd_cycle[24395] = 1'b1;  wr_cycle[24395] = 1'b0;  addr_rom[24395]='h00003d2c;  wr_data_rom[24395]='h00000000;
    rd_cycle[24396] = 1'b1;  wr_cycle[24396] = 1'b0;  addr_rom[24396]='h00003d30;  wr_data_rom[24396]='h00000000;
    rd_cycle[24397] = 1'b1;  wr_cycle[24397] = 1'b0;  addr_rom[24397]='h00003d34;  wr_data_rom[24397]='h00000000;
    rd_cycle[24398] = 1'b1;  wr_cycle[24398] = 1'b0;  addr_rom[24398]='h00003d38;  wr_data_rom[24398]='h00000000;
    rd_cycle[24399] = 1'b1;  wr_cycle[24399] = 1'b0;  addr_rom[24399]='h00003d3c;  wr_data_rom[24399]='h00000000;
    rd_cycle[24400] = 1'b1;  wr_cycle[24400] = 1'b0;  addr_rom[24400]='h00003d40;  wr_data_rom[24400]='h00000000;
    rd_cycle[24401] = 1'b1;  wr_cycle[24401] = 1'b0;  addr_rom[24401]='h00003d44;  wr_data_rom[24401]='h00000000;
    rd_cycle[24402] = 1'b1;  wr_cycle[24402] = 1'b0;  addr_rom[24402]='h00003d48;  wr_data_rom[24402]='h00000000;
    rd_cycle[24403] = 1'b1;  wr_cycle[24403] = 1'b0;  addr_rom[24403]='h00003d4c;  wr_data_rom[24403]='h00000000;
    rd_cycle[24404] = 1'b1;  wr_cycle[24404] = 1'b0;  addr_rom[24404]='h00003d50;  wr_data_rom[24404]='h00000000;
    rd_cycle[24405] = 1'b1;  wr_cycle[24405] = 1'b0;  addr_rom[24405]='h00003d54;  wr_data_rom[24405]='h00000000;
    rd_cycle[24406] = 1'b1;  wr_cycle[24406] = 1'b0;  addr_rom[24406]='h00003d58;  wr_data_rom[24406]='h00000000;
    rd_cycle[24407] = 1'b1;  wr_cycle[24407] = 1'b0;  addr_rom[24407]='h00003d5c;  wr_data_rom[24407]='h00000000;
    rd_cycle[24408] = 1'b1;  wr_cycle[24408] = 1'b0;  addr_rom[24408]='h00003d60;  wr_data_rom[24408]='h00000000;
    rd_cycle[24409] = 1'b1;  wr_cycle[24409] = 1'b0;  addr_rom[24409]='h00003d64;  wr_data_rom[24409]='h00000000;
    rd_cycle[24410] = 1'b1;  wr_cycle[24410] = 1'b0;  addr_rom[24410]='h00003d68;  wr_data_rom[24410]='h00000000;
    rd_cycle[24411] = 1'b1;  wr_cycle[24411] = 1'b0;  addr_rom[24411]='h00003d6c;  wr_data_rom[24411]='h00000000;
    rd_cycle[24412] = 1'b1;  wr_cycle[24412] = 1'b0;  addr_rom[24412]='h00003d70;  wr_data_rom[24412]='h00000000;
    rd_cycle[24413] = 1'b1;  wr_cycle[24413] = 1'b0;  addr_rom[24413]='h00003d74;  wr_data_rom[24413]='h00000000;
    rd_cycle[24414] = 1'b1;  wr_cycle[24414] = 1'b0;  addr_rom[24414]='h00003d78;  wr_data_rom[24414]='h00000000;
    rd_cycle[24415] = 1'b1;  wr_cycle[24415] = 1'b0;  addr_rom[24415]='h00003d7c;  wr_data_rom[24415]='h00000000;
    rd_cycle[24416] = 1'b1;  wr_cycle[24416] = 1'b0;  addr_rom[24416]='h00003d80;  wr_data_rom[24416]='h00000000;
    rd_cycle[24417] = 1'b1;  wr_cycle[24417] = 1'b0;  addr_rom[24417]='h00003d84;  wr_data_rom[24417]='h00000000;
    rd_cycle[24418] = 1'b1;  wr_cycle[24418] = 1'b0;  addr_rom[24418]='h00003d88;  wr_data_rom[24418]='h00000000;
    rd_cycle[24419] = 1'b1;  wr_cycle[24419] = 1'b0;  addr_rom[24419]='h00003d8c;  wr_data_rom[24419]='h00000000;
    rd_cycle[24420] = 1'b1;  wr_cycle[24420] = 1'b0;  addr_rom[24420]='h00003d90;  wr_data_rom[24420]='h00000000;
    rd_cycle[24421] = 1'b1;  wr_cycle[24421] = 1'b0;  addr_rom[24421]='h00003d94;  wr_data_rom[24421]='h00000000;
    rd_cycle[24422] = 1'b1;  wr_cycle[24422] = 1'b0;  addr_rom[24422]='h00003d98;  wr_data_rom[24422]='h00000000;
    rd_cycle[24423] = 1'b1;  wr_cycle[24423] = 1'b0;  addr_rom[24423]='h00003d9c;  wr_data_rom[24423]='h00000000;
    rd_cycle[24424] = 1'b1;  wr_cycle[24424] = 1'b0;  addr_rom[24424]='h00003da0;  wr_data_rom[24424]='h00000000;
    rd_cycle[24425] = 1'b1;  wr_cycle[24425] = 1'b0;  addr_rom[24425]='h00003da4;  wr_data_rom[24425]='h00000000;
    rd_cycle[24426] = 1'b1;  wr_cycle[24426] = 1'b0;  addr_rom[24426]='h00003da8;  wr_data_rom[24426]='h00000000;
    rd_cycle[24427] = 1'b1;  wr_cycle[24427] = 1'b0;  addr_rom[24427]='h00003dac;  wr_data_rom[24427]='h00000000;
    rd_cycle[24428] = 1'b1;  wr_cycle[24428] = 1'b0;  addr_rom[24428]='h00003db0;  wr_data_rom[24428]='h00000000;
    rd_cycle[24429] = 1'b1;  wr_cycle[24429] = 1'b0;  addr_rom[24429]='h00003db4;  wr_data_rom[24429]='h00000000;
    rd_cycle[24430] = 1'b1;  wr_cycle[24430] = 1'b0;  addr_rom[24430]='h00003db8;  wr_data_rom[24430]='h00000000;
    rd_cycle[24431] = 1'b1;  wr_cycle[24431] = 1'b0;  addr_rom[24431]='h00003dbc;  wr_data_rom[24431]='h00000000;
    rd_cycle[24432] = 1'b1;  wr_cycle[24432] = 1'b0;  addr_rom[24432]='h00003dc0;  wr_data_rom[24432]='h00000000;
    rd_cycle[24433] = 1'b1;  wr_cycle[24433] = 1'b0;  addr_rom[24433]='h00003dc4;  wr_data_rom[24433]='h00000000;
    rd_cycle[24434] = 1'b1;  wr_cycle[24434] = 1'b0;  addr_rom[24434]='h00003dc8;  wr_data_rom[24434]='h00000000;
    rd_cycle[24435] = 1'b1;  wr_cycle[24435] = 1'b0;  addr_rom[24435]='h00003dcc;  wr_data_rom[24435]='h00000000;
    rd_cycle[24436] = 1'b1;  wr_cycle[24436] = 1'b0;  addr_rom[24436]='h00003dd0;  wr_data_rom[24436]='h00000000;
    rd_cycle[24437] = 1'b1;  wr_cycle[24437] = 1'b0;  addr_rom[24437]='h00003dd4;  wr_data_rom[24437]='h00000000;
    rd_cycle[24438] = 1'b1;  wr_cycle[24438] = 1'b0;  addr_rom[24438]='h00003dd8;  wr_data_rom[24438]='h00000000;
    rd_cycle[24439] = 1'b1;  wr_cycle[24439] = 1'b0;  addr_rom[24439]='h00003ddc;  wr_data_rom[24439]='h00000000;
    rd_cycle[24440] = 1'b1;  wr_cycle[24440] = 1'b0;  addr_rom[24440]='h00003de0;  wr_data_rom[24440]='h00000000;
    rd_cycle[24441] = 1'b1;  wr_cycle[24441] = 1'b0;  addr_rom[24441]='h00003de4;  wr_data_rom[24441]='h00000000;
    rd_cycle[24442] = 1'b1;  wr_cycle[24442] = 1'b0;  addr_rom[24442]='h00003de8;  wr_data_rom[24442]='h00000000;
    rd_cycle[24443] = 1'b1;  wr_cycle[24443] = 1'b0;  addr_rom[24443]='h00003dec;  wr_data_rom[24443]='h00000000;
    rd_cycle[24444] = 1'b1;  wr_cycle[24444] = 1'b0;  addr_rom[24444]='h00003df0;  wr_data_rom[24444]='h00000000;
    rd_cycle[24445] = 1'b1;  wr_cycle[24445] = 1'b0;  addr_rom[24445]='h00003df4;  wr_data_rom[24445]='h00000000;
    rd_cycle[24446] = 1'b1;  wr_cycle[24446] = 1'b0;  addr_rom[24446]='h00003df8;  wr_data_rom[24446]='h00000000;
    rd_cycle[24447] = 1'b1;  wr_cycle[24447] = 1'b0;  addr_rom[24447]='h00003dfc;  wr_data_rom[24447]='h00000000;
    rd_cycle[24448] = 1'b1;  wr_cycle[24448] = 1'b0;  addr_rom[24448]='h00003e00;  wr_data_rom[24448]='h00000000;
    rd_cycle[24449] = 1'b1;  wr_cycle[24449] = 1'b0;  addr_rom[24449]='h00003e04;  wr_data_rom[24449]='h00000000;
    rd_cycle[24450] = 1'b1;  wr_cycle[24450] = 1'b0;  addr_rom[24450]='h00003e08;  wr_data_rom[24450]='h00000000;
    rd_cycle[24451] = 1'b1;  wr_cycle[24451] = 1'b0;  addr_rom[24451]='h00003e0c;  wr_data_rom[24451]='h00000000;
    rd_cycle[24452] = 1'b1;  wr_cycle[24452] = 1'b0;  addr_rom[24452]='h00003e10;  wr_data_rom[24452]='h00000000;
    rd_cycle[24453] = 1'b1;  wr_cycle[24453] = 1'b0;  addr_rom[24453]='h00003e14;  wr_data_rom[24453]='h00000000;
    rd_cycle[24454] = 1'b1;  wr_cycle[24454] = 1'b0;  addr_rom[24454]='h00003e18;  wr_data_rom[24454]='h00000000;
    rd_cycle[24455] = 1'b1;  wr_cycle[24455] = 1'b0;  addr_rom[24455]='h00003e1c;  wr_data_rom[24455]='h00000000;
    rd_cycle[24456] = 1'b1;  wr_cycle[24456] = 1'b0;  addr_rom[24456]='h00003e20;  wr_data_rom[24456]='h00000000;
    rd_cycle[24457] = 1'b1;  wr_cycle[24457] = 1'b0;  addr_rom[24457]='h00003e24;  wr_data_rom[24457]='h00000000;
    rd_cycle[24458] = 1'b1;  wr_cycle[24458] = 1'b0;  addr_rom[24458]='h00003e28;  wr_data_rom[24458]='h00000000;
    rd_cycle[24459] = 1'b1;  wr_cycle[24459] = 1'b0;  addr_rom[24459]='h00003e2c;  wr_data_rom[24459]='h00000000;
    rd_cycle[24460] = 1'b1;  wr_cycle[24460] = 1'b0;  addr_rom[24460]='h00003e30;  wr_data_rom[24460]='h00000000;
    rd_cycle[24461] = 1'b1;  wr_cycle[24461] = 1'b0;  addr_rom[24461]='h00003e34;  wr_data_rom[24461]='h00000000;
    rd_cycle[24462] = 1'b1;  wr_cycle[24462] = 1'b0;  addr_rom[24462]='h00003e38;  wr_data_rom[24462]='h00000000;
    rd_cycle[24463] = 1'b1;  wr_cycle[24463] = 1'b0;  addr_rom[24463]='h00003e3c;  wr_data_rom[24463]='h00000000;
    rd_cycle[24464] = 1'b1;  wr_cycle[24464] = 1'b0;  addr_rom[24464]='h00003e40;  wr_data_rom[24464]='h00000000;
    rd_cycle[24465] = 1'b1;  wr_cycle[24465] = 1'b0;  addr_rom[24465]='h00003e44;  wr_data_rom[24465]='h00000000;
    rd_cycle[24466] = 1'b1;  wr_cycle[24466] = 1'b0;  addr_rom[24466]='h00003e48;  wr_data_rom[24466]='h00000000;
    rd_cycle[24467] = 1'b1;  wr_cycle[24467] = 1'b0;  addr_rom[24467]='h00003e4c;  wr_data_rom[24467]='h00000000;
    rd_cycle[24468] = 1'b1;  wr_cycle[24468] = 1'b0;  addr_rom[24468]='h00003e50;  wr_data_rom[24468]='h00000000;
    rd_cycle[24469] = 1'b1;  wr_cycle[24469] = 1'b0;  addr_rom[24469]='h00003e54;  wr_data_rom[24469]='h00000000;
    rd_cycle[24470] = 1'b1;  wr_cycle[24470] = 1'b0;  addr_rom[24470]='h00003e58;  wr_data_rom[24470]='h00000000;
    rd_cycle[24471] = 1'b1;  wr_cycle[24471] = 1'b0;  addr_rom[24471]='h00003e5c;  wr_data_rom[24471]='h00000000;
    rd_cycle[24472] = 1'b1;  wr_cycle[24472] = 1'b0;  addr_rom[24472]='h00003e60;  wr_data_rom[24472]='h00000000;
    rd_cycle[24473] = 1'b1;  wr_cycle[24473] = 1'b0;  addr_rom[24473]='h00003e64;  wr_data_rom[24473]='h00000000;
    rd_cycle[24474] = 1'b1;  wr_cycle[24474] = 1'b0;  addr_rom[24474]='h00003e68;  wr_data_rom[24474]='h00000000;
    rd_cycle[24475] = 1'b1;  wr_cycle[24475] = 1'b0;  addr_rom[24475]='h00003e6c;  wr_data_rom[24475]='h00000000;
    rd_cycle[24476] = 1'b1;  wr_cycle[24476] = 1'b0;  addr_rom[24476]='h00003e70;  wr_data_rom[24476]='h00000000;
    rd_cycle[24477] = 1'b1;  wr_cycle[24477] = 1'b0;  addr_rom[24477]='h00003e74;  wr_data_rom[24477]='h00000000;
    rd_cycle[24478] = 1'b1;  wr_cycle[24478] = 1'b0;  addr_rom[24478]='h00003e78;  wr_data_rom[24478]='h00000000;
    rd_cycle[24479] = 1'b1;  wr_cycle[24479] = 1'b0;  addr_rom[24479]='h00003e7c;  wr_data_rom[24479]='h00000000;
    rd_cycle[24480] = 1'b1;  wr_cycle[24480] = 1'b0;  addr_rom[24480]='h00003e80;  wr_data_rom[24480]='h00000000;
    rd_cycle[24481] = 1'b1;  wr_cycle[24481] = 1'b0;  addr_rom[24481]='h00003e84;  wr_data_rom[24481]='h00000000;
    rd_cycle[24482] = 1'b1;  wr_cycle[24482] = 1'b0;  addr_rom[24482]='h00003e88;  wr_data_rom[24482]='h00000000;
    rd_cycle[24483] = 1'b1;  wr_cycle[24483] = 1'b0;  addr_rom[24483]='h00003e8c;  wr_data_rom[24483]='h00000000;
    rd_cycle[24484] = 1'b1;  wr_cycle[24484] = 1'b0;  addr_rom[24484]='h00003e90;  wr_data_rom[24484]='h00000000;
    rd_cycle[24485] = 1'b1;  wr_cycle[24485] = 1'b0;  addr_rom[24485]='h00003e94;  wr_data_rom[24485]='h00000000;
    rd_cycle[24486] = 1'b1;  wr_cycle[24486] = 1'b0;  addr_rom[24486]='h00003e98;  wr_data_rom[24486]='h00000000;
    rd_cycle[24487] = 1'b1;  wr_cycle[24487] = 1'b0;  addr_rom[24487]='h00003e9c;  wr_data_rom[24487]='h00000000;
    rd_cycle[24488] = 1'b1;  wr_cycle[24488] = 1'b0;  addr_rom[24488]='h00003ea0;  wr_data_rom[24488]='h00000000;
    rd_cycle[24489] = 1'b1;  wr_cycle[24489] = 1'b0;  addr_rom[24489]='h00003ea4;  wr_data_rom[24489]='h00000000;
    rd_cycle[24490] = 1'b1;  wr_cycle[24490] = 1'b0;  addr_rom[24490]='h00003ea8;  wr_data_rom[24490]='h00000000;
    rd_cycle[24491] = 1'b1;  wr_cycle[24491] = 1'b0;  addr_rom[24491]='h00003eac;  wr_data_rom[24491]='h00000000;
    rd_cycle[24492] = 1'b1;  wr_cycle[24492] = 1'b0;  addr_rom[24492]='h00003eb0;  wr_data_rom[24492]='h00000000;
    rd_cycle[24493] = 1'b1;  wr_cycle[24493] = 1'b0;  addr_rom[24493]='h00003eb4;  wr_data_rom[24493]='h00000000;
    rd_cycle[24494] = 1'b1;  wr_cycle[24494] = 1'b0;  addr_rom[24494]='h00003eb8;  wr_data_rom[24494]='h00000000;
    rd_cycle[24495] = 1'b1;  wr_cycle[24495] = 1'b0;  addr_rom[24495]='h00003ebc;  wr_data_rom[24495]='h00000000;
    rd_cycle[24496] = 1'b1;  wr_cycle[24496] = 1'b0;  addr_rom[24496]='h00003ec0;  wr_data_rom[24496]='h00000000;
    rd_cycle[24497] = 1'b1;  wr_cycle[24497] = 1'b0;  addr_rom[24497]='h00003ec4;  wr_data_rom[24497]='h00000000;
    rd_cycle[24498] = 1'b1;  wr_cycle[24498] = 1'b0;  addr_rom[24498]='h00003ec8;  wr_data_rom[24498]='h00000000;
    rd_cycle[24499] = 1'b1;  wr_cycle[24499] = 1'b0;  addr_rom[24499]='h00003ecc;  wr_data_rom[24499]='h00000000;
    rd_cycle[24500] = 1'b1;  wr_cycle[24500] = 1'b0;  addr_rom[24500]='h00003ed0;  wr_data_rom[24500]='h00000000;
    rd_cycle[24501] = 1'b1;  wr_cycle[24501] = 1'b0;  addr_rom[24501]='h00003ed4;  wr_data_rom[24501]='h00000000;
    rd_cycle[24502] = 1'b1;  wr_cycle[24502] = 1'b0;  addr_rom[24502]='h00003ed8;  wr_data_rom[24502]='h00000000;
    rd_cycle[24503] = 1'b1;  wr_cycle[24503] = 1'b0;  addr_rom[24503]='h00003edc;  wr_data_rom[24503]='h00000000;
    rd_cycle[24504] = 1'b1;  wr_cycle[24504] = 1'b0;  addr_rom[24504]='h00003ee0;  wr_data_rom[24504]='h00000000;
    rd_cycle[24505] = 1'b1;  wr_cycle[24505] = 1'b0;  addr_rom[24505]='h00003ee4;  wr_data_rom[24505]='h00000000;
    rd_cycle[24506] = 1'b1;  wr_cycle[24506] = 1'b0;  addr_rom[24506]='h00003ee8;  wr_data_rom[24506]='h00000000;
    rd_cycle[24507] = 1'b1;  wr_cycle[24507] = 1'b0;  addr_rom[24507]='h00003eec;  wr_data_rom[24507]='h00000000;
    rd_cycle[24508] = 1'b1;  wr_cycle[24508] = 1'b0;  addr_rom[24508]='h00003ef0;  wr_data_rom[24508]='h00000000;
    rd_cycle[24509] = 1'b1;  wr_cycle[24509] = 1'b0;  addr_rom[24509]='h00003ef4;  wr_data_rom[24509]='h00000000;
    rd_cycle[24510] = 1'b1;  wr_cycle[24510] = 1'b0;  addr_rom[24510]='h00003ef8;  wr_data_rom[24510]='h00000000;
    rd_cycle[24511] = 1'b1;  wr_cycle[24511] = 1'b0;  addr_rom[24511]='h00003efc;  wr_data_rom[24511]='h00000000;
    rd_cycle[24512] = 1'b1;  wr_cycle[24512] = 1'b0;  addr_rom[24512]='h00003f00;  wr_data_rom[24512]='h00000000;
    rd_cycle[24513] = 1'b1;  wr_cycle[24513] = 1'b0;  addr_rom[24513]='h00003f04;  wr_data_rom[24513]='h00000000;
    rd_cycle[24514] = 1'b1;  wr_cycle[24514] = 1'b0;  addr_rom[24514]='h00003f08;  wr_data_rom[24514]='h00000000;
    rd_cycle[24515] = 1'b1;  wr_cycle[24515] = 1'b0;  addr_rom[24515]='h00003f0c;  wr_data_rom[24515]='h00000000;
    rd_cycle[24516] = 1'b1;  wr_cycle[24516] = 1'b0;  addr_rom[24516]='h00003f10;  wr_data_rom[24516]='h00000000;
    rd_cycle[24517] = 1'b1;  wr_cycle[24517] = 1'b0;  addr_rom[24517]='h00003f14;  wr_data_rom[24517]='h00000000;
    rd_cycle[24518] = 1'b1;  wr_cycle[24518] = 1'b0;  addr_rom[24518]='h00003f18;  wr_data_rom[24518]='h00000000;
    rd_cycle[24519] = 1'b1;  wr_cycle[24519] = 1'b0;  addr_rom[24519]='h00003f1c;  wr_data_rom[24519]='h00000000;
    rd_cycle[24520] = 1'b1;  wr_cycle[24520] = 1'b0;  addr_rom[24520]='h00003f20;  wr_data_rom[24520]='h00000000;
    rd_cycle[24521] = 1'b1;  wr_cycle[24521] = 1'b0;  addr_rom[24521]='h00003f24;  wr_data_rom[24521]='h00000000;
    rd_cycle[24522] = 1'b1;  wr_cycle[24522] = 1'b0;  addr_rom[24522]='h00003f28;  wr_data_rom[24522]='h00000000;
    rd_cycle[24523] = 1'b1;  wr_cycle[24523] = 1'b0;  addr_rom[24523]='h00003f2c;  wr_data_rom[24523]='h00000000;
    rd_cycle[24524] = 1'b1;  wr_cycle[24524] = 1'b0;  addr_rom[24524]='h00003f30;  wr_data_rom[24524]='h00000000;
    rd_cycle[24525] = 1'b1;  wr_cycle[24525] = 1'b0;  addr_rom[24525]='h00003f34;  wr_data_rom[24525]='h00000000;
    rd_cycle[24526] = 1'b1;  wr_cycle[24526] = 1'b0;  addr_rom[24526]='h00003f38;  wr_data_rom[24526]='h00000000;
    rd_cycle[24527] = 1'b1;  wr_cycle[24527] = 1'b0;  addr_rom[24527]='h00003f3c;  wr_data_rom[24527]='h00000000;
    rd_cycle[24528] = 1'b1;  wr_cycle[24528] = 1'b0;  addr_rom[24528]='h00003f40;  wr_data_rom[24528]='h00000000;
    rd_cycle[24529] = 1'b1;  wr_cycle[24529] = 1'b0;  addr_rom[24529]='h00003f44;  wr_data_rom[24529]='h00000000;
    rd_cycle[24530] = 1'b1;  wr_cycle[24530] = 1'b0;  addr_rom[24530]='h00003f48;  wr_data_rom[24530]='h00000000;
    rd_cycle[24531] = 1'b1;  wr_cycle[24531] = 1'b0;  addr_rom[24531]='h00003f4c;  wr_data_rom[24531]='h00000000;
    rd_cycle[24532] = 1'b1;  wr_cycle[24532] = 1'b0;  addr_rom[24532]='h00003f50;  wr_data_rom[24532]='h00000000;
    rd_cycle[24533] = 1'b1;  wr_cycle[24533] = 1'b0;  addr_rom[24533]='h00003f54;  wr_data_rom[24533]='h00000000;
    rd_cycle[24534] = 1'b1;  wr_cycle[24534] = 1'b0;  addr_rom[24534]='h00003f58;  wr_data_rom[24534]='h00000000;
    rd_cycle[24535] = 1'b1;  wr_cycle[24535] = 1'b0;  addr_rom[24535]='h00003f5c;  wr_data_rom[24535]='h00000000;
    rd_cycle[24536] = 1'b1;  wr_cycle[24536] = 1'b0;  addr_rom[24536]='h00003f60;  wr_data_rom[24536]='h00000000;
    rd_cycle[24537] = 1'b1;  wr_cycle[24537] = 1'b0;  addr_rom[24537]='h00003f64;  wr_data_rom[24537]='h00000000;
    rd_cycle[24538] = 1'b1;  wr_cycle[24538] = 1'b0;  addr_rom[24538]='h00003f68;  wr_data_rom[24538]='h00000000;
    rd_cycle[24539] = 1'b1;  wr_cycle[24539] = 1'b0;  addr_rom[24539]='h00003f6c;  wr_data_rom[24539]='h00000000;
    rd_cycle[24540] = 1'b1;  wr_cycle[24540] = 1'b0;  addr_rom[24540]='h00003f70;  wr_data_rom[24540]='h00000000;
    rd_cycle[24541] = 1'b1;  wr_cycle[24541] = 1'b0;  addr_rom[24541]='h00003f74;  wr_data_rom[24541]='h00000000;
    rd_cycle[24542] = 1'b1;  wr_cycle[24542] = 1'b0;  addr_rom[24542]='h00003f78;  wr_data_rom[24542]='h00000000;
    rd_cycle[24543] = 1'b1;  wr_cycle[24543] = 1'b0;  addr_rom[24543]='h00003f7c;  wr_data_rom[24543]='h00000000;
    rd_cycle[24544] = 1'b1;  wr_cycle[24544] = 1'b0;  addr_rom[24544]='h00003f80;  wr_data_rom[24544]='h00000000;
    rd_cycle[24545] = 1'b1;  wr_cycle[24545] = 1'b0;  addr_rom[24545]='h00003f84;  wr_data_rom[24545]='h00000000;
    rd_cycle[24546] = 1'b1;  wr_cycle[24546] = 1'b0;  addr_rom[24546]='h00003f88;  wr_data_rom[24546]='h00000000;
    rd_cycle[24547] = 1'b1;  wr_cycle[24547] = 1'b0;  addr_rom[24547]='h00003f8c;  wr_data_rom[24547]='h00000000;
    rd_cycle[24548] = 1'b1;  wr_cycle[24548] = 1'b0;  addr_rom[24548]='h00003f90;  wr_data_rom[24548]='h00000000;
    rd_cycle[24549] = 1'b1;  wr_cycle[24549] = 1'b0;  addr_rom[24549]='h00003f94;  wr_data_rom[24549]='h00000000;
    rd_cycle[24550] = 1'b1;  wr_cycle[24550] = 1'b0;  addr_rom[24550]='h00003f98;  wr_data_rom[24550]='h00000000;
    rd_cycle[24551] = 1'b1;  wr_cycle[24551] = 1'b0;  addr_rom[24551]='h00003f9c;  wr_data_rom[24551]='h00000000;
    rd_cycle[24552] = 1'b1;  wr_cycle[24552] = 1'b0;  addr_rom[24552]='h00003fa0;  wr_data_rom[24552]='h00000000;
    rd_cycle[24553] = 1'b1;  wr_cycle[24553] = 1'b0;  addr_rom[24553]='h00003fa4;  wr_data_rom[24553]='h00000000;
    rd_cycle[24554] = 1'b1;  wr_cycle[24554] = 1'b0;  addr_rom[24554]='h00003fa8;  wr_data_rom[24554]='h00000000;
    rd_cycle[24555] = 1'b1;  wr_cycle[24555] = 1'b0;  addr_rom[24555]='h00003fac;  wr_data_rom[24555]='h00000000;
    rd_cycle[24556] = 1'b1;  wr_cycle[24556] = 1'b0;  addr_rom[24556]='h00003fb0;  wr_data_rom[24556]='h00000000;
    rd_cycle[24557] = 1'b1;  wr_cycle[24557] = 1'b0;  addr_rom[24557]='h00003fb4;  wr_data_rom[24557]='h00000000;
    rd_cycle[24558] = 1'b1;  wr_cycle[24558] = 1'b0;  addr_rom[24558]='h00003fb8;  wr_data_rom[24558]='h00000000;
    rd_cycle[24559] = 1'b1;  wr_cycle[24559] = 1'b0;  addr_rom[24559]='h00003fbc;  wr_data_rom[24559]='h00000000;
    rd_cycle[24560] = 1'b1;  wr_cycle[24560] = 1'b0;  addr_rom[24560]='h00003fc0;  wr_data_rom[24560]='h00000000;
    rd_cycle[24561] = 1'b1;  wr_cycle[24561] = 1'b0;  addr_rom[24561]='h00003fc4;  wr_data_rom[24561]='h00000000;
    rd_cycle[24562] = 1'b1;  wr_cycle[24562] = 1'b0;  addr_rom[24562]='h00003fc8;  wr_data_rom[24562]='h00000000;
    rd_cycle[24563] = 1'b1;  wr_cycle[24563] = 1'b0;  addr_rom[24563]='h00003fcc;  wr_data_rom[24563]='h00000000;
    rd_cycle[24564] = 1'b1;  wr_cycle[24564] = 1'b0;  addr_rom[24564]='h00003fd0;  wr_data_rom[24564]='h00000000;
    rd_cycle[24565] = 1'b1;  wr_cycle[24565] = 1'b0;  addr_rom[24565]='h00003fd4;  wr_data_rom[24565]='h00000000;
    rd_cycle[24566] = 1'b1;  wr_cycle[24566] = 1'b0;  addr_rom[24566]='h00003fd8;  wr_data_rom[24566]='h00000000;
    rd_cycle[24567] = 1'b1;  wr_cycle[24567] = 1'b0;  addr_rom[24567]='h00003fdc;  wr_data_rom[24567]='h00000000;
    rd_cycle[24568] = 1'b1;  wr_cycle[24568] = 1'b0;  addr_rom[24568]='h00003fe0;  wr_data_rom[24568]='h00000000;
    rd_cycle[24569] = 1'b1;  wr_cycle[24569] = 1'b0;  addr_rom[24569]='h00003fe4;  wr_data_rom[24569]='h00000000;
    rd_cycle[24570] = 1'b1;  wr_cycle[24570] = 1'b0;  addr_rom[24570]='h00003fe8;  wr_data_rom[24570]='h00000000;
    rd_cycle[24571] = 1'b1;  wr_cycle[24571] = 1'b0;  addr_rom[24571]='h00003fec;  wr_data_rom[24571]='h00000000;
    rd_cycle[24572] = 1'b1;  wr_cycle[24572] = 1'b0;  addr_rom[24572]='h00003ff0;  wr_data_rom[24572]='h00000000;
    rd_cycle[24573] = 1'b1;  wr_cycle[24573] = 1'b0;  addr_rom[24573]='h00003ff4;  wr_data_rom[24573]='h00000000;
    rd_cycle[24574] = 1'b1;  wr_cycle[24574] = 1'b0;  addr_rom[24574]='h00003ff8;  wr_data_rom[24574]='h00000000;
    rd_cycle[24575] = 1'b1;  wr_cycle[24575] = 1'b0;  addr_rom[24575]='h00003ffc;  wr_data_rom[24575]='h00000000;
end

initial begin
    validation_data[    0] = 'h00003530; 
    validation_data[    1] = 'h000026eb; 
    validation_data[    2] = 'h000020d5; 
    validation_data[    3] = 'h000033d8; 
    validation_data[    4] = 'h00002082; 
    validation_data[    5] = 'h00000fc1; 
    validation_data[    6] = 'h00003a24; 
    validation_data[    7] = 'h00000f46; 
    validation_data[    8] = 'h00001637; 
    validation_data[    9] = 'h000035da; 
    validation_data[   10] = 'h0000121c; 
    validation_data[   11] = 'h000016d9; 
    validation_data[   12] = 'h00001fc2; 
    validation_data[   13] = 'h00002bac; 
    validation_data[   14] = 'h00001aeb; 
    validation_data[   15] = 'h00002d7d; 
    validation_data[   16] = 'h00001b08; 
    validation_data[   17] = 'h00000251; 
    validation_data[   18] = 'h000029d8; 
    validation_data[   19] = 'h00002b1a; 
    validation_data[   20] = 'h00000e19; 
    validation_data[   21] = 'h00001bee; 
    validation_data[   22] = 'h000008d4; 
    validation_data[   23] = 'h00001274; 
    validation_data[   24] = 'h00002416; 
    validation_data[   25] = 'h00001678; 
    validation_data[   26] = 'h00001ae3; 
    validation_data[   27] = 'h000033e3; 
    validation_data[   28] = 'h00000bf0; 
    validation_data[   29] = 'h00001f8d; 
    validation_data[   30] = 'h000011ae; 
    validation_data[   31] = 'h00000f0a; 
    validation_data[   32] = 'h00001948; 
    validation_data[   33] = 'h00002cb6; 
    validation_data[   34] = 'h000031ff; 
    validation_data[   35] = 'h00000b89; 
    validation_data[   36] = 'h00002b8e; 
    validation_data[   37] = 'h00002797; 
    validation_data[   38] = 'h00002cfe; 
    validation_data[   39] = 'h00003090; 
    validation_data[   40] = 'h00001bef; 
    validation_data[   41] = 'h00003bf8; 
    validation_data[   42] = 'h00002c87; 
    validation_data[   43] = 'h00001328; 
    validation_data[   44] = 'h00003c78; 
    validation_data[   45] = 'h00000f5b; 
    validation_data[   46] = 'h00002c91; 
    validation_data[   47] = 'h000012c4; 
    validation_data[   48] = 'h00000ae1; 
    validation_data[   49] = 'h000019bc; 
    validation_data[   50] = 'h000013f3; 
    validation_data[   51] = 'h00001a35; 
    validation_data[   52] = 'h00000c13; 
    validation_data[   53] = 'h00001d2e; 
    validation_data[   54] = 'h00001525; 
    validation_data[   55] = 'h00000ee1; 
    validation_data[   56] = 'h0000137d; 
    validation_data[   57] = 'h00001caa; 
    validation_data[   58] = 'h00003374; 
    validation_data[   59] = 'h0000130e; 
    validation_data[   60] = 'h00000e8c; 
    validation_data[   61] = 'h0000026e; 
    validation_data[   62] = 'h00002be5; 
    validation_data[   63] = 'h00002e09; 
    validation_data[   64] = 'h00000ebf; 
    validation_data[   65] = 'h00003754; 
    validation_data[   66] = 'h00001680; 
    validation_data[   67] = 'h000020b4; 
    validation_data[   68] = 'h000013a6; 
    validation_data[   69] = 'h000029c8; 
    validation_data[   70] = 'h00002c53; 
    validation_data[   71] = 'h00000b56; 
    validation_data[   72] = 'h00002c2c; 
    validation_data[   73] = 'h000025f9; 
    validation_data[   74] = 'h0000352b; 
    validation_data[   75] = 'h000027a7; 
    validation_data[   76] = 'h000027a8; 
    validation_data[   77] = 'h0000293b; 
    validation_data[   78] = 'h00003652; 
    validation_data[   79] = 'h00001f3e; 
    validation_data[   80] = 'h00001772; 
    validation_data[   81] = 'h0000038b; 
    validation_data[   82] = 'h00003af2; 
    validation_data[   83] = 'h00003e3f; 
    validation_data[   84] = 'h00001ee2; 
    validation_data[   85] = 'h000039e6; 
    validation_data[   86] = 'h00003061; 
    validation_data[   87] = 'h00002026; 
    validation_data[   88] = 'h00001406; 
    validation_data[   89] = 'h0000233d; 
    validation_data[   90] = 'h00000c7a; 
    validation_data[   91] = 'h0000255f; 
    validation_data[   92] = 'h0000261c; 
    validation_data[   93] = 'h000023c8; 
    validation_data[   94] = 'h00002b66; 
    validation_data[   95] = 'h000010e9; 
    validation_data[   96] = 'h000019d9; 
    validation_data[   97] = 'h00000471; 
    validation_data[   98] = 'h00001176; 
    validation_data[   99] = 'h00000281; 
    validation_data[  100] = 'h00002fed; 
    validation_data[  101] = 'h000033cc; 
    validation_data[  102] = 'h00000cb2; 
    validation_data[  103] = 'h0000243b; 
    validation_data[  104] = 'h00001cc4; 
    validation_data[  105] = 'h00001d39; 
    validation_data[  106] = 'h00001f10; 
    validation_data[  107] = 'h00000ab8; 
    validation_data[  108] = 'h000009a6; 
    validation_data[  109] = 'h00001532; 
    validation_data[  110] = 'h0000365b; 
    validation_data[  111] = 'h00003932; 
    validation_data[  112] = 'h00000959; 
    validation_data[  113] = 'h00000706; 
    validation_data[  114] = 'h00002b4a; 
    validation_data[  115] = 'h000039f8; 
    validation_data[  116] = 'h00000cc4; 
    validation_data[  117] = 'h00002b50; 
    validation_data[  118] = 'h00001dcc; 
    validation_data[  119] = 'h000005fa; 
    validation_data[  120] = 'h00002131; 
    validation_data[  121] = 'h0000151e; 
    validation_data[  122] = 'h00000cf7; 
    validation_data[  123] = 'h00002ae7; 
    validation_data[  124] = 'h00001692; 
    validation_data[  125] = 'h0000155b; 
    validation_data[  126] = 'h000029da; 
    validation_data[  127] = 'h00003d50; 
    validation_data[  128] = 'h000032b2; 
    validation_data[  129] = 'h00002978; 
    validation_data[  130] = 'h00003359; 
    validation_data[  131] = 'h00002b52; 
    validation_data[  132] = 'h00000fa7; 
    validation_data[  133] = 'h00003c63; 
    validation_data[  134] = 'h00000386; 
    validation_data[  135] = 'h00002853; 
    validation_data[  136] = 'h000023f3; 
    validation_data[  137] = 'h00003540; 
    validation_data[  138] = 'h00001875; 
    validation_data[  139] = 'h000006af; 
    validation_data[  140] = 'h000004a0; 
    validation_data[  141] = 'h0000273b; 
    validation_data[  142] = 'h00003363; 
    validation_data[  143] = 'h00002fe7; 
    validation_data[  144] = 'h00002155; 
    validation_data[  145] = 'h0000221f; 
    validation_data[  146] = 'h00003691; 
    validation_data[  147] = 'h000000e3; 
    validation_data[  148] = 'h00002101; 
    validation_data[  149] = 'h00002e8e; 
    validation_data[  150] = 'h00002f83; 
    validation_data[  151] = 'h00003efa; 
    validation_data[  152] = 'h0000028b; 
    validation_data[  153] = 'h0000308c; 
    validation_data[  154] = 'h00003307; 
    validation_data[  155] = 'h00002e78; 
    validation_data[  156] = 'h0000327b; 
    validation_data[  157] = 'h0000344c; 
    validation_data[  158] = 'h00002bf2; 
    validation_data[  159] = 'h0000349e; 
    validation_data[  160] = 'h00002d8f; 
    validation_data[  161] = 'h00001485; 
    validation_data[  162] = 'h00001d81; 
    validation_data[  163] = 'h0000013d; 
    validation_data[  164] = 'h0000039d; 
    validation_data[  165] = 'h000007a7; 
    validation_data[  166] = 'h00003b4e; 
    validation_data[  167] = 'h00001e9c; 
    validation_data[  168] = 'h0000289c; 
    validation_data[  169] = 'h000006fd; 
    validation_data[  170] = 'h00003bb9; 
    validation_data[  171] = 'h000029e6; 
    validation_data[  172] = 'h000032be; 
    validation_data[  173] = 'h00003100; 
    validation_data[  174] = 'h00002d04; 
    validation_data[  175] = 'h00000c3f; 
    validation_data[  176] = 'h00001088; 
    validation_data[  177] = 'h00001df4; 
    validation_data[  178] = 'h0000221e; 
    validation_data[  179] = 'h000010cd; 
    validation_data[  180] = 'h00001bde; 
    validation_data[  181] = 'h00001353; 
    validation_data[  182] = 'h00002c4f; 
    validation_data[  183] = 'h0000343a; 
    validation_data[  184] = 'h00002a1f; 
    validation_data[  185] = 'h0000090f; 
    validation_data[  186] = 'h00000e4a; 
    validation_data[  187] = 'h00002bd1; 
    validation_data[  188] = 'h00000102; 
    validation_data[  189] = 'h00003603; 
    validation_data[  190] = 'h00000ce6; 
    validation_data[  191] = 'h000037ad; 
    validation_data[  192] = 'h00001bf5; 
    validation_data[  193] = 'h00000a18; 
    validation_data[  194] = 'h000001e5; 
    validation_data[  195] = 'h000002aa; 
    validation_data[  196] = 'h00002a9d; 
    validation_data[  197] = 'h000013b5; 
    validation_data[  198] = 'h00000ee9; 
    validation_data[  199] = 'h0000252d; 
    validation_data[  200] = 'h00003419; 
    validation_data[  201] = 'h00003341; 
    validation_data[  202] = 'h00001dc4; 
    validation_data[  203] = 'h00000a0a; 
    validation_data[  204] = 'h0000373b; 
    validation_data[  205] = 'h00000a4c; 
    validation_data[  206] = 'h000010d4; 
    validation_data[  207] = 'h00002d5d; 
    validation_data[  208] = 'h0000168d; 
    validation_data[  209] = 'h000014f2; 
    validation_data[  210] = 'h0000342d; 
    validation_data[  211] = 'h00003b29; 
    validation_data[  212] = 'h000023c6; 
    validation_data[  213] = 'h00000933; 
    validation_data[  214] = 'h000007fd; 
    validation_data[  215] = 'h0000068d; 
    validation_data[  216] = 'h0000141e; 
    validation_data[  217] = 'h00000624; 
    validation_data[  218] = 'h000028e9; 
    validation_data[  219] = 'h0000024a; 
    validation_data[  220] = 'h00000855; 
    validation_data[  221] = 'h00000d0c; 
    validation_data[  222] = 'h0000002f; 
    validation_data[  223] = 'h000030fc; 
    validation_data[  224] = 'h00000640; 
    validation_data[  225] = 'h00000188; 
    validation_data[  226] = 'h00001bed; 
    validation_data[  227] = 'h00001d15; 
    validation_data[  228] = 'h00002c89; 
    validation_data[  229] = 'h00002dda; 
    validation_data[  230] = 'h000014a4; 
    validation_data[  231] = 'h000025c9; 
    validation_data[  232] = 'h00002b86; 
    validation_data[  233] = 'h00003e1d; 
    validation_data[  234] = 'h00001fe3; 
    validation_data[  235] = 'h000016e5; 
    validation_data[  236] = 'h00001689; 
    validation_data[  237] = 'h000016fb; 
    validation_data[  238] = 'h00002b45; 
    validation_data[  239] = 'h00003033; 
    validation_data[  240] = 'h00001406; 
    validation_data[  241] = 'h0000396b; 
    validation_data[  242] = 'h0000183c; 
    validation_data[  243] = 'h00001500; 
    validation_data[  244] = 'h0000322e; 
    validation_data[  245] = 'h00000ac8; 
    validation_data[  246] = 'h0000056a; 
    validation_data[  247] = 'h00000b69; 
    validation_data[  248] = 'h00003703; 
    validation_data[  249] = 'h0000259f; 
    validation_data[  250] = 'h0000083a; 
    validation_data[  251] = 'h00001025; 
    validation_data[  252] = 'h00001612; 
    validation_data[  253] = 'h00002a7e; 
    validation_data[  254] = 'h000038a0; 
    validation_data[  255] = 'h000036d9; 
    validation_data[  256] = 'h00000540; 
    validation_data[  257] = 'h00001b94; 
    validation_data[  258] = 'h00000ce5; 
    validation_data[  259] = 'h0000171a; 
    validation_data[  260] = 'h00000b0c; 
    validation_data[  261] = 'h00002e1a; 
    validation_data[  262] = 'h00000d1e; 
    validation_data[  263] = 'h00003cbe; 
    validation_data[  264] = 'h00003f5d; 
    validation_data[  265] = 'h00000b88; 
    validation_data[  266] = 'h00000a48; 
    validation_data[  267] = 'h00002afb; 
    validation_data[  268] = 'h00001ac4; 
    validation_data[  269] = 'h00003378; 
    validation_data[  270] = 'h00000e9b; 
    validation_data[  271] = 'h00003553; 
    validation_data[  272] = 'h000021c4; 
    validation_data[  273] = 'h000023b8; 
    validation_data[  274] = 'h00002dda; 
    validation_data[  275] = 'h00001bc2; 
    validation_data[  276] = 'h00002ce5; 
    validation_data[  277] = 'h00001929; 
    validation_data[  278] = 'h000010b4; 
    validation_data[  279] = 'h00002654; 
    validation_data[  280] = 'h000004d1; 
    validation_data[  281] = 'h0000275d; 
    validation_data[  282] = 'h00000858; 
    validation_data[  283] = 'h0000352f; 
    validation_data[  284] = 'h0000090f; 
    validation_data[  285] = 'h00000ed4; 
    validation_data[  286] = 'h00000eb7; 
    validation_data[  287] = 'h00000752; 
    validation_data[  288] = 'h000008ae; 
    validation_data[  289] = 'h00001f18; 
    validation_data[  290] = 'h00002a6e; 
    validation_data[  291] = 'h00001f64; 
    validation_data[  292] = 'h00003020; 
    validation_data[  293] = 'h00003dd0; 
    validation_data[  294] = 'h00000cbe; 
    validation_data[  295] = 'h000009d6; 
    validation_data[  296] = 'h0000112d; 
    validation_data[  297] = 'h00002a6c; 
    validation_data[  298] = 'h000019bf; 
    validation_data[  299] = 'h000016f8; 
    validation_data[  300] = 'h00002d1e; 
    validation_data[  301] = 'h00003b56; 
    validation_data[  302] = 'h00001da9; 
    validation_data[  303] = 'h00003fe7; 
    validation_data[  304] = 'h000034f8; 
    validation_data[  305] = 'h00000cea; 
    validation_data[  306] = 'h00001a9b; 
    validation_data[  307] = 'h00002191; 
    validation_data[  308] = 'h00003f92; 
    validation_data[  309] = 'h000003c3; 
    validation_data[  310] = 'h00003174; 
    validation_data[  311] = 'h00002e86; 
    validation_data[  312] = 'h00003eaf; 
    validation_data[  313] = 'h00001ca4; 
    validation_data[  314] = 'h00003c39; 
    validation_data[  315] = 'h00002bcd; 
    validation_data[  316] = 'h00001fc8; 
    validation_data[  317] = 'h00002f3b; 
    validation_data[  318] = 'h000010f4; 
    validation_data[  319] = 'h00001e0e; 
    validation_data[  320] = 'h00001ebc; 
    validation_data[  321] = 'h000024d7; 
    validation_data[  322] = 'h0000160b; 
    validation_data[  323] = 'h00000f98; 
    validation_data[  324] = 'h000020fe; 
    validation_data[  325] = 'h000021d0; 
    validation_data[  326] = 'h00003978; 
    validation_data[  327] = 'h00001bdc; 
    validation_data[  328] = 'h00001053; 
    validation_data[  329] = 'h00002109; 
    validation_data[  330] = 'h00003e49; 
    validation_data[  331] = 'h000018dc; 
    validation_data[  332] = 'h00000aee; 
    validation_data[  333] = 'h000006ae; 
    validation_data[  334] = 'h0000223d; 
    validation_data[  335] = 'h00000a7c; 
    validation_data[  336] = 'h0000288e; 
    validation_data[  337] = 'h0000195b; 
    validation_data[  338] = 'h00002366; 
    validation_data[  339] = 'h000021cc; 
    validation_data[  340] = 'h00000dfa; 
    validation_data[  341] = 'h000015ea; 
    validation_data[  342] = 'h00002c7f; 
    validation_data[  343] = 'h00000dac; 
    validation_data[  344] = 'h00002c7a; 
    validation_data[  345] = 'h0000257e; 
    validation_data[  346] = 'h0000059f; 
    validation_data[  347] = 'h00002ec7; 
    validation_data[  348] = 'h000015a0; 
    validation_data[  349] = 'h00000182; 
    validation_data[  350] = 'h00003bf0; 
    validation_data[  351] = 'h0000166a; 
    validation_data[  352] = 'h00001aa8; 
    validation_data[  353] = 'h00000931; 
    validation_data[  354] = 'h00001095; 
    validation_data[  355] = 'h00002000; 
    validation_data[  356] = 'h00000e18; 
    validation_data[  357] = 'h00001911; 
    validation_data[  358] = 'h000033e4; 
    validation_data[  359] = 'h000021eb; 
    validation_data[  360] = 'h00000b8f; 
    validation_data[  361] = 'h00001ec2; 
    validation_data[  362] = 'h000024b7; 
    validation_data[  363] = 'h000032c5; 
    validation_data[  364] = 'h00000c63; 
    validation_data[  365] = 'h00002301; 
    validation_data[  366] = 'h000011d3; 
    validation_data[  367] = 'h00000917; 
    validation_data[  368] = 'h0000365c; 
    validation_data[  369] = 'h0000259d; 
    validation_data[  370] = 'h00000e21; 
    validation_data[  371] = 'h0000311c; 
    validation_data[  372] = 'h000013ca; 
    validation_data[  373] = 'h00001a83; 
    validation_data[  374] = 'h00000203; 
    validation_data[  375] = 'h00002c4b; 
    validation_data[  376] = 'h00003ff8; 
    validation_data[  377] = 'h00001efa; 
    validation_data[  378] = 'h00000e76; 
    validation_data[  379] = 'h00000276; 
    validation_data[  380] = 'h00001bc2; 
    validation_data[  381] = 'h00001026; 
    validation_data[  382] = 'h00001785; 
    validation_data[  383] = 'h00003750; 
    validation_data[  384] = 'h00001c64; 
    validation_data[  385] = 'h0000177d; 
    validation_data[  386] = 'h00003b94; 
    validation_data[  387] = 'h000014bf; 
    validation_data[  388] = 'h00003ff3; 
    validation_data[  389] = 'h00002d4d; 
    validation_data[  390] = 'h0000216f; 
    validation_data[  391] = 'h00003266; 
    validation_data[  392] = 'h00002413; 
    validation_data[  393] = 'h00002588; 
    validation_data[  394] = 'h0000180e; 
    validation_data[  395] = 'h00000470; 
    validation_data[  396] = 'h00000eda; 
    validation_data[  397] = 'h00000211; 
    validation_data[  398] = 'h0000219f; 
    validation_data[  399] = 'h00001deb; 
    validation_data[  400] = 'h00002149; 
    validation_data[  401] = 'h000037fb; 
    validation_data[  402] = 'h00001705; 
    validation_data[  403] = 'h00002a82; 
    validation_data[  404] = 'h00001574; 
    validation_data[  405] = 'h00002fc4; 
    validation_data[  406] = 'h00002977; 
    validation_data[  407] = 'h0000241c; 
    validation_data[  408] = 'h00000d6c; 
    validation_data[  409] = 'h00001673; 
    validation_data[  410] = 'h000024eb; 
    validation_data[  411] = 'h000009af; 
    validation_data[  412] = 'h00000ea1; 
    validation_data[  413] = 'h000025e7; 
    validation_data[  414] = 'h00000735; 
    validation_data[  415] = 'h0000179b; 
    validation_data[  416] = 'h000003f4; 
    validation_data[  417] = 'h00002fbd; 
    validation_data[  418] = 'h00001656; 
    validation_data[  419] = 'h00001041; 
    validation_data[  420] = 'h000036f3; 
    validation_data[  421] = 'h0000242b; 
    validation_data[  422] = 'h00000631; 
    validation_data[  423] = 'h00003257; 
    validation_data[  424] = 'h00000521; 
    validation_data[  425] = 'h0000010a; 
    validation_data[  426] = 'h000009df; 
    validation_data[  427] = 'h00001269; 
    validation_data[  428] = 'h00001add; 
    validation_data[  429] = 'h00000028; 
    validation_data[  430] = 'h0000137c; 
    validation_data[  431] = 'h00000e01; 
    validation_data[  432] = 'h0000280b; 
    validation_data[  433] = 'h00003986; 
    validation_data[  434] = 'h00003e80; 
    validation_data[  435] = 'h000033c8; 
    validation_data[  436] = 'h00003166; 
    validation_data[  437] = 'h00000510; 
    validation_data[  438] = 'h00001f1f; 
    validation_data[  439] = 'h00001946; 
    validation_data[  440] = 'h0000137e; 
    validation_data[  441] = 'h00003895; 
    validation_data[  442] = 'h000030d7; 
    validation_data[  443] = 'h000010a3; 
    validation_data[  444] = 'h00002d73; 
    validation_data[  445] = 'h00002a9e; 
    validation_data[  446] = 'h00000c99; 
    validation_data[  447] = 'h00000487; 
    validation_data[  448] = 'h00000529; 
    validation_data[  449] = 'h00003ef8; 
    validation_data[  450] = 'h00000b82; 
    validation_data[  451] = 'h000008a3; 
    validation_data[  452] = 'h00000fa8; 
    validation_data[  453] = 'h00001846; 
    validation_data[  454] = 'h000007ca; 
    validation_data[  455] = 'h00000b0f; 
    validation_data[  456] = 'h00002a1d; 
    validation_data[  457] = 'h00001d15; 
    validation_data[  458] = 'h000037cd; 
    validation_data[  459] = 'h00002288; 
    validation_data[  460] = 'h00000a54; 
    validation_data[  461] = 'h00002009; 
    validation_data[  462] = 'h00000cf5; 
    validation_data[  463] = 'h0000227d; 
    validation_data[  464] = 'h000028a4; 
    validation_data[  465] = 'h00000291; 
    validation_data[  466] = 'h00003a89; 
    validation_data[  467] = 'h00003734; 
    validation_data[  468] = 'h00001ae0; 
    validation_data[  469] = 'h00002766; 
    validation_data[  470] = 'h00000a7f; 
    validation_data[  471] = 'h000036df; 
    validation_data[  472] = 'h00001c44; 
    validation_data[  473] = 'h00002aed; 
    validation_data[  474] = 'h00001de4; 
    validation_data[  475] = 'h000038bb; 
    validation_data[  476] = 'h00003493; 
    validation_data[  477] = 'h00002c8d; 
    validation_data[  478] = 'h00001597; 
    validation_data[  479] = 'h00003622; 
    validation_data[  480] = 'h00003323; 
    validation_data[  481] = 'h000003a7; 
    validation_data[  482] = 'h00002e30; 
    validation_data[  483] = 'h00002512; 
    validation_data[  484] = 'h00000316; 
    validation_data[  485] = 'h000009d9; 
    validation_data[  486] = 'h00002b52; 
    validation_data[  487] = 'h00003b4c; 
    validation_data[  488] = 'h00002db5; 
    validation_data[  489] = 'h00000567; 
    validation_data[  490] = 'h000017b3; 
    validation_data[  491] = 'h000008f3; 
    validation_data[  492] = 'h000031b1; 
    validation_data[  493] = 'h000016b0; 
    validation_data[  494] = 'h00002439; 
    validation_data[  495] = 'h000010b7; 
    validation_data[  496] = 'h00001834; 
    validation_data[  497] = 'h00002917; 
    validation_data[  498] = 'h000029c8; 
    validation_data[  499] = 'h00002705; 
    validation_data[  500] = 'h000030b4; 
    validation_data[  501] = 'h00003050; 
    validation_data[  502] = 'h00003920; 
    validation_data[  503] = 'h00003b15; 
    validation_data[  504] = 'h000033f7; 
    validation_data[  505] = 'h000025e3; 
    validation_data[  506] = 'h00001e01; 
    validation_data[  507] = 'h00003612; 
    validation_data[  508] = 'h00002de4; 
    validation_data[  509] = 'h00002faf; 
    validation_data[  510] = 'h00002a73; 
    validation_data[  511] = 'h00003599; 
    validation_data[  512] = 'h0000335f; 
    validation_data[  513] = 'h000011b4; 
    validation_data[  514] = 'h00003b58; 
    validation_data[  515] = 'h000032f8; 
    validation_data[  516] = 'h00003596; 
    validation_data[  517] = 'h00002dce; 
    validation_data[  518] = 'h000033a2; 
    validation_data[  519] = 'h00000d6c; 
    validation_data[  520] = 'h000021ae; 
    validation_data[  521] = 'h0000190e; 
    validation_data[  522] = 'h00000c2d; 
    validation_data[  523] = 'h00001d2d; 
    validation_data[  524] = 'h00001842; 
    validation_data[  525] = 'h00000fb5; 
    validation_data[  526] = 'h00002b8d; 
    validation_data[  527] = 'h000008a1; 
    validation_data[  528] = 'h0000298b; 
    validation_data[  529] = 'h00001202; 
    validation_data[  530] = 'h00003f31; 
    validation_data[  531] = 'h000013c5; 
    validation_data[  532] = 'h00002336; 
    validation_data[  533] = 'h00002b99; 
    validation_data[  534] = 'h00001623; 
    validation_data[  535] = 'h000035e0; 
    validation_data[  536] = 'h00003493; 
    validation_data[  537] = 'h000000bb; 
    validation_data[  538] = 'h00002958; 
    validation_data[  539] = 'h00002baf; 
    validation_data[  540] = 'h00002063; 
    validation_data[  541] = 'h0000209c; 
    validation_data[  542] = 'h00000761; 
    validation_data[  543] = 'h00002b28; 
    validation_data[  544] = 'h000022fa; 
    validation_data[  545] = 'h00001100; 
    validation_data[  546] = 'h000029d0; 
    validation_data[  547] = 'h00000d30; 
    validation_data[  548] = 'h00002170; 
    validation_data[  549] = 'h000001bf; 
    validation_data[  550] = 'h00000db1; 
    validation_data[  551] = 'h00000f09; 
    validation_data[  552] = 'h0000204f; 
    validation_data[  553] = 'h0000328d; 
    validation_data[  554] = 'h00003ba5; 
    validation_data[  555] = 'h0000275a; 
    validation_data[  556] = 'h00003126; 
    validation_data[  557] = 'h00000613; 
    validation_data[  558] = 'h000024ab; 
    validation_data[  559] = 'h00000ba9; 
    validation_data[  560] = 'h00001f2f; 
    validation_data[  561] = 'h00001d1f; 
    validation_data[  562] = 'h00003333; 
    validation_data[  563] = 'h00002807; 
    validation_data[  564] = 'h000033f5; 
    validation_data[  565] = 'h000019eb; 
    validation_data[  566] = 'h00002855; 
    validation_data[  567] = 'h0000053f; 
    validation_data[  568] = 'h000032d4; 
    validation_data[  569] = 'h00000a4d; 
    validation_data[  570] = 'h00002d83; 
    validation_data[  571] = 'h000026e6; 
    validation_data[  572] = 'h00000236; 
    validation_data[  573] = 'h00000b50; 
    validation_data[  574] = 'h0000119f; 
    validation_data[  575] = 'h000036ec; 
    validation_data[  576] = 'h000019ed; 
    validation_data[  577] = 'h0000145b; 
    validation_data[  578] = 'h00003527; 
    validation_data[  579] = 'h00003452; 
    validation_data[  580] = 'h00000da9; 
    validation_data[  581] = 'h00003f8b; 
    validation_data[  582] = 'h00002533; 
    validation_data[  583] = 'h000008e2; 
    validation_data[  584] = 'h00002689; 
    validation_data[  585] = 'h000027d1; 
    validation_data[  586] = 'h00003f08; 
    validation_data[  587] = 'h00002a28; 
    validation_data[  588] = 'h00003baa; 
    validation_data[  589] = 'h0000260f; 
    validation_data[  590] = 'h000002f5; 
    validation_data[  591] = 'h00001a5b; 
    validation_data[  592] = 'h0000072c; 
    validation_data[  593] = 'h00003bc2; 
    validation_data[  594] = 'h00001b63; 
    validation_data[  595] = 'h00003bd1; 
    validation_data[  596] = 'h00003415; 
    validation_data[  597] = 'h000024b0; 
    validation_data[  598] = 'h0000077d; 
    validation_data[  599] = 'h00001593; 
    validation_data[  600] = 'h00002b62; 
    validation_data[  601] = 'h000037d5; 
    validation_data[  602] = 'h00003753; 
    validation_data[  603] = 'h00000b08; 
    validation_data[  604] = 'h00003617; 
    validation_data[  605] = 'h00003d64; 
    validation_data[  606] = 'h000007b4; 
    validation_data[  607] = 'h0000260a; 
    validation_data[  608] = 'h0000000d; 
    validation_data[  609] = 'h00002db5; 
    validation_data[  610] = 'h00003c86; 
    validation_data[  611] = 'h0000392a; 
    validation_data[  612] = 'h00003cbc; 
    validation_data[  613] = 'h00003161; 
    validation_data[  614] = 'h00003be1; 
    validation_data[  615] = 'h00002cb9; 
    validation_data[  616] = 'h00000706; 
    validation_data[  617] = 'h000027de; 
    validation_data[  618] = 'h0000319a; 
    validation_data[  619] = 'h000027a1; 
    validation_data[  620] = 'h00002f21; 
    validation_data[  621] = 'h0000070a; 
    validation_data[  622] = 'h00000a3e; 
    validation_data[  623] = 'h00001e6e; 
    validation_data[  624] = 'h00002cd4; 
    validation_data[  625] = 'h00000d1c; 
    validation_data[  626] = 'h00001544; 
    validation_data[  627] = 'h0000218e; 
    validation_data[  628] = 'h00000299; 
    validation_data[  629] = 'h00001eaf; 
    validation_data[  630] = 'h00000b8d; 
    validation_data[  631] = 'h00000264; 
    validation_data[  632] = 'h00000f17; 
    validation_data[  633] = 'h000027ea; 
    validation_data[  634] = 'h00002cfe; 
    validation_data[  635] = 'h000002d9; 
    validation_data[  636] = 'h00000d4e; 
    validation_data[  637] = 'h00002e54; 
    validation_data[  638] = 'h00000ff8; 
    validation_data[  639] = 'h000001fe; 
    validation_data[  640] = 'h0000069a; 
    validation_data[  641] = 'h00001f23; 
    validation_data[  642] = 'h000007b9; 
    validation_data[  643] = 'h00003a32; 
    validation_data[  644] = 'h00000682; 
    validation_data[  645] = 'h00000f0c; 
    validation_data[  646] = 'h000001eb; 
    validation_data[  647] = 'h00001f58; 
    validation_data[  648] = 'h00002d31; 
    validation_data[  649] = 'h00001cee; 
    validation_data[  650] = 'h00003a3c; 
    validation_data[  651] = 'h00002124; 
    validation_data[  652] = 'h000029c7; 
    validation_data[  653] = 'h0000151a; 
    validation_data[  654] = 'h000022b0; 
    validation_data[  655] = 'h000039b4; 
    validation_data[  656] = 'h0000310c; 
    validation_data[  657] = 'h00001694; 
    validation_data[  658] = 'h00000b25; 
    validation_data[  659] = 'h000027eb; 
    validation_data[  660] = 'h000001ed; 
    validation_data[  661] = 'h000032fc; 
    validation_data[  662] = 'h000035c0; 
    validation_data[  663] = 'h000037c7; 
    validation_data[  664] = 'h00001a33; 
    validation_data[  665] = 'h0000122e; 
    validation_data[  666] = 'h00000942; 
    validation_data[  667] = 'h00000645; 
    validation_data[  668] = 'h00001030; 
    validation_data[  669] = 'h000035e1; 
    validation_data[  670] = 'h00001895; 
    validation_data[  671] = 'h00003fb6; 
    validation_data[  672] = 'h00002d1b; 
    validation_data[  673] = 'h0000193c; 
    validation_data[  674] = 'h00000d98; 
    validation_data[  675] = 'h0000031f; 
    validation_data[  676] = 'h000017f6; 
    validation_data[  677] = 'h00000cdd; 
    validation_data[  678] = 'h00001730; 
    validation_data[  679] = 'h000006b2; 
    validation_data[  680] = 'h00003382; 
    validation_data[  681] = 'h00000eca; 
    validation_data[  682] = 'h0000316b; 
    validation_data[  683] = 'h00003e94; 
    validation_data[  684] = 'h00001957; 
    validation_data[  685] = 'h00002561; 
    validation_data[  686] = 'h00003494; 
    validation_data[  687] = 'h00003e4b; 
    validation_data[  688] = 'h00000367; 
    validation_data[  689] = 'h0000292b; 
    validation_data[  690] = 'h00001899; 
    validation_data[  691] = 'h0000189d; 
    validation_data[  692] = 'h000035d4; 
    validation_data[  693] = 'h000025c2; 
    validation_data[  694] = 'h00002c71; 
    validation_data[  695] = 'h0000257e; 
    validation_data[  696] = 'h00001501; 
    validation_data[  697] = 'h0000187d; 
    validation_data[  698] = 'h00001690; 
    validation_data[  699] = 'h0000181c; 
    validation_data[  700] = 'h00001841; 
    validation_data[  701] = 'h00002765; 
    validation_data[  702] = 'h0000094f; 
    validation_data[  703] = 'h00001a39; 
    validation_data[  704] = 'h00002673; 
    validation_data[  705] = 'h00003ebf; 
    validation_data[  706] = 'h000010a1; 
    validation_data[  707] = 'h000030e2; 
    validation_data[  708] = 'h0000316f; 
    validation_data[  709] = 'h0000364c; 
    validation_data[  710] = 'h000010af; 
    validation_data[  711] = 'h00001598; 
    validation_data[  712] = 'h000006c7; 
    validation_data[  713] = 'h00003781; 
    validation_data[  714] = 'h00000bfa; 
    validation_data[  715] = 'h00002a6e; 
    validation_data[  716] = 'h00002c6c; 
    validation_data[  717] = 'h000011fe; 
    validation_data[  718] = 'h00003861; 
    validation_data[  719] = 'h00003868; 
    validation_data[  720] = 'h00002cb3; 
    validation_data[  721] = 'h00002314; 
    validation_data[  722] = 'h00003977; 
    validation_data[  723] = 'h00000a0d; 
    validation_data[  724] = 'h00000ea3; 
    validation_data[  725] = 'h00002c3b; 
    validation_data[  726] = 'h00001aa5; 
    validation_data[  727] = 'h000003dc; 
    validation_data[  728] = 'h000009b0; 
    validation_data[  729] = 'h00000a4f; 
    validation_data[  730] = 'h0000306c; 
    validation_data[  731] = 'h00000097; 
    validation_data[  732] = 'h0000104a; 
    validation_data[  733] = 'h00000e53; 
    validation_data[  734] = 'h000012e3; 
    validation_data[  735] = 'h00003c1c; 
    validation_data[  736] = 'h000011cd; 
    validation_data[  737] = 'h0000169d; 
    validation_data[  738] = 'h00002a5e; 
    validation_data[  739] = 'h000037e4; 
    validation_data[  740] = 'h00001f69; 
    validation_data[  741] = 'h000024ff; 
    validation_data[  742] = 'h00000355; 
    validation_data[  743] = 'h00000e68; 
    validation_data[  744] = 'h0000146c; 
    validation_data[  745] = 'h00002ca7; 
    validation_data[  746] = 'h0000273c; 
    validation_data[  747] = 'h00002ca4; 
    validation_data[  748] = 'h00002b21; 
    validation_data[  749] = 'h00003b85; 
    validation_data[  750] = 'h00002c6d; 
    validation_data[  751] = 'h00002241; 
    validation_data[  752] = 'h000020c2; 
    validation_data[  753] = 'h0000179c; 
    validation_data[  754] = 'h000009f4; 
    validation_data[  755] = 'h00002ec7; 
    validation_data[  756] = 'h000037a1; 
    validation_data[  757] = 'h00002223; 
    validation_data[  758] = 'h000038de; 
    validation_data[  759] = 'h00000c9b; 
    validation_data[  760] = 'h00003b3c; 
    validation_data[  761] = 'h00002c16; 
    validation_data[  762] = 'h00003e5b; 
    validation_data[  763] = 'h00002a1b; 
    validation_data[  764] = 'h00003ed0; 
    validation_data[  765] = 'h00001764; 
    validation_data[  766] = 'h000028e4; 
    validation_data[  767] = 'h0000055e; 
    validation_data[  768] = 'h00003db4; 
    validation_data[  769] = 'h00001540; 
    validation_data[  770] = 'h0000173d; 
    validation_data[  771] = 'h000010b6; 
    validation_data[  772] = 'h00000b46; 
    validation_data[  773] = 'h0000232a; 
    validation_data[  774] = 'h0000117e; 
    validation_data[  775] = 'h00002649; 
    validation_data[  776] = 'h0000035a; 
    validation_data[  777] = 'h00001ae3; 
    validation_data[  778] = 'h0000071c; 
    validation_data[  779] = 'h000014cf; 
    validation_data[  780] = 'h00000c6d; 
    validation_data[  781] = 'h00000795; 
    validation_data[  782] = 'h000014d9; 
    validation_data[  783] = 'h00002956; 
    validation_data[  784] = 'h000013f2; 
    validation_data[  785] = 'h00001bd4; 
    validation_data[  786] = 'h000030e3; 
    validation_data[  787] = 'h000003e9; 
    validation_data[  788] = 'h00003af7; 
    validation_data[  789] = 'h000017cb; 
    validation_data[  790] = 'h0000114e; 
    validation_data[  791] = 'h00002b32; 
    validation_data[  792] = 'h00002daa; 
    validation_data[  793] = 'h00003712; 
    validation_data[  794] = 'h0000279a; 
    validation_data[  795] = 'h00000bc2; 
    validation_data[  796] = 'h0000253b; 
    validation_data[  797] = 'h00001a13; 
    validation_data[  798] = 'h00002a7b; 
    validation_data[  799] = 'h00003b83; 
    validation_data[  800] = 'h00001808; 
    validation_data[  801] = 'h00001acc; 
    validation_data[  802] = 'h00003767; 
    validation_data[  803] = 'h000012d7; 
    validation_data[  804] = 'h00000402; 
    validation_data[  805] = 'h00002880; 
    validation_data[  806] = 'h00003345; 
    validation_data[  807] = 'h0000003a; 
    validation_data[  808] = 'h00003833; 
    validation_data[  809] = 'h0000371b; 
    validation_data[  810] = 'h00001149; 
    validation_data[  811] = 'h000032e5; 
    validation_data[  812] = 'h0000385f; 
    validation_data[  813] = 'h00003c28; 
    validation_data[  814] = 'h0000269a; 
    validation_data[  815] = 'h00001524; 
    validation_data[  816] = 'h0000209b; 
    validation_data[  817] = 'h00002944; 
    validation_data[  818] = 'h00002370; 
    validation_data[  819] = 'h00001bc3; 
    validation_data[  820] = 'h00003677; 
    validation_data[  821] = 'h00003da4; 
    validation_data[  822] = 'h00001f2a; 
    validation_data[  823] = 'h00000f10; 
    validation_data[  824] = 'h000026c4; 
    validation_data[  825] = 'h00003ff8; 
    validation_data[  826] = 'h00001410; 
    validation_data[  827] = 'h00000acd; 
    validation_data[  828] = 'h000031a9; 
    validation_data[  829] = 'h000014a7; 
    validation_data[  830] = 'h0000235b; 
    validation_data[  831] = 'h000004a0; 
    validation_data[  832] = 'h0000232a; 
    validation_data[  833] = 'h00000d96; 
    validation_data[  834] = 'h00000cbc; 
    validation_data[  835] = 'h00000ec1; 
    validation_data[  836] = 'h00003fb3; 
    validation_data[  837] = 'h000004cf; 
    validation_data[  838] = 'h00001d8a; 
    validation_data[  839] = 'h00002e6c; 
    validation_data[  840] = 'h00003cdb; 
    validation_data[  841] = 'h00001fb4; 
    validation_data[  842] = 'h0000344b; 
    validation_data[  843] = 'h000008f8; 
    validation_data[  844] = 'h0000245b; 
    validation_data[  845] = 'h0000234a; 
    validation_data[  846] = 'h00002846; 
    validation_data[  847] = 'h00003cf8; 
    validation_data[  848] = 'h0000389a; 
    validation_data[  849] = 'h0000248d; 
    validation_data[  850] = 'h00002e24; 
    validation_data[  851] = 'h00000a3b; 
    validation_data[  852] = 'h000003e3; 
    validation_data[  853] = 'h000000ab; 
    validation_data[  854] = 'h000035f1; 
    validation_data[  855] = 'h000032e7; 
    validation_data[  856] = 'h0000201e; 
    validation_data[  857] = 'h00001a00; 
    validation_data[  858] = 'h00000971; 
    validation_data[  859] = 'h0000209c; 
    validation_data[  860] = 'h0000109a; 
    validation_data[  861] = 'h00002862; 
    validation_data[  862] = 'h000027e6; 
    validation_data[  863] = 'h00002a6b; 
    validation_data[  864] = 'h000000f1; 
    validation_data[  865] = 'h00003992; 
    validation_data[  866] = 'h00002139; 
    validation_data[  867] = 'h00002ac8; 
    validation_data[  868] = 'h000012a7; 
    validation_data[  869] = 'h00003014; 
    validation_data[  870] = 'h00003995; 
    validation_data[  871] = 'h00002468; 
    validation_data[  872] = 'h000026ec; 
    validation_data[  873] = 'h00002ee8; 
    validation_data[  874] = 'h00002e13; 
    validation_data[  875] = 'h00003b9f; 
    validation_data[  876] = 'h00003b37; 
    validation_data[  877] = 'h000002a5; 
    validation_data[  878] = 'h00001c82; 
    validation_data[  879] = 'h000000b5; 
    validation_data[  880] = 'h00003d3b; 
    validation_data[  881] = 'h000012b1; 
    validation_data[  882] = 'h00000703; 
    validation_data[  883] = 'h00000327; 
    validation_data[  884] = 'h0000323d; 
    validation_data[  885] = 'h00002cad; 
    validation_data[  886] = 'h00003d9c; 
    validation_data[  887] = 'h00003900; 
    validation_data[  888] = 'h000028f9; 
    validation_data[  889] = 'h00003757; 
    validation_data[  890] = 'h00003f5e; 
    validation_data[  891] = 'h000006d2; 
    validation_data[  892] = 'h00000133; 
    validation_data[  893] = 'h0000195f; 
    validation_data[  894] = 'h00002beb; 
    validation_data[  895] = 'h00002bfb; 
    validation_data[  896] = 'h00003733; 
    validation_data[  897] = 'h00000ba1; 
    validation_data[  898] = 'h00001f9f; 
    validation_data[  899] = 'h00002aa8; 
    validation_data[  900] = 'h00000659; 
    validation_data[  901] = 'h00001bd9; 
    validation_data[  902] = 'h00001840; 
    validation_data[  903] = 'h00001d71; 
    validation_data[  904] = 'h00002685; 
    validation_data[  905] = 'h00002c3a; 
    validation_data[  906] = 'h00001217; 
    validation_data[  907] = 'h000021cd; 
    validation_data[  908] = 'h00003c06; 
    validation_data[  909] = 'h00002881; 
    validation_data[  910] = 'h0000111a; 
    validation_data[  911] = 'h00003cca; 
    validation_data[  912] = 'h00001d0a; 
    validation_data[  913] = 'h00001ec5; 
    validation_data[  914] = 'h000034d0; 
    validation_data[  915] = 'h000033ac; 
    validation_data[  916] = 'h0000196d; 
    validation_data[  917] = 'h00003267; 
    validation_data[  918] = 'h00002491; 
    validation_data[  919] = 'h00002a81; 
    validation_data[  920] = 'h000039f4; 
    validation_data[  921] = 'h00002295; 
    validation_data[  922] = 'h00003a7b; 
    validation_data[  923] = 'h0000073a; 
    validation_data[  924] = 'h000028f3; 
    validation_data[  925] = 'h0000354b; 
    validation_data[  926] = 'h00001749; 
    validation_data[  927] = 'h00001d5a; 
    validation_data[  928] = 'h0000348c; 
    validation_data[  929] = 'h00000834; 
    validation_data[  930] = 'h00000cd1; 
    validation_data[  931] = 'h00001f44; 
    validation_data[  932] = 'h00002dec; 
    validation_data[  933] = 'h000019b3; 
    validation_data[  934] = 'h0000301d; 
    validation_data[  935] = 'h000036fc; 
    validation_data[  936] = 'h000022dc; 
    validation_data[  937] = 'h00001783; 
    validation_data[  938] = 'h00002094; 
    validation_data[  939] = 'h00000a6f; 
    validation_data[  940] = 'h00003d9b; 
    validation_data[  941] = 'h0000347b; 
    validation_data[  942] = 'h0000034a; 
    validation_data[  943] = 'h000004c9; 
    validation_data[  944] = 'h000021eb; 
    validation_data[  945] = 'h000010a5; 
    validation_data[  946] = 'h00003706; 
    validation_data[  947] = 'h00000056; 
    validation_data[  948] = 'h00001441; 
    validation_data[  949] = 'h000026ef; 
    validation_data[  950] = 'h00001d6d; 
    validation_data[  951] = 'h00001371; 
    validation_data[  952] = 'h00001dad; 
    validation_data[  953] = 'h000036d5; 
    validation_data[  954] = 'h00003118; 
    validation_data[  955] = 'h000039d2; 
    validation_data[  956] = 'h00002357; 
    validation_data[  957] = 'h0000337f; 
    validation_data[  958] = 'h00000c5b; 
    validation_data[  959] = 'h00003ba5; 
    validation_data[  960] = 'h0000353b; 
    validation_data[  961] = 'h00002dfe; 
    validation_data[  962] = 'h00002f14; 
    validation_data[  963] = 'h00003004; 
    validation_data[  964] = 'h00002483; 
    validation_data[  965] = 'h00002db4; 
    validation_data[  966] = 'h000025c7; 
    validation_data[  967] = 'h00003f9f; 
    validation_data[  968] = 'h00000773; 
    validation_data[  969] = 'h00003a1c; 
    validation_data[  970] = 'h00001ed1; 
    validation_data[  971] = 'h00001149; 
    validation_data[  972] = 'h00003fea; 
    validation_data[  973] = 'h00003f6e; 
    validation_data[  974] = 'h00003686; 
    validation_data[  975] = 'h00000206; 
    validation_data[  976] = 'h00002b95; 
    validation_data[  977] = 'h00000b83; 
    validation_data[  978] = 'h000008cd; 
    validation_data[  979] = 'h00003df5; 
    validation_data[  980] = 'h0000158e; 
    validation_data[  981] = 'h000005d9; 
    validation_data[  982] = 'h0000392b; 
    validation_data[  983] = 'h00000a67; 
    validation_data[  984] = 'h00001260; 
    validation_data[  985] = 'h000017fe; 
    validation_data[  986] = 'h00003a2d; 
    validation_data[  987] = 'h00001c18; 
    validation_data[  988] = 'h00002f0a; 
    validation_data[  989] = 'h000009e9; 
    validation_data[  990] = 'h0000304d; 
    validation_data[  991] = 'h00003a8f; 
    validation_data[  992] = 'h000029ac; 
    validation_data[  993] = 'h00000c42; 
    validation_data[  994] = 'h00000a2e; 
    validation_data[  995] = 'h000032b3; 
    validation_data[  996] = 'h000013fb; 
    validation_data[  997] = 'h00001ff0; 
    validation_data[  998] = 'h00000973; 
    validation_data[  999] = 'h00002b2c; 
    validation_data[ 1000] = 'h00000d26; 
    validation_data[ 1001] = 'h0000323a; 
    validation_data[ 1002] = 'h00002581; 
    validation_data[ 1003] = 'h00001aaa; 
    validation_data[ 1004] = 'h00000138; 
    validation_data[ 1005] = 'h00001134; 
    validation_data[ 1006] = 'h00000f2a; 
    validation_data[ 1007] = 'h00001c40; 
    validation_data[ 1008] = 'h00003ec4; 
    validation_data[ 1009] = 'h00003584; 
    validation_data[ 1010] = 'h000037aa; 
    validation_data[ 1011] = 'h00001db1; 
    validation_data[ 1012] = 'h00001876; 
    validation_data[ 1013] = 'h00003f05; 
    validation_data[ 1014] = 'h00003526; 
    validation_data[ 1015] = 'h000033e1; 
    validation_data[ 1016] = 'h00000eb8; 
    validation_data[ 1017] = 'h000011c3; 
    validation_data[ 1018] = 'h00002ce5; 
    validation_data[ 1019] = 'h00003f78; 
    validation_data[ 1020] = 'h00002b25; 
    validation_data[ 1021] = 'h000015df; 
    validation_data[ 1022] = 'h000030ec; 
    validation_data[ 1023] = 'h00002b40; 
    validation_data[ 1024] = 'h00000760; 
    validation_data[ 1025] = 'h00001941; 
    validation_data[ 1026] = 'h00001fd4; 
    validation_data[ 1027] = 'h00000165; 
    validation_data[ 1028] = 'h000013ff; 
    validation_data[ 1029] = 'h00001b8d; 
    validation_data[ 1030] = 'h000002be; 
    validation_data[ 1031] = 'h0000202f; 
    validation_data[ 1032] = 'h000029cf; 
    validation_data[ 1033] = 'h00003c9c; 
    validation_data[ 1034] = 'h0000325c; 
    validation_data[ 1035] = 'h00003fc6; 
    validation_data[ 1036] = 'h0000268b; 
    validation_data[ 1037] = 'h0000282f; 
    validation_data[ 1038] = 'h000036d1; 
    validation_data[ 1039] = 'h0000011b; 
    validation_data[ 1040] = 'h000007db; 
    validation_data[ 1041] = 'h00001854; 
    validation_data[ 1042] = 'h00000dcb; 
    validation_data[ 1043] = 'h00001bc0; 
    validation_data[ 1044] = 'h000038aa; 
    validation_data[ 1045] = 'h00003af5; 
    validation_data[ 1046] = 'h0000203e; 
    validation_data[ 1047] = 'h0000105d; 
    validation_data[ 1048] = 'h00003491; 
    validation_data[ 1049] = 'h0000306f; 
    validation_data[ 1050] = 'h00001a5c; 
    validation_data[ 1051] = 'h00002920; 
    validation_data[ 1052] = 'h00001856; 
    validation_data[ 1053] = 'h00001989; 
    validation_data[ 1054] = 'h0000259a; 
    validation_data[ 1055] = 'h000019da; 
    validation_data[ 1056] = 'h00003f60; 
    validation_data[ 1057] = 'h00003b52; 
    validation_data[ 1058] = 'h00002949; 
    validation_data[ 1059] = 'h000016d4; 
    validation_data[ 1060] = 'h00002188; 
    validation_data[ 1061] = 'h000012fa; 
    validation_data[ 1062] = 'h0000348f; 
    validation_data[ 1063] = 'h0000164c; 
    validation_data[ 1064] = 'h0000381f; 
    validation_data[ 1065] = 'h00001f95; 
    validation_data[ 1066] = 'h000032ee; 
    validation_data[ 1067] = 'h00003e20; 
    validation_data[ 1068] = 'h00000e69; 
    validation_data[ 1069] = 'h00001c21; 
    validation_data[ 1070] = 'h0000006d; 
    validation_data[ 1071] = 'h00001634; 
    validation_data[ 1072] = 'h0000166a; 
    validation_data[ 1073] = 'h00003a8e; 
    validation_data[ 1074] = 'h00003738; 
    validation_data[ 1075] = 'h00001946; 
    validation_data[ 1076] = 'h00002d5f; 
    validation_data[ 1077] = 'h00001963; 
    validation_data[ 1078] = 'h000034c7; 
    validation_data[ 1079] = 'h0000379b; 
    validation_data[ 1080] = 'h000025bc; 
    validation_data[ 1081] = 'h00001a5d; 
    validation_data[ 1082] = 'h00003151; 
    validation_data[ 1083] = 'h00001f91; 
    validation_data[ 1084] = 'h00001d19; 
    validation_data[ 1085] = 'h000027b3; 
    validation_data[ 1086] = 'h0000362c; 
    validation_data[ 1087] = 'h0000268e; 
    validation_data[ 1088] = 'h000021f4; 
    validation_data[ 1089] = 'h00002480; 
    validation_data[ 1090] = 'h00003d3c; 
    validation_data[ 1091] = 'h00001e53; 
    validation_data[ 1092] = 'h0000242b; 
    validation_data[ 1093] = 'h00000812; 
    validation_data[ 1094] = 'h0000068f; 
    validation_data[ 1095] = 'h0000184b; 
    validation_data[ 1096] = 'h00000a21; 
    validation_data[ 1097] = 'h00000cef; 
    validation_data[ 1098] = 'h0000337e; 
    validation_data[ 1099] = 'h0000170c; 
    validation_data[ 1100] = 'h00003001; 
    validation_data[ 1101] = 'h00003bfd; 
    validation_data[ 1102] = 'h00002d68; 
    validation_data[ 1103] = 'h0000109a; 
    validation_data[ 1104] = 'h000014f6; 
    validation_data[ 1105] = 'h00003ab9; 
    validation_data[ 1106] = 'h0000074d; 
    validation_data[ 1107] = 'h000029e4; 
    validation_data[ 1108] = 'h00001466; 
    validation_data[ 1109] = 'h00002ced; 
    validation_data[ 1110] = 'h000010f5; 
    validation_data[ 1111] = 'h00001fbf; 
    validation_data[ 1112] = 'h00001d76; 
    validation_data[ 1113] = 'h0000311a; 
    validation_data[ 1114] = 'h000002d1; 
    validation_data[ 1115] = 'h00003d65; 
    validation_data[ 1116] = 'h00003e50; 
    validation_data[ 1117] = 'h00003e03; 
    validation_data[ 1118] = 'h00003e02; 
    validation_data[ 1119] = 'h00000dd5; 
    validation_data[ 1120] = 'h00003b4c; 
    validation_data[ 1121] = 'h00001f86; 
    validation_data[ 1122] = 'h000033a9; 
    validation_data[ 1123] = 'h0000100a; 
    validation_data[ 1124] = 'h00002986; 
    validation_data[ 1125] = 'h00001963; 
    validation_data[ 1126] = 'h00003f5a; 
    validation_data[ 1127] = 'h00001c03; 
    validation_data[ 1128] = 'h00003b5a; 
    validation_data[ 1129] = 'h00000bf5; 
    validation_data[ 1130] = 'h0000193c; 
    validation_data[ 1131] = 'h00003755; 
    validation_data[ 1132] = 'h00001137; 
    validation_data[ 1133] = 'h0000178b; 
    validation_data[ 1134] = 'h00002201; 
    validation_data[ 1135] = 'h0000282d; 
    validation_data[ 1136] = 'h00002366; 
    validation_data[ 1137] = 'h000004b9; 
    validation_data[ 1138] = 'h00001989; 
    validation_data[ 1139] = 'h00003ee7; 
    validation_data[ 1140] = 'h0000362b; 
    validation_data[ 1141] = 'h00002115; 
    validation_data[ 1142] = 'h00000cd8; 
    validation_data[ 1143] = 'h00000a00; 
    validation_data[ 1144] = 'h00001709; 
    validation_data[ 1145] = 'h000024fe; 
    validation_data[ 1146] = 'h00000b26; 
    validation_data[ 1147] = 'h00003ceb; 
    validation_data[ 1148] = 'h0000379b; 
    validation_data[ 1149] = 'h00003414; 
    validation_data[ 1150] = 'h00001599; 
    validation_data[ 1151] = 'h00001e7d; 
    validation_data[ 1152] = 'h00000dc5; 
    validation_data[ 1153] = 'h00002eba; 
    validation_data[ 1154] = 'h00002305; 
    validation_data[ 1155] = 'h0000165f; 
    validation_data[ 1156] = 'h00001a98; 
    validation_data[ 1157] = 'h00001af0; 
    validation_data[ 1158] = 'h00001d0e; 
    validation_data[ 1159] = 'h00003aed; 
    validation_data[ 1160] = 'h00002135; 
    validation_data[ 1161] = 'h0000331f; 
    validation_data[ 1162] = 'h00002d54; 
    validation_data[ 1163] = 'h00003606; 
    validation_data[ 1164] = 'h00002e73; 
    validation_data[ 1165] = 'h00000673; 
    validation_data[ 1166] = 'h00000f58; 
    validation_data[ 1167] = 'h00001dc7; 
    validation_data[ 1168] = 'h000003ae; 
    validation_data[ 1169] = 'h00001cce; 
    validation_data[ 1170] = 'h00003ecb; 
    validation_data[ 1171] = 'h000031bc; 
    validation_data[ 1172] = 'h0000226f; 
    validation_data[ 1173] = 'h000006a8; 
    validation_data[ 1174] = 'h00002ec1; 
    validation_data[ 1175] = 'h00000a83; 
    validation_data[ 1176] = 'h00003e5e; 
    validation_data[ 1177] = 'h00003ba1; 
    validation_data[ 1178] = 'h00000cdf; 
    validation_data[ 1179] = 'h00003c30; 
    validation_data[ 1180] = 'h00001534; 
    validation_data[ 1181] = 'h0000274e; 
    validation_data[ 1182] = 'h00002047; 
    validation_data[ 1183] = 'h00002a8c; 
    validation_data[ 1184] = 'h000016ea; 
    validation_data[ 1185] = 'h00001cde; 
    validation_data[ 1186] = 'h0000108b; 
    validation_data[ 1187] = 'h000020d5; 
    validation_data[ 1188] = 'h00001f3c; 
    validation_data[ 1189] = 'h00002873; 
    validation_data[ 1190] = 'h000008e7; 
    validation_data[ 1191] = 'h00002dfb; 
    validation_data[ 1192] = 'h00003495; 
    validation_data[ 1193] = 'h00001888; 
    validation_data[ 1194] = 'h0000150a; 
    validation_data[ 1195] = 'h0000373d; 
    validation_data[ 1196] = 'h00003b0c; 
    validation_data[ 1197] = 'h00000965; 
    validation_data[ 1198] = 'h000027e0; 
    validation_data[ 1199] = 'h00001cb7; 
    validation_data[ 1200] = 'h0000053d; 
    validation_data[ 1201] = 'h00001a42; 
    validation_data[ 1202] = 'h00003d36; 
    validation_data[ 1203] = 'h0000131a; 
    validation_data[ 1204] = 'h000003c6; 
    validation_data[ 1205] = 'h0000371b; 
    validation_data[ 1206] = 'h00002572; 
    validation_data[ 1207] = 'h00002da5; 
    validation_data[ 1208] = 'h000020cc; 
    validation_data[ 1209] = 'h00003cd9; 
    validation_data[ 1210] = 'h000020ea; 
    validation_data[ 1211] = 'h000006ae; 
    validation_data[ 1212] = 'h00000e85; 
    validation_data[ 1213] = 'h0000114e; 
    validation_data[ 1214] = 'h00001541; 
    validation_data[ 1215] = 'h0000313d; 
    validation_data[ 1216] = 'h00000e48; 
    validation_data[ 1217] = 'h0000138b; 
    validation_data[ 1218] = 'h0000131b; 
    validation_data[ 1219] = 'h0000151a; 
    validation_data[ 1220] = 'h00000552; 
    validation_data[ 1221] = 'h00000227; 
    validation_data[ 1222] = 'h00002daf; 
    validation_data[ 1223] = 'h00001f7d; 
    validation_data[ 1224] = 'h000034ee; 
    validation_data[ 1225] = 'h00003361; 
    validation_data[ 1226] = 'h0000296b; 
    validation_data[ 1227] = 'h000010d5; 
    validation_data[ 1228] = 'h000005a8; 
    validation_data[ 1229] = 'h000017df; 
    validation_data[ 1230] = 'h00003f76; 
    validation_data[ 1231] = 'h000033c2; 
    validation_data[ 1232] = 'h00003534; 
    validation_data[ 1233] = 'h00000d16; 
    validation_data[ 1234] = 'h00003497; 
    validation_data[ 1235] = 'h00001697; 
    validation_data[ 1236] = 'h00000aba; 
    validation_data[ 1237] = 'h00000b0f; 
    validation_data[ 1238] = 'h000023db; 
    validation_data[ 1239] = 'h00000d84; 
    validation_data[ 1240] = 'h000038ab; 
    validation_data[ 1241] = 'h00003066; 
    validation_data[ 1242] = 'h0000277b; 
    validation_data[ 1243] = 'h000031bb; 
    validation_data[ 1244] = 'h000015b5; 
    validation_data[ 1245] = 'h00002ac4; 
    validation_data[ 1246] = 'h00003758; 
    validation_data[ 1247] = 'h000015bc; 
    validation_data[ 1248] = 'h00001127; 
    validation_data[ 1249] = 'h00000b8b; 
    validation_data[ 1250] = 'h00001581; 
    validation_data[ 1251] = 'h00003451; 
    validation_data[ 1252] = 'h000036dc; 
    validation_data[ 1253] = 'h00003901; 
    validation_data[ 1254] = 'h000019b9; 
    validation_data[ 1255] = 'h0000162b; 
    validation_data[ 1256] = 'h0000346a; 
    validation_data[ 1257] = 'h00002a61; 
    validation_data[ 1258] = 'h00001448; 
    validation_data[ 1259] = 'h00003eb1; 
    validation_data[ 1260] = 'h00002c47; 
    validation_data[ 1261] = 'h00001427; 
    validation_data[ 1262] = 'h000007cd; 
    validation_data[ 1263] = 'h00002b7c; 
    validation_data[ 1264] = 'h000037db; 
    validation_data[ 1265] = 'h00003d21; 
    validation_data[ 1266] = 'h00000cf6; 
    validation_data[ 1267] = 'h00001261; 
    validation_data[ 1268] = 'h00001f03; 
    validation_data[ 1269] = 'h000022ec; 
    validation_data[ 1270] = 'h00003954; 
    validation_data[ 1271] = 'h000034ed; 
    validation_data[ 1272] = 'h00002683; 
    validation_data[ 1273] = 'h00003a36; 
    validation_data[ 1274] = 'h000039db; 
    validation_data[ 1275] = 'h00001ca0; 
    validation_data[ 1276] = 'h0000082b; 
    validation_data[ 1277] = 'h000000a8; 
    validation_data[ 1278] = 'h00002e56; 
    validation_data[ 1279] = 'h0000121f; 
    validation_data[ 1280] = 'h00000598; 
    validation_data[ 1281] = 'h00002764; 
    validation_data[ 1282] = 'h00001d8a; 
    validation_data[ 1283] = 'h00002979; 
    validation_data[ 1284] = 'h00001e89; 
    validation_data[ 1285] = 'h00002590; 
    validation_data[ 1286] = 'h00003ff5; 
    validation_data[ 1287] = 'h00003fc3; 
    validation_data[ 1288] = 'h00001a43; 
    validation_data[ 1289] = 'h00001e7f; 
    validation_data[ 1290] = 'h00002409; 
    validation_data[ 1291] = 'h00003a77; 
    validation_data[ 1292] = 'h00003114; 
    validation_data[ 1293] = 'h000010ba; 
    validation_data[ 1294] = 'h000010dc; 
    validation_data[ 1295] = 'h00000b54; 
    validation_data[ 1296] = 'h00003e28; 
    validation_data[ 1297] = 'h000021ba; 
    validation_data[ 1298] = 'h00001a18; 
    validation_data[ 1299] = 'h0000164b; 
    validation_data[ 1300] = 'h00001c5b; 
    validation_data[ 1301] = 'h000007fa; 
    validation_data[ 1302] = 'h00000553; 
    validation_data[ 1303] = 'h000029c9; 
    validation_data[ 1304] = 'h000012a3; 
    validation_data[ 1305] = 'h0000144d; 
    validation_data[ 1306] = 'h000006d9; 
    validation_data[ 1307] = 'h00000951; 
    validation_data[ 1308] = 'h000037c2; 
    validation_data[ 1309] = 'h00002f15; 
    validation_data[ 1310] = 'h00001be9; 
    validation_data[ 1311] = 'h0000045b; 
    validation_data[ 1312] = 'h00001eeb; 
    validation_data[ 1313] = 'h000023a5; 
    validation_data[ 1314] = 'h00003d52; 
    validation_data[ 1315] = 'h00002500; 
    validation_data[ 1316] = 'h00003561; 
    validation_data[ 1317] = 'h000011c5; 
    validation_data[ 1318] = 'h00000a37; 
    validation_data[ 1319] = 'h00000066; 
    validation_data[ 1320] = 'h00003abc; 
    validation_data[ 1321] = 'h00000eb4; 
    validation_data[ 1322] = 'h00001212; 
    validation_data[ 1323] = 'h000007de; 
    validation_data[ 1324] = 'h00001ca3; 
    validation_data[ 1325] = 'h00001408; 
    validation_data[ 1326] = 'h0000268e; 
    validation_data[ 1327] = 'h00003637; 
    validation_data[ 1328] = 'h00000c9f; 
    validation_data[ 1329] = 'h00001a18; 
    validation_data[ 1330] = 'h000030b3; 
    validation_data[ 1331] = 'h00003cb5; 
    validation_data[ 1332] = 'h0000099a; 
    validation_data[ 1333] = 'h00000772; 
    validation_data[ 1334] = 'h0000034d; 
    validation_data[ 1335] = 'h000016b1; 
    validation_data[ 1336] = 'h00003854; 
    validation_data[ 1337] = 'h000006bc; 
    validation_data[ 1338] = 'h000003ae; 
    validation_data[ 1339] = 'h0000175a; 
    validation_data[ 1340] = 'h00003285; 
    validation_data[ 1341] = 'h000013df; 
    validation_data[ 1342] = 'h00003b7f; 
    validation_data[ 1343] = 'h00002e8d; 
    validation_data[ 1344] = 'h00002ba3; 
    validation_data[ 1345] = 'h00003bcf; 
    validation_data[ 1346] = 'h00001b5c; 
    validation_data[ 1347] = 'h00002100; 
    validation_data[ 1348] = 'h00000e4f; 
    validation_data[ 1349] = 'h00002062; 
    validation_data[ 1350] = 'h000031c7; 
    validation_data[ 1351] = 'h00003812; 
    validation_data[ 1352] = 'h00002a54; 
    validation_data[ 1353] = 'h00000e09; 
    validation_data[ 1354] = 'h000039ec; 
    validation_data[ 1355] = 'h000027c7; 
    validation_data[ 1356] = 'h00000694; 
    validation_data[ 1357] = 'h00002c07; 
    validation_data[ 1358] = 'h00001888; 
    validation_data[ 1359] = 'h00003c34; 
    validation_data[ 1360] = 'h00002227; 
    validation_data[ 1361] = 'h000004ec; 
    validation_data[ 1362] = 'h0000179d; 
    validation_data[ 1363] = 'h00002716; 
    validation_data[ 1364] = 'h00002233; 
    validation_data[ 1365] = 'h00003a7a; 
    validation_data[ 1366] = 'h00001f07; 
    validation_data[ 1367] = 'h00000387; 
    validation_data[ 1368] = 'h000012f5; 
    validation_data[ 1369] = 'h000021ba; 
    validation_data[ 1370] = 'h00003067; 
    validation_data[ 1371] = 'h0000204c; 
    validation_data[ 1372] = 'h00003bdb; 
    validation_data[ 1373] = 'h00001fa6; 
    validation_data[ 1374] = 'h0000255e; 
    validation_data[ 1375] = 'h00002679; 
    validation_data[ 1376] = 'h000036f0; 
    validation_data[ 1377] = 'h00002240; 
    validation_data[ 1378] = 'h0000168a; 
    validation_data[ 1379] = 'h000004c8; 
    validation_data[ 1380] = 'h00003d06; 
    validation_data[ 1381] = 'h00001d4c; 
    validation_data[ 1382] = 'h00003e31; 
    validation_data[ 1383] = 'h00000175; 
    validation_data[ 1384] = 'h00003b3d; 
    validation_data[ 1385] = 'h000008e4; 
    validation_data[ 1386] = 'h000009c0; 
    validation_data[ 1387] = 'h00000799; 
    validation_data[ 1388] = 'h0000015f; 
    validation_data[ 1389] = 'h00001fcd; 
    validation_data[ 1390] = 'h0000110a; 
    validation_data[ 1391] = 'h00003354; 
    validation_data[ 1392] = 'h0000215b; 
    validation_data[ 1393] = 'h00001efe; 
    validation_data[ 1394] = 'h000026c0; 
    validation_data[ 1395] = 'h0000003d; 
    validation_data[ 1396] = 'h00003fa2; 
    validation_data[ 1397] = 'h000019c8; 
    validation_data[ 1398] = 'h0000157e; 
    validation_data[ 1399] = 'h00001351; 
    validation_data[ 1400] = 'h000015e4; 
    validation_data[ 1401] = 'h00002a30; 
    validation_data[ 1402] = 'h000004a6; 
    validation_data[ 1403] = 'h00000607; 
    validation_data[ 1404] = 'h000011b5; 
    validation_data[ 1405] = 'h00001f48; 
    validation_data[ 1406] = 'h0000004a; 
    validation_data[ 1407] = 'h00003d31; 
    validation_data[ 1408] = 'h00002e63; 
    validation_data[ 1409] = 'h00002f24; 
    validation_data[ 1410] = 'h000031d2; 
    validation_data[ 1411] = 'h00001015; 
    validation_data[ 1412] = 'h00000c28; 
    validation_data[ 1413] = 'h000029d7; 
    validation_data[ 1414] = 'h00002a06; 
    validation_data[ 1415] = 'h00000bfe; 
    validation_data[ 1416] = 'h00003178; 
    validation_data[ 1417] = 'h0000295b; 
    validation_data[ 1418] = 'h00002909; 
    validation_data[ 1419] = 'h000027c3; 
    validation_data[ 1420] = 'h00001c38; 
    validation_data[ 1421] = 'h00000550; 
    validation_data[ 1422] = 'h0000294d; 
    validation_data[ 1423] = 'h00001130; 
    validation_data[ 1424] = 'h000004c1; 
    validation_data[ 1425] = 'h000015a3; 
    validation_data[ 1426] = 'h000023e8; 
    validation_data[ 1427] = 'h00003ee5; 
    validation_data[ 1428] = 'h00002b0e; 
    validation_data[ 1429] = 'h00000a0d; 
    validation_data[ 1430] = 'h00001ded; 
    validation_data[ 1431] = 'h00001822; 
    validation_data[ 1432] = 'h00003e22; 
    validation_data[ 1433] = 'h000028be; 
    validation_data[ 1434] = 'h00000431; 
    validation_data[ 1435] = 'h00001af7; 
    validation_data[ 1436] = 'h000002f8; 
    validation_data[ 1437] = 'h0000028b; 
    validation_data[ 1438] = 'h00000b47; 
    validation_data[ 1439] = 'h0000040e; 
    validation_data[ 1440] = 'h00001f89; 
    validation_data[ 1441] = 'h00001f6d; 
    validation_data[ 1442] = 'h00003a6c; 
    validation_data[ 1443] = 'h000033bc; 
    validation_data[ 1444] = 'h00001fab; 
    validation_data[ 1445] = 'h00000292; 
    validation_data[ 1446] = 'h00003815; 
    validation_data[ 1447] = 'h00001b12; 
    validation_data[ 1448] = 'h00003ff7; 
    validation_data[ 1449] = 'h00001199; 
    validation_data[ 1450] = 'h00003f90; 
    validation_data[ 1451] = 'h00002144; 
    validation_data[ 1452] = 'h00001149; 
    validation_data[ 1453] = 'h00001bca; 
    validation_data[ 1454] = 'h00001eba; 
    validation_data[ 1455] = 'h00003665; 
    validation_data[ 1456] = 'h00000a5c; 
    validation_data[ 1457] = 'h00001c1c; 
    validation_data[ 1458] = 'h00003719; 
    validation_data[ 1459] = 'h00001299; 
    validation_data[ 1460] = 'h00003419; 
    validation_data[ 1461] = 'h0000043f; 
    validation_data[ 1462] = 'h00000cd4; 
    validation_data[ 1463] = 'h000004a6; 
    validation_data[ 1464] = 'h000008b8; 
    validation_data[ 1465] = 'h000011c6; 
    validation_data[ 1466] = 'h00001f26; 
    validation_data[ 1467] = 'h00001e30; 
    validation_data[ 1468] = 'h0000013d; 
    validation_data[ 1469] = 'h000003ae; 
    validation_data[ 1470] = 'h00001c3a; 
    validation_data[ 1471] = 'h00000695; 
    validation_data[ 1472] = 'h000030e1; 
    validation_data[ 1473] = 'h00000cb9; 
    validation_data[ 1474] = 'h00002f06; 
    validation_data[ 1475] = 'h000032b9; 
    validation_data[ 1476] = 'h000012f2; 
    validation_data[ 1477] = 'h00002abc; 
    validation_data[ 1478] = 'h00001311; 
    validation_data[ 1479] = 'h000037b4; 
    validation_data[ 1480] = 'h00001a53; 
    validation_data[ 1481] = 'h0000230b; 
    validation_data[ 1482] = 'h00001789; 
    validation_data[ 1483] = 'h0000388e; 
    validation_data[ 1484] = 'h00001cd7; 
    validation_data[ 1485] = 'h0000295e; 
    validation_data[ 1486] = 'h00003f06; 
    validation_data[ 1487] = 'h00002a1a; 
    validation_data[ 1488] = 'h00000713; 
    validation_data[ 1489] = 'h000005e4; 
    validation_data[ 1490] = 'h00003fb3; 
    validation_data[ 1491] = 'h0000100a; 
    validation_data[ 1492] = 'h00003d68; 
    validation_data[ 1493] = 'h00000b72; 
    validation_data[ 1494] = 'h00003a21; 
    validation_data[ 1495] = 'h00002449; 
    validation_data[ 1496] = 'h000031b3; 
    validation_data[ 1497] = 'h000004fb; 
    validation_data[ 1498] = 'h00002025; 
    validation_data[ 1499] = 'h00000e19; 
    validation_data[ 1500] = 'h00003d32; 
    validation_data[ 1501] = 'h00001bec; 
    validation_data[ 1502] = 'h000006f6; 
    validation_data[ 1503] = 'h00001819; 
    validation_data[ 1504] = 'h00000886; 
    validation_data[ 1505] = 'h00003863; 
    validation_data[ 1506] = 'h000003d0; 
    validation_data[ 1507] = 'h00000878; 
    validation_data[ 1508] = 'h0000253c; 
    validation_data[ 1509] = 'h0000075a; 
    validation_data[ 1510] = 'h0000253d; 
    validation_data[ 1511] = 'h000020ce; 
    validation_data[ 1512] = 'h00001902; 
    validation_data[ 1513] = 'h0000220d; 
    validation_data[ 1514] = 'h000033d2; 
    validation_data[ 1515] = 'h0000168b; 
    validation_data[ 1516] = 'h00003ae9; 
    validation_data[ 1517] = 'h000001b0; 
    validation_data[ 1518] = 'h00003d6e; 
    validation_data[ 1519] = 'h00001864; 
    validation_data[ 1520] = 'h000028d4; 
    validation_data[ 1521] = 'h0000054d; 
    validation_data[ 1522] = 'h00003f5b; 
    validation_data[ 1523] = 'h00001cae; 
    validation_data[ 1524] = 'h00001f48; 
    validation_data[ 1525] = 'h00002f54; 
    validation_data[ 1526] = 'h00000988; 
    validation_data[ 1527] = 'h0000279d; 
    validation_data[ 1528] = 'h0000399c; 
    validation_data[ 1529] = 'h00001f8f; 
    validation_data[ 1530] = 'h00001c31; 
    validation_data[ 1531] = 'h000013f8; 
    validation_data[ 1532] = 'h00002da5; 
    validation_data[ 1533] = 'h00003926; 
    validation_data[ 1534] = 'h00001cc9; 
    validation_data[ 1535] = 'h000017eb; 
    validation_data[ 1536] = 'h0000259c; 
    validation_data[ 1537] = 'h00003ab1; 
    validation_data[ 1538] = 'h00003cd4; 
    validation_data[ 1539] = 'h000002c9; 
    validation_data[ 1540] = 'h00000c3f; 
    validation_data[ 1541] = 'h00003e78; 
    validation_data[ 1542] = 'h00002984; 
    validation_data[ 1543] = 'h00001b30; 
    validation_data[ 1544] = 'h00003d0c; 
    validation_data[ 1545] = 'h000027e2; 
    validation_data[ 1546] = 'h00002f9a; 
    validation_data[ 1547] = 'h000021a7; 
    validation_data[ 1548] = 'h00000b5a; 
    validation_data[ 1549] = 'h000004b5; 
    validation_data[ 1550] = 'h0000057c; 
    validation_data[ 1551] = 'h000022ec; 
    validation_data[ 1552] = 'h00002d3c; 
    validation_data[ 1553] = 'h00002cb6; 
    validation_data[ 1554] = 'h00003f41; 
    validation_data[ 1555] = 'h00002460; 
    validation_data[ 1556] = 'h00000edf; 
    validation_data[ 1557] = 'h0000086d; 
    validation_data[ 1558] = 'h0000106a; 
    validation_data[ 1559] = 'h000035e3; 
    validation_data[ 1560] = 'h00003f18; 
    validation_data[ 1561] = 'h00002c16; 
    validation_data[ 1562] = 'h00002a71; 
    validation_data[ 1563] = 'h00000ca0; 
    validation_data[ 1564] = 'h000020a8; 
    validation_data[ 1565] = 'h00003d55; 
    validation_data[ 1566] = 'h00001d12; 
    validation_data[ 1567] = 'h0000081c; 
    validation_data[ 1568] = 'h00002df3; 
    validation_data[ 1569] = 'h000022d9; 
    validation_data[ 1570] = 'h0000088d; 
    validation_data[ 1571] = 'h000009bd; 
    validation_data[ 1572] = 'h00000a6c; 
    validation_data[ 1573] = 'h00000442; 
    validation_data[ 1574] = 'h000006cf; 
    validation_data[ 1575] = 'h00002b4d; 
    validation_data[ 1576] = 'h000003c6; 
    validation_data[ 1577] = 'h000037a9; 
    validation_data[ 1578] = 'h00000632; 
    validation_data[ 1579] = 'h000001b9; 
    validation_data[ 1580] = 'h00002d1e; 
    validation_data[ 1581] = 'h00000e0f; 
    validation_data[ 1582] = 'h00002cc7; 
    validation_data[ 1583] = 'h0000383a; 
    validation_data[ 1584] = 'h000037a0; 
    validation_data[ 1585] = 'h000005e7; 
    validation_data[ 1586] = 'h000012e6; 
    validation_data[ 1587] = 'h000028e9; 
    validation_data[ 1588] = 'h000006f2; 
    validation_data[ 1589] = 'h000020f1; 
    validation_data[ 1590] = 'h00002ddf; 
    validation_data[ 1591] = 'h00002721; 
    validation_data[ 1592] = 'h00001af3; 
    validation_data[ 1593] = 'h00002104; 
    validation_data[ 1594] = 'h00000be7; 
    validation_data[ 1595] = 'h00002fce; 
    validation_data[ 1596] = 'h00000523; 
    validation_data[ 1597] = 'h00003967; 
    validation_data[ 1598] = 'h00000644; 
    validation_data[ 1599] = 'h00001c67; 
    validation_data[ 1600] = 'h000031af; 
    validation_data[ 1601] = 'h00001967; 
    validation_data[ 1602] = 'h000010b9; 
    validation_data[ 1603] = 'h00001777; 
    validation_data[ 1604] = 'h000009a6; 
    validation_data[ 1605] = 'h00001858; 
    validation_data[ 1606] = 'h00001ad8; 
    validation_data[ 1607] = 'h000016d5; 
    validation_data[ 1608] = 'h0000050c; 
    validation_data[ 1609] = 'h000009ed; 
    validation_data[ 1610] = 'h00001ab3; 
    validation_data[ 1611] = 'h000031b3; 
    validation_data[ 1612] = 'h000004b6; 
    validation_data[ 1613] = 'h000007f7; 
    validation_data[ 1614] = 'h000036aa; 
    validation_data[ 1615] = 'h00003989; 
    validation_data[ 1616] = 'h00003867; 
    validation_data[ 1617] = 'h0000090f; 
    validation_data[ 1618] = 'h00003165; 
    validation_data[ 1619] = 'h00003f1f; 
    validation_data[ 1620] = 'h00002337; 
    validation_data[ 1621] = 'h00002ba5; 
    validation_data[ 1622] = 'h0000142b; 
    validation_data[ 1623] = 'h0000217f; 
    validation_data[ 1624] = 'h0000352d; 
    validation_data[ 1625] = 'h000010e2; 
    validation_data[ 1626] = 'h0000169c; 
    validation_data[ 1627] = 'h00003b5b; 
    validation_data[ 1628] = 'h00001813; 
    validation_data[ 1629] = 'h00001a2f; 
    validation_data[ 1630] = 'h000036ef; 
    validation_data[ 1631] = 'h00002d7b; 
    validation_data[ 1632] = 'h0000049e; 
    validation_data[ 1633] = 'h00002978; 
    validation_data[ 1634] = 'h0000175b; 
    validation_data[ 1635] = 'h00001558; 
    validation_data[ 1636] = 'h00002ee6; 
    validation_data[ 1637] = 'h00000c50; 
    validation_data[ 1638] = 'h00000422; 
    validation_data[ 1639] = 'h000003cb; 
    validation_data[ 1640] = 'h00002e79; 
    validation_data[ 1641] = 'h00003406; 
    validation_data[ 1642] = 'h00000579; 
    validation_data[ 1643] = 'h000017d8; 
    validation_data[ 1644] = 'h00002ad6; 
    validation_data[ 1645] = 'h00002840; 
    validation_data[ 1646] = 'h00003615; 
    validation_data[ 1647] = 'h00000e22; 
    validation_data[ 1648] = 'h000037fd; 
    validation_data[ 1649] = 'h000010dd; 
    validation_data[ 1650] = 'h000030a5; 
    validation_data[ 1651] = 'h00001b69; 
    validation_data[ 1652] = 'h00002e60; 
    validation_data[ 1653] = 'h00001aa0; 
    validation_data[ 1654] = 'h00000972; 
    validation_data[ 1655] = 'h0000095f; 
    validation_data[ 1656] = 'h00003d42; 
    validation_data[ 1657] = 'h00002226; 
    validation_data[ 1658] = 'h00002526; 
    validation_data[ 1659] = 'h000032ce; 
    validation_data[ 1660] = 'h0000338e; 
    validation_data[ 1661] = 'h000015f6; 
    validation_data[ 1662] = 'h00003219; 
    validation_data[ 1663] = 'h000008b6; 
    validation_data[ 1664] = 'h00003975; 
    validation_data[ 1665] = 'h00000667; 
    validation_data[ 1666] = 'h00003d6b; 
    validation_data[ 1667] = 'h00000dde; 
    validation_data[ 1668] = 'h00001d05; 
    validation_data[ 1669] = 'h00003f11; 
    validation_data[ 1670] = 'h00002d1d; 
    validation_data[ 1671] = 'h0000201e; 
    validation_data[ 1672] = 'h000002f1; 
    validation_data[ 1673] = 'h000017a3; 
    validation_data[ 1674] = 'h00003100; 
    validation_data[ 1675] = 'h00001724; 
    validation_data[ 1676] = 'h000034f1; 
    validation_data[ 1677] = 'h00000cc1; 
    validation_data[ 1678] = 'h00003407; 
    validation_data[ 1679] = 'h000028fc; 
    validation_data[ 1680] = 'h00002bff; 
    validation_data[ 1681] = 'h00003d9d; 
    validation_data[ 1682] = 'h000027d3; 
    validation_data[ 1683] = 'h00000df1; 
    validation_data[ 1684] = 'h00001408; 
    validation_data[ 1685] = 'h0000289b; 
    validation_data[ 1686] = 'h00002a29; 
    validation_data[ 1687] = 'h000033be; 
    validation_data[ 1688] = 'h00000236; 
    validation_data[ 1689] = 'h00003aaa; 
    validation_data[ 1690] = 'h00001254; 
    validation_data[ 1691] = 'h00001591; 
    validation_data[ 1692] = 'h0000078f; 
    validation_data[ 1693] = 'h000003c1; 
    validation_data[ 1694] = 'h0000038d; 
    validation_data[ 1695] = 'h00001e53; 
    validation_data[ 1696] = 'h000033ef; 
    validation_data[ 1697] = 'h000000c0; 
    validation_data[ 1698] = 'h00001bf7; 
    validation_data[ 1699] = 'h00002bbd; 
    validation_data[ 1700] = 'h0000397f; 
    validation_data[ 1701] = 'h00000b97; 
    validation_data[ 1702] = 'h00003fe1; 
    validation_data[ 1703] = 'h00000129; 
    validation_data[ 1704] = 'h00000680; 
    validation_data[ 1705] = 'h00001db5; 
    validation_data[ 1706] = 'h00002d72; 
    validation_data[ 1707] = 'h00002990; 
    validation_data[ 1708] = 'h000000ff; 
    validation_data[ 1709] = 'h00002b22; 
    validation_data[ 1710] = 'h00000de4; 
    validation_data[ 1711] = 'h000020d0; 
    validation_data[ 1712] = 'h000034d5; 
    validation_data[ 1713] = 'h00003276; 
    validation_data[ 1714] = 'h00000189; 
    validation_data[ 1715] = 'h0000232e; 
    validation_data[ 1716] = 'h00003ec4; 
    validation_data[ 1717] = 'h0000385b; 
    validation_data[ 1718] = 'h0000323f; 
    validation_data[ 1719] = 'h00000edd; 
    validation_data[ 1720] = 'h0000093f; 
    validation_data[ 1721] = 'h00000a70; 
    validation_data[ 1722] = 'h000034a8; 
    validation_data[ 1723] = 'h00001cd6; 
    validation_data[ 1724] = 'h00002e7d; 
    validation_data[ 1725] = 'h00003570; 
    validation_data[ 1726] = 'h00003b51; 
    validation_data[ 1727] = 'h00000067; 
    validation_data[ 1728] = 'h00000992; 
    validation_data[ 1729] = 'h00001a02; 
    validation_data[ 1730] = 'h000007e0; 
    validation_data[ 1731] = 'h00000009; 
    validation_data[ 1732] = 'h00000f17; 
    validation_data[ 1733] = 'h0000324d; 
    validation_data[ 1734] = 'h00000025; 
    validation_data[ 1735] = 'h00000a5e; 
    validation_data[ 1736] = 'h00000241; 
    validation_data[ 1737] = 'h00002e68; 
    validation_data[ 1738] = 'h00002110; 
    validation_data[ 1739] = 'h0000064e; 
    validation_data[ 1740] = 'h00003534; 
    validation_data[ 1741] = 'h00001d06; 
    validation_data[ 1742] = 'h000029d5; 
    validation_data[ 1743] = 'h000037b6; 
    validation_data[ 1744] = 'h000001af; 
    validation_data[ 1745] = 'h0000041b; 
    validation_data[ 1746] = 'h000023f8; 
    validation_data[ 1747] = 'h00003632; 
    validation_data[ 1748] = 'h000006e0; 
    validation_data[ 1749] = 'h000028a3; 
    validation_data[ 1750] = 'h00003ab2; 
    validation_data[ 1751] = 'h00000db8; 
    validation_data[ 1752] = 'h00002f99; 
    validation_data[ 1753] = 'h00003cb0; 
    validation_data[ 1754] = 'h000003a8; 
    validation_data[ 1755] = 'h0000347e; 
    validation_data[ 1756] = 'h00000724; 
    validation_data[ 1757] = 'h000002ac; 
    validation_data[ 1758] = 'h000007f9; 
    validation_data[ 1759] = 'h00000d8e; 
    validation_data[ 1760] = 'h0000080b; 
    validation_data[ 1761] = 'h0000264e; 
    validation_data[ 1762] = 'h00002e88; 
    validation_data[ 1763] = 'h00003527; 
    validation_data[ 1764] = 'h000004b2; 
    validation_data[ 1765] = 'h00002731; 
    validation_data[ 1766] = 'h0000211f; 
    validation_data[ 1767] = 'h00002802; 
    validation_data[ 1768] = 'h00000547; 
    validation_data[ 1769] = 'h00003249; 
    validation_data[ 1770] = 'h00003fa6; 
    validation_data[ 1771] = 'h00003476; 
    validation_data[ 1772] = 'h00000bb1; 
    validation_data[ 1773] = 'h000002a1; 
    validation_data[ 1774] = 'h00002598; 
    validation_data[ 1775] = 'h000025b4; 
    validation_data[ 1776] = 'h0000118b; 
    validation_data[ 1777] = 'h00001318; 
    validation_data[ 1778] = 'h00003007; 
    validation_data[ 1779] = 'h00001fbf; 
    validation_data[ 1780] = 'h000036f0; 
    validation_data[ 1781] = 'h00002f0a; 
    validation_data[ 1782] = 'h000015de; 
    validation_data[ 1783] = 'h000002ec; 
    validation_data[ 1784] = 'h0000365a; 
    validation_data[ 1785] = 'h0000121a; 
    validation_data[ 1786] = 'h00000625; 
    validation_data[ 1787] = 'h000027a9; 
    validation_data[ 1788] = 'h00002fc2; 
    validation_data[ 1789] = 'h00003e94; 
    validation_data[ 1790] = 'h00002ada; 
    validation_data[ 1791] = 'h000036a9; 
    validation_data[ 1792] = 'h0000308c; 
    validation_data[ 1793] = 'h00002e75; 
    validation_data[ 1794] = 'h00000def; 
    validation_data[ 1795] = 'h00003aed; 
    validation_data[ 1796] = 'h0000063e; 
    validation_data[ 1797] = 'h00000e26; 
    validation_data[ 1798] = 'h00002ea1; 
    validation_data[ 1799] = 'h00000f83; 
    validation_data[ 1800] = 'h00000e59; 
    validation_data[ 1801] = 'h000039c3; 
    validation_data[ 1802] = 'h00002385; 
    validation_data[ 1803] = 'h00003f65; 
    validation_data[ 1804] = 'h00000f00; 
    validation_data[ 1805] = 'h00002bcb; 
    validation_data[ 1806] = 'h00002e80; 
    validation_data[ 1807] = 'h000015e1; 
    validation_data[ 1808] = 'h000034bb; 
    validation_data[ 1809] = 'h00000ee1; 
    validation_data[ 1810] = 'h00003a13; 
    validation_data[ 1811] = 'h00002cf4; 
    validation_data[ 1812] = 'h00001dcc; 
    validation_data[ 1813] = 'h00003afd; 
    validation_data[ 1814] = 'h00001638; 
    validation_data[ 1815] = 'h00003556; 
    validation_data[ 1816] = 'h00003ca1; 
    validation_data[ 1817] = 'h0000367c; 
    validation_data[ 1818] = 'h00002b44; 
    validation_data[ 1819] = 'h00002c70; 
    validation_data[ 1820] = 'h00001f73; 
    validation_data[ 1821] = 'h00000dda; 
    validation_data[ 1822] = 'h00001088; 
    validation_data[ 1823] = 'h00000441; 
    validation_data[ 1824] = 'h00002d9d; 
    validation_data[ 1825] = 'h000003be; 
    validation_data[ 1826] = 'h00000b6c; 
    validation_data[ 1827] = 'h00000b79; 
    validation_data[ 1828] = 'h000015f7; 
    validation_data[ 1829] = 'h00001d23; 
    validation_data[ 1830] = 'h00001a8b; 
    validation_data[ 1831] = 'h00001d46; 
    validation_data[ 1832] = 'h00002684; 
    validation_data[ 1833] = 'h00003882; 
    validation_data[ 1834] = 'h000036af; 
    validation_data[ 1835] = 'h00001dd1; 
    validation_data[ 1836] = 'h00001131; 
    validation_data[ 1837] = 'h0000213b; 
    validation_data[ 1838] = 'h00001baf; 
    validation_data[ 1839] = 'h00000b54; 
    validation_data[ 1840] = 'h00001243; 
    validation_data[ 1841] = 'h00001ca9; 
    validation_data[ 1842] = 'h00001b41; 
    validation_data[ 1843] = 'h00001536; 
    validation_data[ 1844] = 'h00001638; 
    validation_data[ 1845] = 'h00000a5a; 
    validation_data[ 1846] = 'h00003b26; 
    validation_data[ 1847] = 'h00002244; 
    validation_data[ 1848] = 'h00000f8c; 
    validation_data[ 1849] = 'h00003544; 
    validation_data[ 1850] = 'h00001572; 
    validation_data[ 1851] = 'h00001c4c; 
    validation_data[ 1852] = 'h00003a79; 
    validation_data[ 1853] = 'h00003859; 
    validation_data[ 1854] = 'h000001f9; 
    validation_data[ 1855] = 'h00000f49; 
    validation_data[ 1856] = 'h000007bb; 
    validation_data[ 1857] = 'h0000163b; 
    validation_data[ 1858] = 'h00002e64; 
    validation_data[ 1859] = 'h000020a9; 
    validation_data[ 1860] = 'h00002616; 
    validation_data[ 1861] = 'h00003678; 
    validation_data[ 1862] = 'h00002df1; 
    validation_data[ 1863] = 'h00000942; 
    validation_data[ 1864] = 'h00001abd; 
    validation_data[ 1865] = 'h000029e7; 
    validation_data[ 1866] = 'h00001b85; 
    validation_data[ 1867] = 'h00000ff4; 
    validation_data[ 1868] = 'h000018f6; 
    validation_data[ 1869] = 'h00002ee6; 
    validation_data[ 1870] = 'h00000fcb; 
    validation_data[ 1871] = 'h00002912; 
    validation_data[ 1872] = 'h00003388; 
    validation_data[ 1873] = 'h000009c4; 
    validation_data[ 1874] = 'h00002ba9; 
    validation_data[ 1875] = 'h0000347e; 
    validation_data[ 1876] = 'h0000364c; 
    validation_data[ 1877] = 'h000010d3; 
    validation_data[ 1878] = 'h00000eb7; 
    validation_data[ 1879] = 'h00001b9c; 
    validation_data[ 1880] = 'h00003883; 
    validation_data[ 1881] = 'h0000139c; 
    validation_data[ 1882] = 'h00003eae; 
    validation_data[ 1883] = 'h00002251; 
    validation_data[ 1884] = 'h000020b8; 
    validation_data[ 1885] = 'h000022bc; 
    validation_data[ 1886] = 'h00001219; 
    validation_data[ 1887] = 'h00003cc8; 
    validation_data[ 1888] = 'h000032d0; 
    validation_data[ 1889] = 'h00001677; 
    validation_data[ 1890] = 'h000021fd; 
    validation_data[ 1891] = 'h0000253d; 
    validation_data[ 1892] = 'h000012b0; 
    validation_data[ 1893] = 'h00001957; 
    validation_data[ 1894] = 'h00000932; 
    validation_data[ 1895] = 'h00003c9f; 
    validation_data[ 1896] = 'h00000fc9; 
    validation_data[ 1897] = 'h00001121; 
    validation_data[ 1898] = 'h00000234; 
    validation_data[ 1899] = 'h00000824; 
    validation_data[ 1900] = 'h000036c9; 
    validation_data[ 1901] = 'h00001f0c; 
    validation_data[ 1902] = 'h0000349b; 
    validation_data[ 1903] = 'h00003aab; 
    validation_data[ 1904] = 'h00003ba6; 
    validation_data[ 1905] = 'h00002ff9; 
    validation_data[ 1906] = 'h00001314; 
    validation_data[ 1907] = 'h00003b4c; 
    validation_data[ 1908] = 'h00001340; 
    validation_data[ 1909] = 'h00003028; 
    validation_data[ 1910] = 'h00000cd7; 
    validation_data[ 1911] = 'h00000acd; 
    validation_data[ 1912] = 'h00001ca4; 
    validation_data[ 1913] = 'h00001b0d; 
    validation_data[ 1914] = 'h00000881; 
    validation_data[ 1915] = 'h000026c3; 
    validation_data[ 1916] = 'h00003a19; 
    validation_data[ 1917] = 'h00003329; 
    validation_data[ 1918] = 'h0000385f; 
    validation_data[ 1919] = 'h00001523; 
    validation_data[ 1920] = 'h00002963; 
    validation_data[ 1921] = 'h00000ee0; 
    validation_data[ 1922] = 'h00000791; 
    validation_data[ 1923] = 'h00003ebf; 
    validation_data[ 1924] = 'h00000bef; 
    validation_data[ 1925] = 'h00000436; 
    validation_data[ 1926] = 'h00003a7f; 
    validation_data[ 1927] = 'h00001b27; 
    validation_data[ 1928] = 'h000018fc; 
    validation_data[ 1929] = 'h00003369; 
    validation_data[ 1930] = 'h0000092d; 
    validation_data[ 1931] = 'h0000315a; 
    validation_data[ 1932] = 'h00000d37; 
    validation_data[ 1933] = 'h00001a85; 
    validation_data[ 1934] = 'h000036c2; 
    validation_data[ 1935] = 'h00001ab8; 
    validation_data[ 1936] = 'h00001157; 
    validation_data[ 1937] = 'h00003157; 
    validation_data[ 1938] = 'h00003f8e; 
    validation_data[ 1939] = 'h000017fe; 
    validation_data[ 1940] = 'h00003d25; 
    validation_data[ 1941] = 'h00001dad; 
    validation_data[ 1942] = 'h000021ef; 
    validation_data[ 1943] = 'h00002c66; 
    validation_data[ 1944] = 'h00003882; 
    validation_data[ 1945] = 'h00000453; 
    validation_data[ 1946] = 'h00003075; 
    validation_data[ 1947] = 'h00000d3f; 
    validation_data[ 1948] = 'h00001d4e; 
    validation_data[ 1949] = 'h00001f55; 
    validation_data[ 1950] = 'h00000ec0; 
    validation_data[ 1951] = 'h00002535; 
    validation_data[ 1952] = 'h000037d8; 
    validation_data[ 1953] = 'h00003cb0; 
    validation_data[ 1954] = 'h0000094a; 
    validation_data[ 1955] = 'h0000283b; 
    validation_data[ 1956] = 'h00001d4d; 
    validation_data[ 1957] = 'h00000170; 
    validation_data[ 1958] = 'h00001848; 
    validation_data[ 1959] = 'h00003c6f; 
    validation_data[ 1960] = 'h00003804; 
    validation_data[ 1961] = 'h00003b64; 
    validation_data[ 1962] = 'h000019ea; 
    validation_data[ 1963] = 'h000019da; 
    validation_data[ 1964] = 'h000006e7; 
    validation_data[ 1965] = 'h00000eec; 
    validation_data[ 1966] = 'h00001995; 
    validation_data[ 1967] = 'h000032ab; 
    validation_data[ 1968] = 'h000022ea; 
    validation_data[ 1969] = 'h000016c9; 
    validation_data[ 1970] = 'h00001e48; 
    validation_data[ 1971] = 'h0000346d; 
    validation_data[ 1972] = 'h000021d8; 
    validation_data[ 1973] = 'h00001b44; 
    validation_data[ 1974] = 'h000038ae; 
    validation_data[ 1975] = 'h00002d6a; 
    validation_data[ 1976] = 'h000030ef; 
    validation_data[ 1977] = 'h0000032f; 
    validation_data[ 1978] = 'h000002d5; 
    validation_data[ 1979] = 'h00002cb3; 
    validation_data[ 1980] = 'h000036fb; 
    validation_data[ 1981] = 'h000009fb; 
    validation_data[ 1982] = 'h000006ff; 
    validation_data[ 1983] = 'h00000c26; 
    validation_data[ 1984] = 'h0000212c; 
    validation_data[ 1985] = 'h000035d2; 
    validation_data[ 1986] = 'h0000000d; 
    validation_data[ 1987] = 'h00003d02; 
    validation_data[ 1988] = 'h000007b6; 
    validation_data[ 1989] = 'h00003fdd; 
    validation_data[ 1990] = 'h00001de6; 
    validation_data[ 1991] = 'h00000faa; 
    validation_data[ 1992] = 'h00002cb2; 
    validation_data[ 1993] = 'h00002b28; 
    validation_data[ 1994] = 'h0000232d; 
    validation_data[ 1995] = 'h0000372a; 
    validation_data[ 1996] = 'h0000127f; 
    validation_data[ 1997] = 'h00002aa0; 
    validation_data[ 1998] = 'h00000631; 
    validation_data[ 1999] = 'h00003296; 
    validation_data[ 2000] = 'h000035cb; 
    validation_data[ 2001] = 'h00001734; 
    validation_data[ 2002] = 'h00003f74; 
    validation_data[ 2003] = 'h000034dc; 
    validation_data[ 2004] = 'h00003060; 
    validation_data[ 2005] = 'h00002d1d; 
    validation_data[ 2006] = 'h0000330d; 
    validation_data[ 2007] = 'h00001236; 
    validation_data[ 2008] = 'h00003ef9; 
    validation_data[ 2009] = 'h00001dde; 
    validation_data[ 2010] = 'h000017f0; 
    validation_data[ 2011] = 'h00003961; 
    validation_data[ 2012] = 'h00002923; 
    validation_data[ 2013] = 'h00003e6b; 
    validation_data[ 2014] = 'h000030a0; 
    validation_data[ 2015] = 'h0000087f; 
    validation_data[ 2016] = 'h000033a9; 
    validation_data[ 2017] = 'h00000789; 
    validation_data[ 2018] = 'h00000441; 
    validation_data[ 2019] = 'h00001d9d; 
    validation_data[ 2020] = 'h00002511; 
    validation_data[ 2021] = 'h00002b77; 
    validation_data[ 2022] = 'h000023e1; 
    validation_data[ 2023] = 'h00002757; 
    validation_data[ 2024] = 'h000010d5; 
    validation_data[ 2025] = 'h00000595; 
    validation_data[ 2026] = 'h00003295; 
    validation_data[ 2027] = 'h0000025d; 
    validation_data[ 2028] = 'h0000037f; 
    validation_data[ 2029] = 'h00002bab; 
    validation_data[ 2030] = 'h000036a5; 
    validation_data[ 2031] = 'h00001411; 
    validation_data[ 2032] = 'h00001cdc; 
    validation_data[ 2033] = 'h000038be; 
    validation_data[ 2034] = 'h000030d9; 
    validation_data[ 2035] = 'h00002a4f; 
    validation_data[ 2036] = 'h000000f9; 
    validation_data[ 2037] = 'h000028bc; 
    validation_data[ 2038] = 'h000009df; 
    validation_data[ 2039] = 'h00000f05; 
    validation_data[ 2040] = 'h00000746; 
    validation_data[ 2041] = 'h00002b23; 
    validation_data[ 2042] = 'h00003442; 
    validation_data[ 2043] = 'h0000307e; 
    validation_data[ 2044] = 'h0000011b; 
    validation_data[ 2045] = 'h00003e62; 
    validation_data[ 2046] = 'h00001981; 
    validation_data[ 2047] = 'h000004dc; 
    validation_data[ 2048] = 'h00001858; 
    validation_data[ 2049] = 'h000015a4; 
    validation_data[ 2050] = 'h00002d00; 
    validation_data[ 2051] = 'h00003afc; 
    validation_data[ 2052] = 'h000030e3; 
    validation_data[ 2053] = 'h0000207b; 
    validation_data[ 2054] = 'h00001337; 
    validation_data[ 2055] = 'h000024f9; 
    validation_data[ 2056] = 'h00000fde; 
    validation_data[ 2057] = 'h00003e84; 
    validation_data[ 2058] = 'h0000202c; 
    validation_data[ 2059] = 'h00002494; 
    validation_data[ 2060] = 'h00001e2b; 
    validation_data[ 2061] = 'h00003a9a; 
    validation_data[ 2062] = 'h000002c1; 
    validation_data[ 2063] = 'h00000f98; 
    validation_data[ 2064] = 'h00001b62; 
    validation_data[ 2065] = 'h00003b15; 
    validation_data[ 2066] = 'h00001c35; 
    validation_data[ 2067] = 'h000031f8; 
    validation_data[ 2068] = 'h00002a0f; 
    validation_data[ 2069] = 'h00000708; 
    validation_data[ 2070] = 'h00000623; 
    validation_data[ 2071] = 'h00000488; 
    validation_data[ 2072] = 'h0000192e; 
    validation_data[ 2073] = 'h00002dd6; 
    validation_data[ 2074] = 'h00000209; 
    validation_data[ 2075] = 'h00003b59; 
    validation_data[ 2076] = 'h00001857; 
    validation_data[ 2077] = 'h0000100e; 
    validation_data[ 2078] = 'h00003eff; 
    validation_data[ 2079] = 'h00000e11; 
    validation_data[ 2080] = 'h000017f7; 
    validation_data[ 2081] = 'h00000e58; 
    validation_data[ 2082] = 'h00000649; 
    validation_data[ 2083] = 'h00002c33; 
    validation_data[ 2084] = 'h000029b4; 
    validation_data[ 2085] = 'h00003b2c; 
    validation_data[ 2086] = 'h000031e6; 
    validation_data[ 2087] = 'h00002851; 
    validation_data[ 2088] = 'h000038d5; 
    validation_data[ 2089] = 'h000038e1; 
    validation_data[ 2090] = 'h00001254; 
    validation_data[ 2091] = 'h0000261b; 
    validation_data[ 2092] = 'h00002c28; 
    validation_data[ 2093] = 'h00000233; 
    validation_data[ 2094] = 'h00000067; 
    validation_data[ 2095] = 'h00001927; 
    validation_data[ 2096] = 'h00000874; 
    validation_data[ 2097] = 'h00003969; 
    validation_data[ 2098] = 'h00000688; 
    validation_data[ 2099] = 'h0000156c; 
    validation_data[ 2100] = 'h00002993; 
    validation_data[ 2101] = 'h00002c53; 
    validation_data[ 2102] = 'h00000ec1; 
    validation_data[ 2103] = 'h00000602; 
    validation_data[ 2104] = 'h00000dce; 
    validation_data[ 2105] = 'h0000305f; 
    validation_data[ 2106] = 'h00003a3d; 
    validation_data[ 2107] = 'h00003aea; 
    validation_data[ 2108] = 'h00000fe5; 
    validation_data[ 2109] = 'h0000130f; 
    validation_data[ 2110] = 'h00001c6b; 
    validation_data[ 2111] = 'h00002d8a; 
    validation_data[ 2112] = 'h00001d8b; 
    validation_data[ 2113] = 'h00001616; 
    validation_data[ 2114] = 'h0000397b; 
    validation_data[ 2115] = 'h00002b05; 
    validation_data[ 2116] = 'h000023ca; 
    validation_data[ 2117] = 'h0000366f; 
    validation_data[ 2118] = 'h00001c91; 
    validation_data[ 2119] = 'h000019ac; 
    validation_data[ 2120] = 'h0000014f; 
    validation_data[ 2121] = 'h00001478; 
    validation_data[ 2122] = 'h00002d62; 
    validation_data[ 2123] = 'h000027cd; 
    validation_data[ 2124] = 'h00003d37; 
    validation_data[ 2125] = 'h00002e7c; 
    validation_data[ 2126] = 'h00001322; 
    validation_data[ 2127] = 'h00001399; 
    validation_data[ 2128] = 'h00002560; 
    validation_data[ 2129] = 'h00000377; 
    validation_data[ 2130] = 'h00002da8; 
    validation_data[ 2131] = 'h00001adc; 
    validation_data[ 2132] = 'h000013a5; 
    validation_data[ 2133] = 'h000023b0; 
    validation_data[ 2134] = 'h00000271; 
    validation_data[ 2135] = 'h00001d75; 
    validation_data[ 2136] = 'h00003777; 
    validation_data[ 2137] = 'h0000325d; 
    validation_data[ 2138] = 'h00002c20; 
    validation_data[ 2139] = 'h000017b9; 
    validation_data[ 2140] = 'h000022b7; 
    validation_data[ 2141] = 'h000004a6; 
    validation_data[ 2142] = 'h0000039d; 
    validation_data[ 2143] = 'h00001e01; 
    validation_data[ 2144] = 'h00002f44; 
    validation_data[ 2145] = 'h00001ce0; 
    validation_data[ 2146] = 'h000002e3; 
    validation_data[ 2147] = 'h000014d0; 
    validation_data[ 2148] = 'h000021b2; 
    validation_data[ 2149] = 'h00003320; 
    validation_data[ 2150] = 'h000013e7; 
    validation_data[ 2151] = 'h00003ec6; 
    validation_data[ 2152] = 'h00001f35; 
    validation_data[ 2153] = 'h00001685; 
    validation_data[ 2154] = 'h000017e7; 
    validation_data[ 2155] = 'h00003595; 
    validation_data[ 2156] = 'h00000f8b; 
    validation_data[ 2157] = 'h000031ad; 
    validation_data[ 2158] = 'h00003d3a; 
    validation_data[ 2159] = 'h00002d20; 
    validation_data[ 2160] = 'h0000231d; 
    validation_data[ 2161] = 'h00003b22; 
    validation_data[ 2162] = 'h0000291d; 
    validation_data[ 2163] = 'h00001d6c; 
    validation_data[ 2164] = 'h0000276a; 
    validation_data[ 2165] = 'h000008ae; 
    validation_data[ 2166] = 'h00000c37; 
    validation_data[ 2167] = 'h00000bee; 
    validation_data[ 2168] = 'h0000130c; 
    validation_data[ 2169] = 'h00001552; 
    validation_data[ 2170] = 'h00000584; 
    validation_data[ 2171] = 'h0000193e; 
    validation_data[ 2172] = 'h0000108e; 
    validation_data[ 2173] = 'h000013f8; 
    validation_data[ 2174] = 'h00001f6f; 
    validation_data[ 2175] = 'h000032fb; 
    validation_data[ 2176] = 'h000000b2; 
    validation_data[ 2177] = 'h00000827; 
    validation_data[ 2178] = 'h00000a98; 
    validation_data[ 2179] = 'h00002bfe; 
    validation_data[ 2180] = 'h0000037a; 
    validation_data[ 2181] = 'h00000fb5; 
    validation_data[ 2182] = 'h000035e0; 
    validation_data[ 2183] = 'h00002878; 
    validation_data[ 2184] = 'h00003a6f; 
    validation_data[ 2185] = 'h00002acb; 
    validation_data[ 2186] = 'h00000b3a; 
    validation_data[ 2187] = 'h0000048d; 
    validation_data[ 2188] = 'h000039b9; 
    validation_data[ 2189] = 'h00001f5e; 
    validation_data[ 2190] = 'h000015e4; 
    validation_data[ 2191] = 'h000019de; 
    validation_data[ 2192] = 'h000012ad; 
    validation_data[ 2193] = 'h000025a5; 
    validation_data[ 2194] = 'h00002797; 
    validation_data[ 2195] = 'h00003a48; 
    validation_data[ 2196] = 'h00003883; 
    validation_data[ 2197] = 'h00000159; 
    validation_data[ 2198] = 'h00003acb; 
    validation_data[ 2199] = 'h00003cab; 
    validation_data[ 2200] = 'h0000349e; 
    validation_data[ 2201] = 'h00001647; 
    validation_data[ 2202] = 'h0000335d; 
    validation_data[ 2203] = 'h00001859; 
    validation_data[ 2204] = 'h00000163; 
    validation_data[ 2205] = 'h00001b38; 
    validation_data[ 2206] = 'h0000224b; 
    validation_data[ 2207] = 'h0000091e; 
    validation_data[ 2208] = 'h000019a8; 
    validation_data[ 2209] = 'h00003ec5; 
    validation_data[ 2210] = 'h00003897; 
    validation_data[ 2211] = 'h00000d24; 
    validation_data[ 2212] = 'h00000bd9; 
    validation_data[ 2213] = 'h00000a36; 
    validation_data[ 2214] = 'h00001e16; 
    validation_data[ 2215] = 'h00003d55; 
    validation_data[ 2216] = 'h000017b1; 
    validation_data[ 2217] = 'h0000221d; 
    validation_data[ 2218] = 'h000000b0; 
    validation_data[ 2219] = 'h00003fd4; 
    validation_data[ 2220] = 'h000037f7; 
    validation_data[ 2221] = 'h00003c4e; 
    validation_data[ 2222] = 'h00002943; 
    validation_data[ 2223] = 'h000021ec; 
    validation_data[ 2224] = 'h00003571; 
    validation_data[ 2225] = 'h000020ac; 
    validation_data[ 2226] = 'h00002e80; 
    validation_data[ 2227] = 'h00000ec4; 
    validation_data[ 2228] = 'h0000065c; 
    validation_data[ 2229] = 'h00001fcf; 
    validation_data[ 2230] = 'h00000032; 
    validation_data[ 2231] = 'h0000309d; 
    validation_data[ 2232] = 'h00003f46; 
    validation_data[ 2233] = 'h00002495; 
    validation_data[ 2234] = 'h00000c8f; 
    validation_data[ 2235] = 'h000027b2; 
    validation_data[ 2236] = 'h0000238f; 
    validation_data[ 2237] = 'h00000597; 
    validation_data[ 2238] = 'h00000f54; 
    validation_data[ 2239] = 'h00000e85; 
    validation_data[ 2240] = 'h00003bbc; 
    validation_data[ 2241] = 'h0000116f; 
    validation_data[ 2242] = 'h00002bf9; 
    validation_data[ 2243] = 'h000001dd; 
    validation_data[ 2244] = 'h00003333; 
    validation_data[ 2245] = 'h00003440; 
    validation_data[ 2246] = 'h000016e9; 
    validation_data[ 2247] = 'h00001251; 
    validation_data[ 2248] = 'h000000f7; 
    validation_data[ 2249] = 'h00003642; 
    validation_data[ 2250] = 'h000018a1; 
    validation_data[ 2251] = 'h00003604; 
    validation_data[ 2252] = 'h000011d9; 
    validation_data[ 2253] = 'h000031a3; 
    validation_data[ 2254] = 'h00001dda; 
    validation_data[ 2255] = 'h000037b1; 
    validation_data[ 2256] = 'h00000d48; 
    validation_data[ 2257] = 'h0000381b; 
    validation_data[ 2258] = 'h00003689; 
    validation_data[ 2259] = 'h00003059; 
    validation_data[ 2260] = 'h000000a9; 
    validation_data[ 2261] = 'h00001c5f; 
    validation_data[ 2262] = 'h0000327a; 
    validation_data[ 2263] = 'h0000064f; 
    validation_data[ 2264] = 'h00003574; 
    validation_data[ 2265] = 'h000021f5; 
    validation_data[ 2266] = 'h0000372d; 
    validation_data[ 2267] = 'h00003cf9; 
    validation_data[ 2268] = 'h00000464; 
    validation_data[ 2269] = 'h0000190c; 
    validation_data[ 2270] = 'h00000235; 
    validation_data[ 2271] = 'h0000260d; 
    validation_data[ 2272] = 'h00001254; 
    validation_data[ 2273] = 'h00000991; 
    validation_data[ 2274] = 'h0000268d; 
    validation_data[ 2275] = 'h000029b9; 
    validation_data[ 2276] = 'h000034aa; 
    validation_data[ 2277] = 'h000030f7; 
    validation_data[ 2278] = 'h000000a3; 
    validation_data[ 2279] = 'h0000030d; 
    validation_data[ 2280] = 'h00003a99; 
    validation_data[ 2281] = 'h00003156; 
    validation_data[ 2282] = 'h000015e9; 
    validation_data[ 2283] = 'h00003b4f; 
    validation_data[ 2284] = 'h00002626; 
    validation_data[ 2285] = 'h000020a5; 
    validation_data[ 2286] = 'h000036be; 
    validation_data[ 2287] = 'h00003266; 
    validation_data[ 2288] = 'h00003145; 
    validation_data[ 2289] = 'h0000241a; 
    validation_data[ 2290] = 'h00000c06; 
    validation_data[ 2291] = 'h000030da; 
    validation_data[ 2292] = 'h00003b0e; 
    validation_data[ 2293] = 'h00003f8e; 
    validation_data[ 2294] = 'h00001fa5; 
    validation_data[ 2295] = 'h00001133; 
    validation_data[ 2296] = 'h00003d93; 
    validation_data[ 2297] = 'h00003bcb; 
    validation_data[ 2298] = 'h00002047; 
    validation_data[ 2299] = 'h00001115; 
    validation_data[ 2300] = 'h00001e57; 
    validation_data[ 2301] = 'h00002d32; 
    validation_data[ 2302] = 'h00001fd7; 
    validation_data[ 2303] = 'h00001228; 
    validation_data[ 2304] = 'h00000d16; 
    validation_data[ 2305] = 'h0000282c; 
    validation_data[ 2306] = 'h000009c4; 
    validation_data[ 2307] = 'h0000277a; 
    validation_data[ 2308] = 'h00003ee2; 
    validation_data[ 2309] = 'h000003fe; 
    validation_data[ 2310] = 'h00002991; 
    validation_data[ 2311] = 'h0000129f; 
    validation_data[ 2312] = 'h00003bc2; 
    validation_data[ 2313] = 'h000011de; 
    validation_data[ 2314] = 'h00000a05; 
    validation_data[ 2315] = 'h00000638; 
    validation_data[ 2316] = 'h000035d3; 
    validation_data[ 2317] = 'h000034cc; 
    validation_data[ 2318] = 'h00001cee; 
    validation_data[ 2319] = 'h00000dc8; 
    validation_data[ 2320] = 'h000035b5; 
    validation_data[ 2321] = 'h0000144a; 
    validation_data[ 2322] = 'h0000157a; 
    validation_data[ 2323] = 'h00003e98; 
    validation_data[ 2324] = 'h000031ba; 
    validation_data[ 2325] = 'h0000229c; 
    validation_data[ 2326] = 'h00002420; 
    validation_data[ 2327] = 'h00002051; 
    validation_data[ 2328] = 'h000005bf; 
    validation_data[ 2329] = 'h00001a7c; 
    validation_data[ 2330] = 'h00002a55; 
    validation_data[ 2331] = 'h0000399b; 
    validation_data[ 2332] = 'h00000976; 
    validation_data[ 2333] = 'h00001417; 
    validation_data[ 2334] = 'h00001b83; 
    validation_data[ 2335] = 'h0000365d; 
    validation_data[ 2336] = 'h00000083; 
    validation_data[ 2337] = 'h00002b0b; 
    validation_data[ 2338] = 'h0000216b; 
    validation_data[ 2339] = 'h00002e2f; 
    validation_data[ 2340] = 'h00000796; 
    validation_data[ 2341] = 'h000029ad; 
    validation_data[ 2342] = 'h00003ddf; 
    validation_data[ 2343] = 'h00002b71; 
    validation_data[ 2344] = 'h0000217e; 
    validation_data[ 2345] = 'h00003d9e; 
    validation_data[ 2346] = 'h000032f4; 
    validation_data[ 2347] = 'h00000a9d; 
    validation_data[ 2348] = 'h000016e9; 
    validation_data[ 2349] = 'h00002bc8; 
    validation_data[ 2350] = 'h00000188; 
    validation_data[ 2351] = 'h00000714; 
    validation_data[ 2352] = 'h000039f8; 
    validation_data[ 2353] = 'h00000ec0; 
    validation_data[ 2354] = 'h0000371b; 
    validation_data[ 2355] = 'h0000050e; 
    validation_data[ 2356] = 'h00000557; 
    validation_data[ 2357] = 'h000009c8; 
    validation_data[ 2358] = 'h00003a1e; 
    validation_data[ 2359] = 'h000026a5; 
    validation_data[ 2360] = 'h00002605; 
    validation_data[ 2361] = 'h000020d6; 
    validation_data[ 2362] = 'h0000066d; 
    validation_data[ 2363] = 'h000027b0; 
    validation_data[ 2364] = 'h0000110d; 
    validation_data[ 2365] = 'h000005fc; 
    validation_data[ 2366] = 'h00002968; 
    validation_data[ 2367] = 'h000038c6; 
    validation_data[ 2368] = 'h00001a91; 
    validation_data[ 2369] = 'h000016f7; 
    validation_data[ 2370] = 'h00000d42; 
    validation_data[ 2371] = 'h00000625; 
    validation_data[ 2372] = 'h00000686; 
    validation_data[ 2373] = 'h00001454; 
    validation_data[ 2374] = 'h000017eb; 
    validation_data[ 2375] = 'h00001693; 
    validation_data[ 2376] = 'h00003b9e; 
    validation_data[ 2377] = 'h00003b20; 
    validation_data[ 2378] = 'h00001e56; 
    validation_data[ 2379] = 'h00001461; 
    validation_data[ 2380] = 'h00002046; 
    validation_data[ 2381] = 'h00000aa8; 
    validation_data[ 2382] = 'h0000167f; 
    validation_data[ 2383] = 'h00003fd8; 
    validation_data[ 2384] = 'h00001c82; 
    validation_data[ 2385] = 'h00003d73; 
    validation_data[ 2386] = 'h000023d2; 
    validation_data[ 2387] = 'h000010c7; 
    validation_data[ 2388] = 'h000003d9; 
    validation_data[ 2389] = 'h000021e4; 
    validation_data[ 2390] = 'h00003594; 
    validation_data[ 2391] = 'h00001969; 
    validation_data[ 2392] = 'h00003188; 
    validation_data[ 2393] = 'h00003a2e; 
    validation_data[ 2394] = 'h00003272; 
    validation_data[ 2395] = 'h00002223; 
    validation_data[ 2396] = 'h00000563; 
    validation_data[ 2397] = 'h000036c6; 
    validation_data[ 2398] = 'h00000a9b; 
    validation_data[ 2399] = 'h00000aa9; 
    validation_data[ 2400] = 'h00000d02; 
    validation_data[ 2401] = 'h0000348e; 
    validation_data[ 2402] = 'h00000217; 
    validation_data[ 2403] = 'h00003971; 
    validation_data[ 2404] = 'h00001b32; 
    validation_data[ 2405] = 'h0000349d; 
    validation_data[ 2406] = 'h00003d5a; 
    validation_data[ 2407] = 'h00001187; 
    validation_data[ 2408] = 'h00001538; 
    validation_data[ 2409] = 'h00001bd0; 
    validation_data[ 2410] = 'h00000e11; 
    validation_data[ 2411] = 'h00001604; 
    validation_data[ 2412] = 'h00001be7; 
    validation_data[ 2413] = 'h00002357; 
    validation_data[ 2414] = 'h000011e4; 
    validation_data[ 2415] = 'h00001bea; 
    validation_data[ 2416] = 'h00002400; 
    validation_data[ 2417] = 'h00003c0c; 
    validation_data[ 2418] = 'h0000202e; 
    validation_data[ 2419] = 'h00000dd0; 
    validation_data[ 2420] = 'h00003381; 
    validation_data[ 2421] = 'h00000418; 
    validation_data[ 2422] = 'h000035f7; 
    validation_data[ 2423] = 'h00002b6b; 
    validation_data[ 2424] = 'h000020c8; 
    validation_data[ 2425] = 'h00002db8; 
    validation_data[ 2426] = 'h00002316; 
    validation_data[ 2427] = 'h00001888; 
    validation_data[ 2428] = 'h0000324f; 
    validation_data[ 2429] = 'h000036e8; 
    validation_data[ 2430] = 'h00002fed; 
    validation_data[ 2431] = 'h000036c3; 
    validation_data[ 2432] = 'h0000354b; 
    validation_data[ 2433] = 'h00001e6f; 
    validation_data[ 2434] = 'h00003742; 
    validation_data[ 2435] = 'h00003fb7; 
    validation_data[ 2436] = 'h000038f3; 
    validation_data[ 2437] = 'h000003b7; 
    validation_data[ 2438] = 'h00003b22; 
    validation_data[ 2439] = 'h00001a07; 
    validation_data[ 2440] = 'h0000115a; 
    validation_data[ 2441] = 'h000033a8; 
    validation_data[ 2442] = 'h000022e5; 
    validation_data[ 2443] = 'h00003b13; 
    validation_data[ 2444] = 'h00002142; 
    validation_data[ 2445] = 'h000009d5; 
    validation_data[ 2446] = 'h000006ff; 
    validation_data[ 2447] = 'h000036b4; 
    validation_data[ 2448] = 'h000010f9; 
    validation_data[ 2449] = 'h00000484; 
    validation_data[ 2450] = 'h000038f8; 
    validation_data[ 2451] = 'h00002358; 
    validation_data[ 2452] = 'h00001863; 
    validation_data[ 2453] = 'h0000341d; 
    validation_data[ 2454] = 'h00003200; 
    validation_data[ 2455] = 'h00002a5a; 
    validation_data[ 2456] = 'h0000057a; 
    validation_data[ 2457] = 'h00001b9b; 
    validation_data[ 2458] = 'h0000047c; 
    validation_data[ 2459] = 'h000012e3; 
    validation_data[ 2460] = 'h000015f3; 
    validation_data[ 2461] = 'h00001587; 
    validation_data[ 2462] = 'h00002b6a; 
    validation_data[ 2463] = 'h00000a4b; 
    validation_data[ 2464] = 'h00001ebd; 
    validation_data[ 2465] = 'h00000f91; 
    validation_data[ 2466] = 'h000038b7; 
    validation_data[ 2467] = 'h000001be; 
    validation_data[ 2468] = 'h0000318d; 
    validation_data[ 2469] = 'h0000330f; 
    validation_data[ 2470] = 'h000002cf; 
    validation_data[ 2471] = 'h000012d5; 
    validation_data[ 2472] = 'h00001c95; 
    validation_data[ 2473] = 'h00003096; 
    validation_data[ 2474] = 'h00001ee6; 
    validation_data[ 2475] = 'h0000217a; 
    validation_data[ 2476] = 'h0000018b; 
    validation_data[ 2477] = 'h00000629; 
    validation_data[ 2478] = 'h0000239f; 
    validation_data[ 2479] = 'h00000a01; 
    validation_data[ 2480] = 'h00000edc; 
    validation_data[ 2481] = 'h00001832; 
    validation_data[ 2482] = 'h000006dc; 
    validation_data[ 2483] = 'h000023ff; 
    validation_data[ 2484] = 'h000037e9; 
    validation_data[ 2485] = 'h00003bba; 
    validation_data[ 2486] = 'h0000114d; 
    validation_data[ 2487] = 'h000014b6; 
    validation_data[ 2488] = 'h000010d4; 
    validation_data[ 2489] = 'h00002560; 
    validation_data[ 2490] = 'h00003fc1; 
    validation_data[ 2491] = 'h00000990; 
    validation_data[ 2492] = 'h0000098c; 
    validation_data[ 2493] = 'h000037fd; 
    validation_data[ 2494] = 'h00000615; 
    validation_data[ 2495] = 'h000036aa; 
    validation_data[ 2496] = 'h0000107f; 
    validation_data[ 2497] = 'h00000317; 
    validation_data[ 2498] = 'h00000b02; 
    validation_data[ 2499] = 'h00000167; 
    validation_data[ 2500] = 'h00001c6f; 
    validation_data[ 2501] = 'h000019cb; 
    validation_data[ 2502] = 'h0000318a; 
    validation_data[ 2503] = 'h00000005; 
    validation_data[ 2504] = 'h0000382a; 
    validation_data[ 2505] = 'h00001a73; 
    validation_data[ 2506] = 'h000036e6; 
    validation_data[ 2507] = 'h00002e6c; 
    validation_data[ 2508] = 'h00003610; 
    validation_data[ 2509] = 'h00001f6b; 
    validation_data[ 2510] = 'h00002b1a; 
    validation_data[ 2511] = 'h000021ca; 
    validation_data[ 2512] = 'h00003a70; 
    validation_data[ 2513] = 'h00002933; 
    validation_data[ 2514] = 'h000012ea; 
    validation_data[ 2515] = 'h000016eb; 
    validation_data[ 2516] = 'h00001c82; 
    validation_data[ 2517] = 'h00003808; 
    validation_data[ 2518] = 'h000022ee; 
    validation_data[ 2519] = 'h00001f2d; 
    validation_data[ 2520] = 'h000008b3; 
    validation_data[ 2521] = 'h00003231; 
    validation_data[ 2522] = 'h000023de; 
    validation_data[ 2523] = 'h000034d6; 
    validation_data[ 2524] = 'h00003928; 
    validation_data[ 2525] = 'h000039fe; 
    validation_data[ 2526] = 'h0000053a; 
    validation_data[ 2527] = 'h000021c7; 
    validation_data[ 2528] = 'h0000186c; 
    validation_data[ 2529] = 'h000022d0; 
    validation_data[ 2530] = 'h00003816; 
    validation_data[ 2531] = 'h0000191d; 
    validation_data[ 2532] = 'h00001483; 
    validation_data[ 2533] = 'h000037d9; 
    validation_data[ 2534] = 'h00000a4d; 
    validation_data[ 2535] = 'h00000cfa; 
    validation_data[ 2536] = 'h0000260e; 
    validation_data[ 2537] = 'h00003b8c; 
    validation_data[ 2538] = 'h000032d2; 
    validation_data[ 2539] = 'h000000f8; 
    validation_data[ 2540] = 'h00003f5a; 
    validation_data[ 2541] = 'h0000154a; 
    validation_data[ 2542] = 'h00001e35; 
    validation_data[ 2543] = 'h000017cf; 
    validation_data[ 2544] = 'h0000073f; 
    validation_data[ 2545] = 'h00001756; 
    validation_data[ 2546] = 'h000007ff; 
    validation_data[ 2547] = 'h00001302; 
    validation_data[ 2548] = 'h00003eff; 
    validation_data[ 2549] = 'h000029e1; 
    validation_data[ 2550] = 'h00003416; 
    validation_data[ 2551] = 'h00001bf2; 
    validation_data[ 2552] = 'h000020c6; 
    validation_data[ 2553] = 'h00002967; 
    validation_data[ 2554] = 'h000014f1; 
    validation_data[ 2555] = 'h000038cf; 
    validation_data[ 2556] = 'h00003cb2; 
    validation_data[ 2557] = 'h00003fec; 
    validation_data[ 2558] = 'h00003c8b; 
    validation_data[ 2559] = 'h0000109b; 
    validation_data[ 2560] = 'h00001727; 
    validation_data[ 2561] = 'h000013e9; 
    validation_data[ 2562] = 'h0000052b; 
    validation_data[ 2563] = 'h00001811; 
    validation_data[ 2564] = 'h00001097; 
    validation_data[ 2565] = 'h00001503; 
    validation_data[ 2566] = 'h000011f0; 
    validation_data[ 2567] = 'h000008b0; 
    validation_data[ 2568] = 'h0000310f; 
    validation_data[ 2569] = 'h0000166e; 
    validation_data[ 2570] = 'h00002fbc; 
    validation_data[ 2571] = 'h00002172; 
    validation_data[ 2572] = 'h00000ce1; 
    validation_data[ 2573] = 'h00000e55; 
    validation_data[ 2574] = 'h00002b34; 
    validation_data[ 2575] = 'h000000b6; 
    validation_data[ 2576] = 'h00001056; 
    validation_data[ 2577] = 'h00000133; 
    validation_data[ 2578] = 'h00000e2f; 
    validation_data[ 2579] = 'h00001792; 
    validation_data[ 2580] = 'h00003546; 
    validation_data[ 2581] = 'h00003a8d; 
    validation_data[ 2582] = 'h000018e0; 
    validation_data[ 2583] = 'h00003b86; 
    validation_data[ 2584] = 'h00002f94; 
    validation_data[ 2585] = 'h00003333; 
    validation_data[ 2586] = 'h0000163c; 
    validation_data[ 2587] = 'h000010d6; 
    validation_data[ 2588] = 'h00002781; 
    validation_data[ 2589] = 'h000039a5; 
    validation_data[ 2590] = 'h0000337f; 
    validation_data[ 2591] = 'h000027a3; 
    validation_data[ 2592] = 'h000008f2; 
    validation_data[ 2593] = 'h00003a8c; 
    validation_data[ 2594] = 'h000025af; 
    validation_data[ 2595] = 'h00001d76; 
    validation_data[ 2596] = 'h000023d8; 
    validation_data[ 2597] = 'h0000215b; 
    validation_data[ 2598] = 'h00001a12; 
    validation_data[ 2599] = 'h000036f9; 
    validation_data[ 2600] = 'h00000ea0; 
    validation_data[ 2601] = 'h00001e18; 
    validation_data[ 2602] = 'h000029bb; 
    validation_data[ 2603] = 'h00003ca3; 
    validation_data[ 2604] = 'h00001f70; 
    validation_data[ 2605] = 'h000006de; 
    validation_data[ 2606] = 'h0000349d; 
    validation_data[ 2607] = 'h000009fd; 
    validation_data[ 2608] = 'h00003401; 
    validation_data[ 2609] = 'h000024f0; 
    validation_data[ 2610] = 'h00003f47; 
    validation_data[ 2611] = 'h00003b76; 
    validation_data[ 2612] = 'h000018fe; 
    validation_data[ 2613] = 'h00003d9b; 
    validation_data[ 2614] = 'h000038b7; 
    validation_data[ 2615] = 'h000015a2; 
    validation_data[ 2616] = 'h00001216; 
    validation_data[ 2617] = 'h000033a0; 
    validation_data[ 2618] = 'h00001ed0; 
    validation_data[ 2619] = 'h000019e4; 
    validation_data[ 2620] = 'h0000262c; 
    validation_data[ 2621] = 'h000036c9; 
    validation_data[ 2622] = 'h00003e86; 
    validation_data[ 2623] = 'h00002c8e; 
    validation_data[ 2624] = 'h00003277; 
    validation_data[ 2625] = 'h000036b2; 
    validation_data[ 2626] = 'h00002da6; 
    validation_data[ 2627] = 'h000025ec; 
    validation_data[ 2628] = 'h0000276f; 
    validation_data[ 2629] = 'h00002f91; 
    validation_data[ 2630] = 'h000008b6; 
    validation_data[ 2631] = 'h00001cbf; 
    validation_data[ 2632] = 'h00002381; 
    validation_data[ 2633] = 'h000029cf; 
    validation_data[ 2634] = 'h00000f9d; 
    validation_data[ 2635] = 'h00003ab7; 
    validation_data[ 2636] = 'h00001a8a; 
    validation_data[ 2637] = 'h00003770; 
    validation_data[ 2638] = 'h000029b3; 
    validation_data[ 2639] = 'h00000a3e; 
    validation_data[ 2640] = 'h00003250; 
    validation_data[ 2641] = 'h0000362f; 
    validation_data[ 2642] = 'h00000d7c; 
    validation_data[ 2643] = 'h00003dee; 
    validation_data[ 2644] = 'h000009b8; 
    validation_data[ 2645] = 'h000022c3; 
    validation_data[ 2646] = 'h00002bcd; 
    validation_data[ 2647] = 'h000007f2; 
    validation_data[ 2648] = 'h00000a8a; 
    validation_data[ 2649] = 'h00000454; 
    validation_data[ 2650] = 'h0000310e; 
    validation_data[ 2651] = 'h00001a87; 
    validation_data[ 2652] = 'h00000e61; 
    validation_data[ 2653] = 'h000033de; 
    validation_data[ 2654] = 'h00003fd2; 
    validation_data[ 2655] = 'h00001cff; 
    validation_data[ 2656] = 'h00003bf0; 
    validation_data[ 2657] = 'h0000384f; 
    validation_data[ 2658] = 'h00003997; 
    validation_data[ 2659] = 'h000005a3; 
    validation_data[ 2660] = 'h00002ffb; 
    validation_data[ 2661] = 'h0000317c; 
    validation_data[ 2662] = 'h00002771; 
    validation_data[ 2663] = 'h00002343; 
    validation_data[ 2664] = 'h000016bd; 
    validation_data[ 2665] = 'h00001c89; 
    validation_data[ 2666] = 'h00003b94; 
    validation_data[ 2667] = 'h00003806; 
    validation_data[ 2668] = 'h00001ea6; 
    validation_data[ 2669] = 'h00001b7c; 
    validation_data[ 2670] = 'h00000998; 
    validation_data[ 2671] = 'h0000317d; 
    validation_data[ 2672] = 'h00002b0a; 
    validation_data[ 2673] = 'h00003b68; 
    validation_data[ 2674] = 'h00003389; 
    validation_data[ 2675] = 'h00001c79; 
    validation_data[ 2676] = 'h000033f8; 
    validation_data[ 2677] = 'h00002fef; 
    validation_data[ 2678] = 'h000030fc; 
    validation_data[ 2679] = 'h000028cb; 
    validation_data[ 2680] = 'h0000024a; 
    validation_data[ 2681] = 'h00002a48; 
    validation_data[ 2682] = 'h00003fac; 
    validation_data[ 2683] = 'h00002dad; 
    validation_data[ 2684] = 'h00001077; 
    validation_data[ 2685] = 'h000039bd; 
    validation_data[ 2686] = 'h00002f47; 
    validation_data[ 2687] = 'h00003ba5; 
    validation_data[ 2688] = 'h00000c09; 
    validation_data[ 2689] = 'h00003802; 
    validation_data[ 2690] = 'h000031c2; 
    validation_data[ 2691] = 'h000010e8; 
    validation_data[ 2692] = 'h00001812; 
    validation_data[ 2693] = 'h000002c9; 
    validation_data[ 2694] = 'h00002aab; 
    validation_data[ 2695] = 'h00000d65; 
    validation_data[ 2696] = 'h00002ac6; 
    validation_data[ 2697] = 'h000020f7; 
    validation_data[ 2698] = 'h00001c57; 
    validation_data[ 2699] = 'h000024bb; 
    validation_data[ 2700] = 'h000015d3; 
    validation_data[ 2701] = 'h0000286f; 
    validation_data[ 2702] = 'h0000209b; 
    validation_data[ 2703] = 'h00000698; 
    validation_data[ 2704] = 'h00000a75; 
    validation_data[ 2705] = 'h00001832; 
    validation_data[ 2706] = 'h000000ff; 
    validation_data[ 2707] = 'h000023ff; 
    validation_data[ 2708] = 'h00002ea0; 
    validation_data[ 2709] = 'h000018eb; 
    validation_data[ 2710] = 'h0000013b; 
    validation_data[ 2711] = 'h00003a50; 
    validation_data[ 2712] = 'h000030cb; 
    validation_data[ 2713] = 'h00001bd2; 
    validation_data[ 2714] = 'h000001ae; 
    validation_data[ 2715] = 'h00001673; 
    validation_data[ 2716] = 'h000039bb; 
    validation_data[ 2717] = 'h00001aeb; 
    validation_data[ 2718] = 'h000030e5; 
    validation_data[ 2719] = 'h0000383b; 
    validation_data[ 2720] = 'h00002a0c; 
    validation_data[ 2721] = 'h00003791; 
    validation_data[ 2722] = 'h00000a9e; 
    validation_data[ 2723] = 'h000033af; 
    validation_data[ 2724] = 'h00003a41; 
    validation_data[ 2725] = 'h000007ad; 
    validation_data[ 2726] = 'h00003638; 
    validation_data[ 2727] = 'h00002188; 
    validation_data[ 2728] = 'h0000220d; 
    validation_data[ 2729] = 'h000039a4; 
    validation_data[ 2730] = 'h00001b14; 
    validation_data[ 2731] = 'h00002636; 
    validation_data[ 2732] = 'h0000107f; 
    validation_data[ 2733] = 'h000032e8; 
    validation_data[ 2734] = 'h0000181d; 
    validation_data[ 2735] = 'h00003bb6; 
    validation_data[ 2736] = 'h000024ad; 
    validation_data[ 2737] = 'h0000182a; 
    validation_data[ 2738] = 'h0000245f; 
    validation_data[ 2739] = 'h0000022e; 
    validation_data[ 2740] = 'h0000101b; 
    validation_data[ 2741] = 'h00002974; 
    validation_data[ 2742] = 'h00002d51; 
    validation_data[ 2743] = 'h00002d76; 
    validation_data[ 2744] = 'h00001ab8; 
    validation_data[ 2745] = 'h000022a4; 
    validation_data[ 2746] = 'h00000c2b; 
    validation_data[ 2747] = 'h00000c36; 
    validation_data[ 2748] = 'h00002bb8; 
    validation_data[ 2749] = 'h000012e5; 
    validation_data[ 2750] = 'h0000345f; 
    validation_data[ 2751] = 'h00002447; 
    validation_data[ 2752] = 'h0000364d; 
    validation_data[ 2753] = 'h00000cca; 
    validation_data[ 2754] = 'h00003e8e; 
    validation_data[ 2755] = 'h00001e55; 
    validation_data[ 2756] = 'h000023d9; 
    validation_data[ 2757] = 'h00003ce1; 
    validation_data[ 2758] = 'h00000bda; 
    validation_data[ 2759] = 'h00002b71; 
    validation_data[ 2760] = 'h00002595; 
    validation_data[ 2761] = 'h00001037; 
    validation_data[ 2762] = 'h000018ef; 
    validation_data[ 2763] = 'h000014b0; 
    validation_data[ 2764] = 'h00001565; 
    validation_data[ 2765] = 'h00003b27; 
    validation_data[ 2766] = 'h00002cf5; 
    validation_data[ 2767] = 'h000011f0; 
    validation_data[ 2768] = 'h00002b29; 
    validation_data[ 2769] = 'h00000d72; 
    validation_data[ 2770] = 'h000002c6; 
    validation_data[ 2771] = 'h00001d75; 
    validation_data[ 2772] = 'h00001cf0; 
    validation_data[ 2773] = 'h00001114; 
    validation_data[ 2774] = 'h0000366f; 
    validation_data[ 2775] = 'h000031c3; 
    validation_data[ 2776] = 'h000005c1; 
    validation_data[ 2777] = 'h000007d4; 
    validation_data[ 2778] = 'h00001238; 
    validation_data[ 2779] = 'h000004a2; 
    validation_data[ 2780] = 'h00001ad0; 
    validation_data[ 2781] = 'h000023b6; 
    validation_data[ 2782] = 'h00000bec; 
    validation_data[ 2783] = 'h00002401; 
    validation_data[ 2784] = 'h00002f6b; 
    validation_data[ 2785] = 'h00002eab; 
    validation_data[ 2786] = 'h0000243f; 
    validation_data[ 2787] = 'h00001dbc; 
    validation_data[ 2788] = 'h00002d0c; 
    validation_data[ 2789] = 'h00002580; 
    validation_data[ 2790] = 'h000001e0; 
    validation_data[ 2791] = 'h000021a5; 
    validation_data[ 2792] = 'h000034a3; 
    validation_data[ 2793] = 'h00001383; 
    validation_data[ 2794] = 'h0000219c; 
    validation_data[ 2795] = 'h000032d4; 
    validation_data[ 2796] = 'h00003b16; 
    validation_data[ 2797] = 'h00002667; 
    validation_data[ 2798] = 'h0000365c; 
    validation_data[ 2799] = 'h00001745; 
    validation_data[ 2800] = 'h00003ef1; 
    validation_data[ 2801] = 'h00002095; 
    validation_data[ 2802] = 'h00002c62; 
    validation_data[ 2803] = 'h0000343c; 
    validation_data[ 2804] = 'h00001fe6; 
    validation_data[ 2805] = 'h00003778; 
    validation_data[ 2806] = 'h00000704; 
    validation_data[ 2807] = 'h0000187e; 
    validation_data[ 2808] = 'h000002f6; 
    validation_data[ 2809] = 'h000025e9; 
    validation_data[ 2810] = 'h000018db; 
    validation_data[ 2811] = 'h00002fd3; 
    validation_data[ 2812] = 'h00003baa; 
    validation_data[ 2813] = 'h00001a90; 
    validation_data[ 2814] = 'h00001a3f; 
    validation_data[ 2815] = 'h00003044; 
    validation_data[ 2816] = 'h00002f31; 
    validation_data[ 2817] = 'h0000223b; 
    validation_data[ 2818] = 'h00000a55; 
    validation_data[ 2819] = 'h00002040; 
    validation_data[ 2820] = 'h0000312f; 
    validation_data[ 2821] = 'h00001b31; 
    validation_data[ 2822] = 'h00003532; 
    validation_data[ 2823] = 'h000024f4; 
    validation_data[ 2824] = 'h00003d65; 
    validation_data[ 2825] = 'h00001a96; 
    validation_data[ 2826] = 'h00003c9f; 
    validation_data[ 2827] = 'h00001b82; 
    validation_data[ 2828] = 'h0000008e; 
    validation_data[ 2829] = 'h00002334; 
    validation_data[ 2830] = 'h00000a6a; 
    validation_data[ 2831] = 'h00000dd9; 
    validation_data[ 2832] = 'h00002df3; 
    validation_data[ 2833] = 'h0000315d; 
    validation_data[ 2834] = 'h0000078b; 
    validation_data[ 2835] = 'h00000b00; 
    validation_data[ 2836] = 'h00000bba; 
    validation_data[ 2837] = 'h000023fb; 
    validation_data[ 2838] = 'h000035bf; 
    validation_data[ 2839] = 'h00003ac4; 
    validation_data[ 2840] = 'h000011b6; 
    validation_data[ 2841] = 'h000014a3; 
    validation_data[ 2842] = 'h000025f9; 
    validation_data[ 2843] = 'h00003ef7; 
    validation_data[ 2844] = 'h000016c0; 
    validation_data[ 2845] = 'h000020f2; 
    validation_data[ 2846] = 'h0000074b; 
    validation_data[ 2847] = 'h0000231d; 
    validation_data[ 2848] = 'h00000196; 
    validation_data[ 2849] = 'h00003acf; 
    validation_data[ 2850] = 'h00003d56; 
    validation_data[ 2851] = 'h0000234b; 
    validation_data[ 2852] = 'h0000002e; 
    validation_data[ 2853] = 'h00002f8f; 
    validation_data[ 2854] = 'h00000ae0; 
    validation_data[ 2855] = 'h00001d20; 
    validation_data[ 2856] = 'h0000395f; 
    validation_data[ 2857] = 'h000025f2; 
    validation_data[ 2858] = 'h00000aa1; 
    validation_data[ 2859] = 'h00002eaf; 
    validation_data[ 2860] = 'h00003a74; 
    validation_data[ 2861] = 'h00000526; 
    validation_data[ 2862] = 'h00001d15; 
    validation_data[ 2863] = 'h000010d3; 
    validation_data[ 2864] = 'h000025fe; 
    validation_data[ 2865] = 'h00001da6; 
    validation_data[ 2866] = 'h000010aa; 
    validation_data[ 2867] = 'h00002b9c; 
    validation_data[ 2868] = 'h0000040d; 
    validation_data[ 2869] = 'h000011ca; 
    validation_data[ 2870] = 'h000006a4; 
    validation_data[ 2871] = 'h000015e1; 
    validation_data[ 2872] = 'h00001939; 
    validation_data[ 2873] = 'h00001a34; 
    validation_data[ 2874] = 'h0000034f; 
    validation_data[ 2875] = 'h000024c8; 
    validation_data[ 2876] = 'h000026d7; 
    validation_data[ 2877] = 'h0000120b; 
    validation_data[ 2878] = 'h0000080e; 
    validation_data[ 2879] = 'h00000ab9; 
    validation_data[ 2880] = 'h0000363f; 
    validation_data[ 2881] = 'h00001a55; 
    validation_data[ 2882] = 'h00000c8b; 
    validation_data[ 2883] = 'h000020e8; 
    validation_data[ 2884] = 'h00000d3b; 
    validation_data[ 2885] = 'h00001f10; 
    validation_data[ 2886] = 'h000039f0; 
    validation_data[ 2887] = 'h000022da; 
    validation_data[ 2888] = 'h000014bf; 
    validation_data[ 2889] = 'h00000215; 
    validation_data[ 2890] = 'h0000025d; 
    validation_data[ 2891] = 'h00000c9e; 
    validation_data[ 2892] = 'h000020ee; 
    validation_data[ 2893] = 'h00002593; 
    validation_data[ 2894] = 'h0000212c; 
    validation_data[ 2895] = 'h000013f4; 
    validation_data[ 2896] = 'h00001193; 
    validation_data[ 2897] = 'h00001f44; 
    validation_data[ 2898] = 'h00003484; 
    validation_data[ 2899] = 'h000014ba; 
    validation_data[ 2900] = 'h00000894; 
    validation_data[ 2901] = 'h00000be8; 
    validation_data[ 2902] = 'h00003d18; 
    validation_data[ 2903] = 'h0000288b; 
    validation_data[ 2904] = 'h00003bc3; 
    validation_data[ 2905] = 'h000039a3; 
    validation_data[ 2906] = 'h0000021e; 
    validation_data[ 2907] = 'h00003265; 
    validation_data[ 2908] = 'h00003066; 
    validation_data[ 2909] = 'h0000351f; 
    validation_data[ 2910] = 'h000024ee; 
    validation_data[ 2911] = 'h00002f3c; 
    validation_data[ 2912] = 'h00003a2e; 
    validation_data[ 2913] = 'h00000a06; 
    validation_data[ 2914] = 'h00001914; 
    validation_data[ 2915] = 'h000018f4; 
    validation_data[ 2916] = 'h000011e9; 
    validation_data[ 2917] = 'h00003c88; 
    validation_data[ 2918] = 'h00000cb7; 
    validation_data[ 2919] = 'h00001a74; 
    validation_data[ 2920] = 'h00001f57; 
    validation_data[ 2921] = 'h000024c4; 
    validation_data[ 2922] = 'h0000358b; 
    validation_data[ 2923] = 'h000024c3; 
    validation_data[ 2924] = 'h00002618; 
    validation_data[ 2925] = 'h00002bc6; 
    validation_data[ 2926] = 'h0000204b; 
    validation_data[ 2927] = 'h00002e40; 
    validation_data[ 2928] = 'h00001587; 
    validation_data[ 2929] = 'h000025d5; 
    validation_data[ 2930] = 'h000008cb; 
    validation_data[ 2931] = 'h00003451; 
    validation_data[ 2932] = 'h00002b35; 
    validation_data[ 2933] = 'h0000329c; 
    validation_data[ 2934] = 'h00001a11; 
    validation_data[ 2935] = 'h00003c5e; 
    validation_data[ 2936] = 'h00001860; 
    validation_data[ 2937] = 'h00001966; 
    validation_data[ 2938] = 'h00001842; 
    validation_data[ 2939] = 'h000035d7; 
    validation_data[ 2940] = 'h00001902; 
    validation_data[ 2941] = 'h0000399c; 
    validation_data[ 2942] = 'h0000207b; 
    validation_data[ 2943] = 'h000029ae; 
    validation_data[ 2944] = 'h00000064; 
    validation_data[ 2945] = 'h00003d6d; 
    validation_data[ 2946] = 'h00002bc6; 
    validation_data[ 2947] = 'h00001710; 
    validation_data[ 2948] = 'h00003ad8; 
    validation_data[ 2949] = 'h000001bb; 
    validation_data[ 2950] = 'h000001a7; 
    validation_data[ 2951] = 'h0000222d; 
    validation_data[ 2952] = 'h000031cb; 
    validation_data[ 2953] = 'h0000255a; 
    validation_data[ 2954] = 'h0000324f; 
    validation_data[ 2955] = 'h00002f30; 
    validation_data[ 2956] = 'h0000098d; 
    validation_data[ 2957] = 'h00003213; 
    validation_data[ 2958] = 'h00001e27; 
    validation_data[ 2959] = 'h00002883; 
    validation_data[ 2960] = 'h00003dd2; 
    validation_data[ 2961] = 'h00003546; 
    validation_data[ 2962] = 'h00001513; 
    validation_data[ 2963] = 'h000035c8; 
    validation_data[ 2964] = 'h00001be3; 
    validation_data[ 2965] = 'h00002f50; 
    validation_data[ 2966] = 'h000015d9; 
    validation_data[ 2967] = 'h00001a1b; 
    validation_data[ 2968] = 'h00003762; 
    validation_data[ 2969] = 'h000009db; 
    validation_data[ 2970] = 'h00001604; 
    validation_data[ 2971] = 'h000011b2; 
    validation_data[ 2972] = 'h000000fc; 
    validation_data[ 2973] = 'h00003559; 
    validation_data[ 2974] = 'h00002815; 
    validation_data[ 2975] = 'h00000e09; 
    validation_data[ 2976] = 'h00001a1d; 
    validation_data[ 2977] = 'h00003248; 
    validation_data[ 2978] = 'h000038ea; 
    validation_data[ 2979] = 'h00002c2d; 
    validation_data[ 2980] = 'h00003f72; 
    validation_data[ 2981] = 'h0000059b; 
    validation_data[ 2982] = 'h00003157; 
    validation_data[ 2983] = 'h00003d30; 
    validation_data[ 2984] = 'h000015ff; 
    validation_data[ 2985] = 'h00003fa9; 
    validation_data[ 2986] = 'h000002b2; 
    validation_data[ 2987] = 'h0000178b; 
    validation_data[ 2988] = 'h000006b8; 
    validation_data[ 2989] = 'h000001af; 
    validation_data[ 2990] = 'h00000475; 
    validation_data[ 2991] = 'h000010db; 
    validation_data[ 2992] = 'h00002874; 
    validation_data[ 2993] = 'h00001b76; 
    validation_data[ 2994] = 'h000012ac; 
    validation_data[ 2995] = 'h00002bde; 
    validation_data[ 2996] = 'h000017fc; 
    validation_data[ 2997] = 'h00001573; 
    validation_data[ 2998] = 'h00002219; 
    validation_data[ 2999] = 'h000009ce; 
    validation_data[ 3000] = 'h00000452; 
    validation_data[ 3001] = 'h0000040b; 
    validation_data[ 3002] = 'h00002b0a; 
    validation_data[ 3003] = 'h00002cbf; 
    validation_data[ 3004] = 'h00001a13; 
    validation_data[ 3005] = 'h000013cf; 
    validation_data[ 3006] = 'h00000674; 
    validation_data[ 3007] = 'h0000227a; 
    validation_data[ 3008] = 'h00001a25; 
    validation_data[ 3009] = 'h00000a00; 
    validation_data[ 3010] = 'h00001a3c; 
    validation_data[ 3011] = 'h000000e3; 
    validation_data[ 3012] = 'h00003d1a; 
    validation_data[ 3013] = 'h00000ef0; 
    validation_data[ 3014] = 'h00003800; 
    validation_data[ 3015] = 'h000020d7; 
    validation_data[ 3016] = 'h00003c39; 
    validation_data[ 3017] = 'h0000016e; 
    validation_data[ 3018] = 'h00003662; 
    validation_data[ 3019] = 'h00000e76; 
    validation_data[ 3020] = 'h00002a17; 
    validation_data[ 3021] = 'h00000271; 
    validation_data[ 3022] = 'h00000386; 
    validation_data[ 3023] = 'h00002a08; 
    validation_data[ 3024] = 'h000017b9; 
    validation_data[ 3025] = 'h000007a0; 
    validation_data[ 3026] = 'h000006f9; 
    validation_data[ 3027] = 'h000006ac; 
    validation_data[ 3028] = 'h00002c38; 
    validation_data[ 3029] = 'h00003531; 
    validation_data[ 3030] = 'h000022e3; 
    validation_data[ 3031] = 'h00002a8d; 
    validation_data[ 3032] = 'h0000377c; 
    validation_data[ 3033] = 'h00000003; 
    validation_data[ 3034] = 'h00002645; 
    validation_data[ 3035] = 'h00002941; 
    validation_data[ 3036] = 'h00002b68; 
    validation_data[ 3037] = 'h00000823; 
    validation_data[ 3038] = 'h00000cc9; 
    validation_data[ 3039] = 'h00002fac; 
    validation_data[ 3040] = 'h00001e2c; 
    validation_data[ 3041] = 'h00001191; 
    validation_data[ 3042] = 'h00003716; 
    validation_data[ 3043] = 'h00001707; 
    validation_data[ 3044] = 'h0000145a; 
    validation_data[ 3045] = 'h00003d3b; 
    validation_data[ 3046] = 'h000027e7; 
    validation_data[ 3047] = 'h00001658; 
    validation_data[ 3048] = 'h000012d4; 
    validation_data[ 3049] = 'h000013e0; 
    validation_data[ 3050] = 'h000017cf; 
    validation_data[ 3051] = 'h00003ca3; 
    validation_data[ 3052] = 'h000026de; 
    validation_data[ 3053] = 'h00002064; 
    validation_data[ 3054] = 'h00001648; 
    validation_data[ 3055] = 'h0000171d; 
    validation_data[ 3056] = 'h000001b2; 
    validation_data[ 3057] = 'h00001069; 
    validation_data[ 3058] = 'h00000f19; 
    validation_data[ 3059] = 'h00000d76; 
    validation_data[ 3060] = 'h00000c92; 
    validation_data[ 3061] = 'h0000070a; 
    validation_data[ 3062] = 'h00000c09; 
    validation_data[ 3063] = 'h00001b88; 
    validation_data[ 3064] = 'h00001844; 
    validation_data[ 3065] = 'h0000221e; 
    validation_data[ 3066] = 'h00000fa5; 
    validation_data[ 3067] = 'h00003d48; 
    validation_data[ 3068] = 'h000000d9; 
    validation_data[ 3069] = 'h00003fe9; 
    validation_data[ 3070] = 'h0000072f; 
    validation_data[ 3071] = 'h000029f6; 
    validation_data[ 3072] = 'h00000eec; 
    validation_data[ 3073] = 'h000011ff; 
    validation_data[ 3074] = 'h000006f9; 
    validation_data[ 3075] = 'h000006a6; 
    validation_data[ 3076] = 'h000017a9; 
    validation_data[ 3077] = 'h00001f7e; 
    validation_data[ 3078] = 'h00003e71; 
    validation_data[ 3079] = 'h00000d01; 
    validation_data[ 3080] = 'h000015dc; 
    validation_data[ 3081] = 'h00002ff4; 
    validation_data[ 3082] = 'h000013be; 
    validation_data[ 3083] = 'h00003465; 
    validation_data[ 3084] = 'h00001349; 
    validation_data[ 3085] = 'h00003d3c; 
    validation_data[ 3086] = 'h00003cb5; 
    validation_data[ 3087] = 'h00000ea0; 
    validation_data[ 3088] = 'h0000226d; 
    validation_data[ 3089] = 'h00002a50; 
    validation_data[ 3090] = 'h000038a7; 
    validation_data[ 3091] = 'h00001070; 
    validation_data[ 3092] = 'h000020d8; 
    validation_data[ 3093] = 'h00000525; 
    validation_data[ 3094] = 'h0000124d; 
    validation_data[ 3095] = 'h00002247; 
    validation_data[ 3096] = 'h000009c4; 
    validation_data[ 3097] = 'h000037d4; 
    validation_data[ 3098] = 'h0000275b; 
    validation_data[ 3099] = 'h00000611; 
    validation_data[ 3100] = 'h00000303; 
    validation_data[ 3101] = 'h000026df; 
    validation_data[ 3102] = 'h00003ea0; 
    validation_data[ 3103] = 'h00002cdf; 
    validation_data[ 3104] = 'h0000000f; 
    validation_data[ 3105] = 'h00000fa8; 
    validation_data[ 3106] = 'h00002ab6; 
    validation_data[ 3107] = 'h00001ae8; 
    validation_data[ 3108] = 'h0000071f; 
    validation_data[ 3109] = 'h000019a0; 
    validation_data[ 3110] = 'h00002df6; 
    validation_data[ 3111] = 'h000028c1; 
    validation_data[ 3112] = 'h000009d0; 
    validation_data[ 3113] = 'h00000b27; 
    validation_data[ 3114] = 'h0000362d; 
    validation_data[ 3115] = 'h000017c7; 
    validation_data[ 3116] = 'h000006a3; 
    validation_data[ 3117] = 'h00002bd7; 
    validation_data[ 3118] = 'h00003481; 
    validation_data[ 3119] = 'h00001702; 
    validation_data[ 3120] = 'h000015fe; 
    validation_data[ 3121] = 'h00001db5; 
    validation_data[ 3122] = 'h00003ea2; 
    validation_data[ 3123] = 'h0000103d; 
    validation_data[ 3124] = 'h000017ad; 
    validation_data[ 3125] = 'h00001cd2; 
    validation_data[ 3126] = 'h00001f4b; 
    validation_data[ 3127] = 'h00000eed; 
    validation_data[ 3128] = 'h000031eb; 
    validation_data[ 3129] = 'h0000287e; 
    validation_data[ 3130] = 'h00000d4e; 
    validation_data[ 3131] = 'h000015ee; 
    validation_data[ 3132] = 'h000006cc; 
    validation_data[ 3133] = 'h00002b5d; 
    validation_data[ 3134] = 'h00000783; 
    validation_data[ 3135] = 'h000013f5; 
    validation_data[ 3136] = 'h0000162b; 
    validation_data[ 3137] = 'h000013f6; 
    validation_data[ 3138] = 'h00000daf; 
    validation_data[ 3139] = 'h00001fa5; 
    validation_data[ 3140] = 'h000017ca; 
    validation_data[ 3141] = 'h00001e4f; 
    validation_data[ 3142] = 'h000015a7; 
    validation_data[ 3143] = 'h00001a57; 
    validation_data[ 3144] = 'h000012fe; 
    validation_data[ 3145] = 'h0000117b; 
    validation_data[ 3146] = 'h00003aae; 
    validation_data[ 3147] = 'h00000e3f; 
    validation_data[ 3148] = 'h00000a83; 
    validation_data[ 3149] = 'h00001622; 
    validation_data[ 3150] = 'h000013d7; 
    validation_data[ 3151] = 'h000018a5; 
    validation_data[ 3152] = 'h00000a56; 
    validation_data[ 3153] = 'h000028e8; 
    validation_data[ 3154] = 'h00003e2a; 
    validation_data[ 3155] = 'h000004e2; 
    validation_data[ 3156] = 'h00002996; 
    validation_data[ 3157] = 'h00002306; 
    validation_data[ 3158] = 'h00003476; 
    validation_data[ 3159] = 'h00002c62; 
    validation_data[ 3160] = 'h000029ca; 
    validation_data[ 3161] = 'h00002008; 
    validation_data[ 3162] = 'h000006f2; 
    validation_data[ 3163] = 'h00000a4b; 
    validation_data[ 3164] = 'h00003ee7; 
    validation_data[ 3165] = 'h00001a3d; 
    validation_data[ 3166] = 'h00001997; 
    validation_data[ 3167] = 'h00002e9f; 
    validation_data[ 3168] = 'h00001370; 
    validation_data[ 3169] = 'h000026ff; 
    validation_data[ 3170] = 'h000012e3; 
    validation_data[ 3171] = 'h000017ef; 
    validation_data[ 3172] = 'h000012c8; 
    validation_data[ 3173] = 'h000035ef; 
    validation_data[ 3174] = 'h00003a61; 
    validation_data[ 3175] = 'h00002550; 
    validation_data[ 3176] = 'h00003271; 
    validation_data[ 3177] = 'h000023d2; 
    validation_data[ 3178] = 'h000039c8; 
    validation_data[ 3179] = 'h000038f3; 
    validation_data[ 3180] = 'h000012bd; 
    validation_data[ 3181] = 'h000016b8; 
    validation_data[ 3182] = 'h000005a5; 
    validation_data[ 3183] = 'h000021e3; 
    validation_data[ 3184] = 'h00003c8e; 
    validation_data[ 3185] = 'h00003151; 
    validation_data[ 3186] = 'h0000214d; 
    validation_data[ 3187] = 'h00001c9d; 
    validation_data[ 3188] = 'h00003f31; 
    validation_data[ 3189] = 'h0000345e; 
    validation_data[ 3190] = 'h000027c7; 
    validation_data[ 3191] = 'h00003883; 
    validation_data[ 3192] = 'h000009a6; 
    validation_data[ 3193] = 'h00001d3d; 
    validation_data[ 3194] = 'h00000f6e; 
    validation_data[ 3195] = 'h00000c9e; 
    validation_data[ 3196] = 'h00000e0d; 
    validation_data[ 3197] = 'h00002c0e; 
    validation_data[ 3198] = 'h0000279f; 
    validation_data[ 3199] = 'h00002232; 
    validation_data[ 3200] = 'h0000296c; 
    validation_data[ 3201] = 'h00001dd8; 
    validation_data[ 3202] = 'h00001c78; 
    validation_data[ 3203] = 'h00003b66; 
    validation_data[ 3204] = 'h00001a87; 
    validation_data[ 3205] = 'h00003a00; 
    validation_data[ 3206] = 'h00000f23; 
    validation_data[ 3207] = 'h00000776; 
    validation_data[ 3208] = 'h00000d6a; 
    validation_data[ 3209] = 'h00000775; 
    validation_data[ 3210] = 'h00000431; 
    validation_data[ 3211] = 'h00001046; 
    validation_data[ 3212] = 'h00003bd7; 
    validation_data[ 3213] = 'h00003c1e; 
    validation_data[ 3214] = 'h00002be9; 
    validation_data[ 3215] = 'h00000203; 
    validation_data[ 3216] = 'h00003a03; 
    validation_data[ 3217] = 'h00002c53; 
    validation_data[ 3218] = 'h00000cba; 
    validation_data[ 3219] = 'h0000146a; 
    validation_data[ 3220] = 'h00003d8d; 
    validation_data[ 3221] = 'h00001091; 
    validation_data[ 3222] = 'h00003302; 
    validation_data[ 3223] = 'h00003941; 
    validation_data[ 3224] = 'h00002818; 
    validation_data[ 3225] = 'h00001aa2; 
    validation_data[ 3226] = 'h000001ec; 
    validation_data[ 3227] = 'h00000e08; 
    validation_data[ 3228] = 'h00003c8f; 
    validation_data[ 3229] = 'h00001dbd; 
    validation_data[ 3230] = 'h0000275f; 
    validation_data[ 3231] = 'h00003b0f; 
    validation_data[ 3232] = 'h00000889; 
    validation_data[ 3233] = 'h000035d6; 
    validation_data[ 3234] = 'h00002484; 
    validation_data[ 3235] = 'h00000370; 
    validation_data[ 3236] = 'h0000266f; 
    validation_data[ 3237] = 'h00003596; 
    validation_data[ 3238] = 'h0000114b; 
    validation_data[ 3239] = 'h000005e8; 
    validation_data[ 3240] = 'h000027fa; 
    validation_data[ 3241] = 'h00002178; 
    validation_data[ 3242] = 'h0000174a; 
    validation_data[ 3243] = 'h000020bd; 
    validation_data[ 3244] = 'h00003cde; 
    validation_data[ 3245] = 'h00000f2d; 
    validation_data[ 3246] = 'h000013d0; 
    validation_data[ 3247] = 'h00000202; 
    validation_data[ 3248] = 'h00002f9f; 
    validation_data[ 3249] = 'h00002040; 
    validation_data[ 3250] = 'h00001ebe; 
    validation_data[ 3251] = 'h00000f19; 
    validation_data[ 3252] = 'h00002a1f; 
    validation_data[ 3253] = 'h0000209d; 
    validation_data[ 3254] = 'h000003a5; 
    validation_data[ 3255] = 'h00003832; 
    validation_data[ 3256] = 'h0000336a; 
    validation_data[ 3257] = 'h000035ed; 
    validation_data[ 3258] = 'h0000352e; 
    validation_data[ 3259] = 'h000034aa; 
    validation_data[ 3260] = 'h000017d7; 
    validation_data[ 3261] = 'h00000bba; 
    validation_data[ 3262] = 'h000000fd; 
    validation_data[ 3263] = 'h00001fe7; 
    validation_data[ 3264] = 'h00002abb; 
    validation_data[ 3265] = 'h0000397c; 
    validation_data[ 3266] = 'h00003177; 
    validation_data[ 3267] = 'h0000165d; 
    validation_data[ 3268] = 'h00001a05; 
    validation_data[ 3269] = 'h00000ddd; 
    validation_data[ 3270] = 'h00002fca; 
    validation_data[ 3271] = 'h00002dd5; 
    validation_data[ 3272] = 'h00002026; 
    validation_data[ 3273] = 'h000009fc; 
    validation_data[ 3274] = 'h000002bc; 
    validation_data[ 3275] = 'h00000e58; 
    validation_data[ 3276] = 'h00000768; 
    validation_data[ 3277] = 'h00001f9b; 
    validation_data[ 3278] = 'h000013aa; 
    validation_data[ 3279] = 'h000012ba; 
    validation_data[ 3280] = 'h000001cd; 
    validation_data[ 3281] = 'h00002caf; 
    validation_data[ 3282] = 'h00003707; 
    validation_data[ 3283] = 'h000037de; 
    validation_data[ 3284] = 'h000026ba; 
    validation_data[ 3285] = 'h000036a8; 
    validation_data[ 3286] = 'h00002b04; 
    validation_data[ 3287] = 'h00002e70; 
    validation_data[ 3288] = 'h000017f1; 
    validation_data[ 3289] = 'h0000389a; 
    validation_data[ 3290] = 'h00001303; 
    validation_data[ 3291] = 'h000030b2; 
    validation_data[ 3292] = 'h00002488; 
    validation_data[ 3293] = 'h0000256e; 
    validation_data[ 3294] = 'h00002a60; 
    validation_data[ 3295] = 'h00003ccd; 
    validation_data[ 3296] = 'h000037b9; 
    validation_data[ 3297] = 'h000032a0; 
    validation_data[ 3298] = 'h00000788; 
    validation_data[ 3299] = 'h000023b5; 
    validation_data[ 3300] = 'h00001b01; 
    validation_data[ 3301] = 'h0000258c; 
    validation_data[ 3302] = 'h00002d94; 
    validation_data[ 3303] = 'h00003d68; 
    validation_data[ 3304] = 'h00001f1a; 
    validation_data[ 3305] = 'h000034f9; 
    validation_data[ 3306] = 'h000023c2; 
    validation_data[ 3307] = 'h00001914; 
    validation_data[ 3308] = 'h000028d4; 
    validation_data[ 3309] = 'h00000f6d; 
    validation_data[ 3310] = 'h00000081; 
    validation_data[ 3311] = 'h00001d04; 
    validation_data[ 3312] = 'h00000cb1; 
    validation_data[ 3313] = 'h000013ff; 
    validation_data[ 3314] = 'h000005e1; 
    validation_data[ 3315] = 'h00002b8b; 
    validation_data[ 3316] = 'h00002acc; 
    validation_data[ 3317] = 'h000003d9; 
    validation_data[ 3318] = 'h00000fb7; 
    validation_data[ 3319] = 'h000003f7; 
    validation_data[ 3320] = 'h00000f6e; 
    validation_data[ 3321] = 'h00000af5; 
    validation_data[ 3322] = 'h00003ea5; 
    validation_data[ 3323] = 'h000020bd; 
    validation_data[ 3324] = 'h00003fbc; 
    validation_data[ 3325] = 'h00002f5a; 
    validation_data[ 3326] = 'h0000094c; 
    validation_data[ 3327] = 'h00000b32; 
    validation_data[ 3328] = 'h00002195; 
    validation_data[ 3329] = 'h0000359c; 
    validation_data[ 3330] = 'h00002a00; 
    validation_data[ 3331] = 'h0000092d; 
    validation_data[ 3332] = 'h00002df8; 
    validation_data[ 3333] = 'h000007d9; 
    validation_data[ 3334] = 'h00003342; 
    validation_data[ 3335] = 'h00002e55; 
    validation_data[ 3336] = 'h00000919; 
    validation_data[ 3337] = 'h00000b7d; 
    validation_data[ 3338] = 'h0000253f; 
    validation_data[ 3339] = 'h00001010; 
    validation_data[ 3340] = 'h00003ef9; 
    validation_data[ 3341] = 'h00003421; 
    validation_data[ 3342] = 'h0000290e; 
    validation_data[ 3343] = 'h0000355d; 
    validation_data[ 3344] = 'h00002cde; 
    validation_data[ 3345] = 'h000027c2; 
    validation_data[ 3346] = 'h00002f21; 
    validation_data[ 3347] = 'h00002c61; 
    validation_data[ 3348] = 'h00001cd9; 
    validation_data[ 3349] = 'h000030b6; 
    validation_data[ 3350] = 'h000026bb; 
    validation_data[ 3351] = 'h00001199; 
    validation_data[ 3352] = 'h0000037a; 
    validation_data[ 3353] = 'h00001abf; 
    validation_data[ 3354] = 'h000001ed; 
    validation_data[ 3355] = 'h00003660; 
    validation_data[ 3356] = 'h00003639; 
    validation_data[ 3357] = 'h00002c4e; 
    validation_data[ 3358] = 'h00001f15; 
    validation_data[ 3359] = 'h0000149f; 
    validation_data[ 3360] = 'h000006cd; 
    validation_data[ 3361] = 'h00000245; 
    validation_data[ 3362] = 'h00002a0c; 
    validation_data[ 3363] = 'h000037be; 
    validation_data[ 3364] = 'h0000134b; 
    validation_data[ 3365] = 'h00000a60; 
    validation_data[ 3366] = 'h00002590; 
    validation_data[ 3367] = 'h000027da; 
    validation_data[ 3368] = 'h0000111e; 
    validation_data[ 3369] = 'h000017f2; 
    validation_data[ 3370] = 'h00001bab; 
    validation_data[ 3371] = 'h00000cb4; 
    validation_data[ 3372] = 'h00001db8; 
    validation_data[ 3373] = 'h00003937; 
    validation_data[ 3374] = 'h00003323; 
    validation_data[ 3375] = 'h00003b9c; 
    validation_data[ 3376] = 'h00001dab; 
    validation_data[ 3377] = 'h00003a8d; 
    validation_data[ 3378] = 'h00001182; 
    validation_data[ 3379] = 'h00001b0e; 
    validation_data[ 3380] = 'h000032f1; 
    validation_data[ 3381] = 'h00002e25; 
    validation_data[ 3382] = 'h00000529; 
    validation_data[ 3383] = 'h00002f5a; 
    validation_data[ 3384] = 'h00000c0a; 
    validation_data[ 3385] = 'h00002bf3; 
    validation_data[ 3386] = 'h00001216; 
    validation_data[ 3387] = 'h000026c5; 
    validation_data[ 3388] = 'h00003320; 
    validation_data[ 3389] = 'h00001dec; 
    validation_data[ 3390] = 'h00002a4c; 
    validation_data[ 3391] = 'h00003868; 
    validation_data[ 3392] = 'h0000274c; 
    validation_data[ 3393] = 'h0000158d; 
    validation_data[ 3394] = 'h00003025; 
    validation_data[ 3395] = 'h00003557; 
    validation_data[ 3396] = 'h00003740; 
    validation_data[ 3397] = 'h000033f0; 
    validation_data[ 3398] = 'h00000b6a; 
    validation_data[ 3399] = 'h000004c6; 
    validation_data[ 3400] = 'h000027d5; 
    validation_data[ 3401] = 'h000005ff; 
    validation_data[ 3402] = 'h00001fb8; 
    validation_data[ 3403] = 'h00001510; 
    validation_data[ 3404] = 'h00003800; 
    validation_data[ 3405] = 'h00002f57; 
    validation_data[ 3406] = 'h00003be2; 
    validation_data[ 3407] = 'h0000303f; 
    validation_data[ 3408] = 'h00003bc2; 
    validation_data[ 3409] = 'h000000fb; 
    validation_data[ 3410] = 'h00000cb7; 
    validation_data[ 3411] = 'h00000bd6; 
    validation_data[ 3412] = 'h00002fe8; 
    validation_data[ 3413] = 'h00003133; 
    validation_data[ 3414] = 'h000013d1; 
    validation_data[ 3415] = 'h00000e89; 
    validation_data[ 3416] = 'h000023ae; 
    validation_data[ 3417] = 'h00000f99; 
    validation_data[ 3418] = 'h000032d4; 
    validation_data[ 3419] = 'h0000239c; 
    validation_data[ 3420] = 'h00002e69; 
    validation_data[ 3421] = 'h00001704; 
    validation_data[ 3422] = 'h00003732; 
    validation_data[ 3423] = 'h00002128; 
    validation_data[ 3424] = 'h00003752; 
    validation_data[ 3425] = 'h00002100; 
    validation_data[ 3426] = 'h00001e3a; 
    validation_data[ 3427] = 'h00000d1a; 
    validation_data[ 3428] = 'h00000662; 
    validation_data[ 3429] = 'h0000185c; 
    validation_data[ 3430] = 'h00000103; 
    validation_data[ 3431] = 'h00001211; 
    validation_data[ 3432] = 'h00000bb4; 
    validation_data[ 3433] = 'h00000cdc; 
    validation_data[ 3434] = 'h000023d9; 
    validation_data[ 3435] = 'h00003cf3; 
    validation_data[ 3436] = 'h000003f5; 
    validation_data[ 3437] = 'h000022b4; 
    validation_data[ 3438] = 'h00001147; 
    validation_data[ 3439] = 'h00001789; 
    validation_data[ 3440] = 'h00002428; 
    validation_data[ 3441] = 'h00001bb0; 
    validation_data[ 3442] = 'h0000236d; 
    validation_data[ 3443] = 'h00000aa5; 
    validation_data[ 3444] = 'h00000788; 
    validation_data[ 3445] = 'h00002f94; 
    validation_data[ 3446] = 'h00000597; 
    validation_data[ 3447] = 'h00001891; 
    validation_data[ 3448] = 'h00002611; 
    validation_data[ 3449] = 'h0000118e; 
    validation_data[ 3450] = 'h00002e6f; 
    validation_data[ 3451] = 'h0000075c; 
    validation_data[ 3452] = 'h0000052b; 
    validation_data[ 3453] = 'h00002ad8; 
    validation_data[ 3454] = 'h00003311; 
    validation_data[ 3455] = 'h00002a67; 
    validation_data[ 3456] = 'h00001b4f; 
    validation_data[ 3457] = 'h0000372f; 
    validation_data[ 3458] = 'h00001c5e; 
    validation_data[ 3459] = 'h00001c7c; 
    validation_data[ 3460] = 'h00002625; 
    validation_data[ 3461] = 'h00000121; 
    validation_data[ 3462] = 'h00001ca5; 
    validation_data[ 3463] = 'h000015cd; 
    validation_data[ 3464] = 'h00001266; 
    validation_data[ 3465] = 'h0000024f; 
    validation_data[ 3466] = 'h00003941; 
    validation_data[ 3467] = 'h00002f1c; 
    validation_data[ 3468] = 'h00000a48; 
    validation_data[ 3469] = 'h000036e8; 
    validation_data[ 3470] = 'h00002f45; 
    validation_data[ 3471] = 'h00001a83; 
    validation_data[ 3472] = 'h0000002b; 
    validation_data[ 3473] = 'h00003677; 
    validation_data[ 3474] = 'h00000ff5; 
    validation_data[ 3475] = 'h0000121e; 
    validation_data[ 3476] = 'h000017b9; 
    validation_data[ 3477] = 'h00000fbd; 
    validation_data[ 3478] = 'h000017de; 
    validation_data[ 3479] = 'h00002eec; 
    validation_data[ 3480] = 'h00000274; 
    validation_data[ 3481] = 'h0000369f; 
    validation_data[ 3482] = 'h00003be0; 
    validation_data[ 3483] = 'h00003019; 
    validation_data[ 3484] = 'h0000071d; 
    validation_data[ 3485] = 'h00001d03; 
    validation_data[ 3486] = 'h00000a3b; 
    validation_data[ 3487] = 'h00001980; 
    validation_data[ 3488] = 'h0000031c; 
    validation_data[ 3489] = 'h00002b54; 
    validation_data[ 3490] = 'h00003f9d; 
    validation_data[ 3491] = 'h000002c1; 
    validation_data[ 3492] = 'h00003db3; 
    validation_data[ 3493] = 'h00002b51; 
    validation_data[ 3494] = 'h00000ce3; 
    validation_data[ 3495] = 'h00001200; 
    validation_data[ 3496] = 'h00000515; 
    validation_data[ 3497] = 'h00003448; 
    validation_data[ 3498] = 'h00003510; 
    validation_data[ 3499] = 'h0000011b; 
    validation_data[ 3500] = 'h00002dd6; 
    validation_data[ 3501] = 'h000010de; 
    validation_data[ 3502] = 'h00002382; 
    validation_data[ 3503] = 'h00003044; 
    validation_data[ 3504] = 'h000005a2; 
    validation_data[ 3505] = 'h00002985; 
    validation_data[ 3506] = 'h00002916; 
    validation_data[ 3507] = 'h000032a3; 
    validation_data[ 3508] = 'h0000194b; 
    validation_data[ 3509] = 'h000008ef; 
    validation_data[ 3510] = 'h000026c4; 
    validation_data[ 3511] = 'h00001fb3; 
    validation_data[ 3512] = 'h000018d5; 
    validation_data[ 3513] = 'h00003ebc; 
    validation_data[ 3514] = 'h000001f3; 
    validation_data[ 3515] = 'h00002f19; 
    validation_data[ 3516] = 'h00000f1b; 
    validation_data[ 3517] = 'h0000080f; 
    validation_data[ 3518] = 'h00002cdc; 
    validation_data[ 3519] = 'h000023df; 
    validation_data[ 3520] = 'h00000cc6; 
    validation_data[ 3521] = 'h00003b45; 
    validation_data[ 3522] = 'h00000dcb; 
    validation_data[ 3523] = 'h000005d7; 
    validation_data[ 3524] = 'h00003406; 
    validation_data[ 3525] = 'h00000218; 
    validation_data[ 3526] = 'h00000928; 
    validation_data[ 3527] = 'h00001e7f; 
    validation_data[ 3528] = 'h000036fb; 
    validation_data[ 3529] = 'h00003e16; 
    validation_data[ 3530] = 'h00003af4; 
    validation_data[ 3531] = 'h0000132e; 
    validation_data[ 3532] = 'h00000c77; 
    validation_data[ 3533] = 'h00003772; 
    validation_data[ 3534] = 'h0000095b; 
    validation_data[ 3535] = 'h00002b56; 
    validation_data[ 3536] = 'h0000378a; 
    validation_data[ 3537] = 'h0000395b; 
    validation_data[ 3538] = 'h00000aad; 
    validation_data[ 3539] = 'h0000305c; 
    validation_data[ 3540] = 'h00000670; 
    validation_data[ 3541] = 'h00001136; 
    validation_data[ 3542] = 'h00002073; 
    validation_data[ 3543] = 'h00000372; 
    validation_data[ 3544] = 'h0000246a; 
    validation_data[ 3545] = 'h00001509; 
    validation_data[ 3546] = 'h00000f22; 
    validation_data[ 3547] = 'h00000362; 
    validation_data[ 3548] = 'h00003841; 
    validation_data[ 3549] = 'h0000227f; 
    validation_data[ 3550] = 'h00002b00; 
    validation_data[ 3551] = 'h00003bab; 
    validation_data[ 3552] = 'h0000328a; 
    validation_data[ 3553] = 'h00002dd8; 
    validation_data[ 3554] = 'h00002c10; 
    validation_data[ 3555] = 'h000015c7; 
    validation_data[ 3556] = 'h000013b9; 
    validation_data[ 3557] = 'h00000393; 
    validation_data[ 3558] = 'h00003b9d; 
    validation_data[ 3559] = 'h00002702; 
    validation_data[ 3560] = 'h00001276; 
    validation_data[ 3561] = 'h000029b5; 
    validation_data[ 3562] = 'h0000265b; 
    validation_data[ 3563] = 'h000021c4; 
    validation_data[ 3564] = 'h000021b8; 
    validation_data[ 3565] = 'h00003a2a; 
    validation_data[ 3566] = 'h00003baf; 
    validation_data[ 3567] = 'h00000f4c; 
    validation_data[ 3568] = 'h00002832; 
    validation_data[ 3569] = 'h000015b5; 
    validation_data[ 3570] = 'h00000637; 
    validation_data[ 3571] = 'h00000f4c; 
    validation_data[ 3572] = 'h00002d5d; 
    validation_data[ 3573] = 'h00001663; 
    validation_data[ 3574] = 'h0000252b; 
    validation_data[ 3575] = 'h00001762; 
    validation_data[ 3576] = 'h00002de4; 
    validation_data[ 3577] = 'h00001cd4; 
    validation_data[ 3578] = 'h00001a13; 
    validation_data[ 3579] = 'h00002c45; 
    validation_data[ 3580] = 'h00001c06; 
    validation_data[ 3581] = 'h000039db; 
    validation_data[ 3582] = 'h0000102c; 
    validation_data[ 3583] = 'h00001f5d; 
    validation_data[ 3584] = 'h0000334f; 
    validation_data[ 3585] = 'h000036e0; 
    validation_data[ 3586] = 'h00002a17; 
    validation_data[ 3587] = 'h00000ef3; 
    validation_data[ 3588] = 'h0000043b; 
    validation_data[ 3589] = 'h00002b36; 
    validation_data[ 3590] = 'h000021ba; 
    validation_data[ 3591] = 'h000005ec; 
    validation_data[ 3592] = 'h000016e0; 
    validation_data[ 3593] = 'h00002b4b; 
    validation_data[ 3594] = 'h000008c2; 
    validation_data[ 3595] = 'h000007f3; 
    validation_data[ 3596] = 'h0000154b; 
    validation_data[ 3597] = 'h000029ae; 
    validation_data[ 3598] = 'h000034ab; 
    validation_data[ 3599] = 'h00001e32; 
    validation_data[ 3600] = 'h000025cf; 
    validation_data[ 3601] = 'h00000120; 
    validation_data[ 3602] = 'h0000025d; 
    validation_data[ 3603] = 'h00000706; 
    validation_data[ 3604] = 'h00002218; 
    validation_data[ 3605] = 'h00002404; 
    validation_data[ 3606] = 'h00001951; 
    validation_data[ 3607] = 'h0000206c; 
    validation_data[ 3608] = 'h000010d2; 
    validation_data[ 3609] = 'h00002ddd; 
    validation_data[ 3610] = 'h00002040; 
    validation_data[ 3611] = 'h00001786; 
    validation_data[ 3612] = 'h000006e2; 
    validation_data[ 3613] = 'h00000ae2; 
    validation_data[ 3614] = 'h000006e6; 
    validation_data[ 3615] = 'h00000b7c; 
    validation_data[ 3616] = 'h00000ecc; 
    validation_data[ 3617] = 'h0000045a; 
    validation_data[ 3618] = 'h0000253e; 
    validation_data[ 3619] = 'h0000011d; 
    validation_data[ 3620] = 'h0000232d; 
    validation_data[ 3621] = 'h0000150e; 
    validation_data[ 3622] = 'h0000370f; 
    validation_data[ 3623] = 'h00001290; 
    validation_data[ 3624] = 'h000018ac; 
    validation_data[ 3625] = 'h00003397; 
    validation_data[ 3626] = 'h00001365; 
    validation_data[ 3627] = 'h00000237; 
    validation_data[ 3628] = 'h00002769; 
    validation_data[ 3629] = 'h00000f45; 
    validation_data[ 3630] = 'h000035dd; 
    validation_data[ 3631] = 'h0000202e; 
    validation_data[ 3632] = 'h0000003a; 
    validation_data[ 3633] = 'h0000291b; 
    validation_data[ 3634] = 'h00000a41; 
    validation_data[ 3635] = 'h00001aad; 
    validation_data[ 3636] = 'h00002373; 
    validation_data[ 3637] = 'h00000e93; 
    validation_data[ 3638] = 'h00000e3e; 
    validation_data[ 3639] = 'h000004ff; 
    validation_data[ 3640] = 'h00000ad9; 
    validation_data[ 3641] = 'h0000246c; 
    validation_data[ 3642] = 'h000037d3; 
    validation_data[ 3643] = 'h00002d00; 
    validation_data[ 3644] = 'h00001ac4; 
    validation_data[ 3645] = 'h000017e2; 
    validation_data[ 3646] = 'h00002428; 
    validation_data[ 3647] = 'h00000656; 
    validation_data[ 3648] = 'h00000df7; 
    validation_data[ 3649] = 'h0000021f; 
    validation_data[ 3650] = 'h00000106; 
    validation_data[ 3651] = 'h00001cd0; 
    validation_data[ 3652] = 'h000005e2; 
    validation_data[ 3653] = 'h00000434; 
    validation_data[ 3654] = 'h00003f5f; 
    validation_data[ 3655] = 'h00002142; 
    validation_data[ 3656] = 'h00001183; 
    validation_data[ 3657] = 'h00003ed2; 
    validation_data[ 3658] = 'h000003fa; 
    validation_data[ 3659] = 'h00003c09; 
    validation_data[ 3660] = 'h0000176a; 
    validation_data[ 3661] = 'h00003717; 
    validation_data[ 3662] = 'h000034f6; 
    validation_data[ 3663] = 'h0000342a; 
    validation_data[ 3664] = 'h00000358; 
    validation_data[ 3665] = 'h00001c38; 
    validation_data[ 3666] = 'h00003e55; 
    validation_data[ 3667] = 'h000005fe; 
    validation_data[ 3668] = 'h0000199f; 
    validation_data[ 3669] = 'h0000057c; 
    validation_data[ 3670] = 'h0000103b; 
    validation_data[ 3671] = 'h000021c7; 
    validation_data[ 3672] = 'h00003c6f; 
    validation_data[ 3673] = 'h000028c0; 
    validation_data[ 3674] = 'h0000066d; 
    validation_data[ 3675] = 'h000003c6; 
    validation_data[ 3676] = 'h00003b2d; 
    validation_data[ 3677] = 'h00003fdd; 
    validation_data[ 3678] = 'h00003d51; 
    validation_data[ 3679] = 'h00001c09; 
    validation_data[ 3680] = 'h000028bb; 
    validation_data[ 3681] = 'h0000000c; 
    validation_data[ 3682] = 'h00001381; 
    validation_data[ 3683] = 'h00003f17; 
    validation_data[ 3684] = 'h00003528; 
    validation_data[ 3685] = 'h00000be2; 
    validation_data[ 3686] = 'h00003d4f; 
    validation_data[ 3687] = 'h00002b03; 
    validation_data[ 3688] = 'h00002ab6; 
    validation_data[ 3689] = 'h00001e4c; 
    validation_data[ 3690] = 'h00000621; 
    validation_data[ 3691] = 'h00003ac3; 
    validation_data[ 3692] = 'h00001e05; 
    validation_data[ 3693] = 'h0000161a; 
    validation_data[ 3694] = 'h000004b7; 
    validation_data[ 3695] = 'h00000e67; 
    validation_data[ 3696] = 'h0000130a; 
    validation_data[ 3697] = 'h00003a8d; 
    validation_data[ 3698] = 'h00000d73; 
    validation_data[ 3699] = 'h00000653; 
    validation_data[ 3700] = 'h00002813; 
    validation_data[ 3701] = 'h00003e9c; 
    validation_data[ 3702] = 'h00001ec0; 
    validation_data[ 3703] = 'h00002d97; 
    validation_data[ 3704] = 'h000025ae; 
    validation_data[ 3705] = 'h00000054; 
    validation_data[ 3706] = 'h00002fe3; 
    validation_data[ 3707] = 'h00003974; 
    validation_data[ 3708] = 'h00001c9b; 
    validation_data[ 3709] = 'h000003da; 
    validation_data[ 3710] = 'h000019fa; 
    validation_data[ 3711] = 'h0000226b; 
    validation_data[ 3712] = 'h00002f27; 
    validation_data[ 3713] = 'h000007f7; 
    validation_data[ 3714] = 'h00000b91; 
    validation_data[ 3715] = 'h000012ff; 
    validation_data[ 3716] = 'h000031d0; 
    validation_data[ 3717] = 'h00001f6a; 
    validation_data[ 3718] = 'h00003270; 
    validation_data[ 3719] = 'h000008b5; 
    validation_data[ 3720] = 'h00002714; 
    validation_data[ 3721] = 'h00002480; 
    validation_data[ 3722] = 'h00002ed9; 
    validation_data[ 3723] = 'h000014b9; 
    validation_data[ 3724] = 'h00003283; 
    validation_data[ 3725] = 'h00002eb7; 
    validation_data[ 3726] = 'h0000260d; 
    validation_data[ 3727] = 'h00000394; 
    validation_data[ 3728] = 'h00001d0c; 
    validation_data[ 3729] = 'h00002913; 
    validation_data[ 3730] = 'h00001323; 
    validation_data[ 3731] = 'h00000c25; 
    validation_data[ 3732] = 'h00001552; 
    validation_data[ 3733] = 'h00003dd8; 
    validation_data[ 3734] = 'h00001ec5; 
    validation_data[ 3735] = 'h00000948; 
    validation_data[ 3736] = 'h000030e4; 
    validation_data[ 3737] = 'h00003636; 
    validation_data[ 3738] = 'h00003294; 
    validation_data[ 3739] = 'h000032e7; 
    validation_data[ 3740] = 'h000033d8; 
    validation_data[ 3741] = 'h00000b77; 
    validation_data[ 3742] = 'h00002a67; 
    validation_data[ 3743] = 'h00003185; 
    validation_data[ 3744] = 'h00001394; 
    validation_data[ 3745] = 'h00000d62; 
    validation_data[ 3746] = 'h000007dc; 
    validation_data[ 3747] = 'h000022bb; 
    validation_data[ 3748] = 'h00000845; 
    validation_data[ 3749] = 'h0000261a; 
    validation_data[ 3750] = 'h00003846; 
    validation_data[ 3751] = 'h00001a06; 
    validation_data[ 3752] = 'h0000341a; 
    validation_data[ 3753] = 'h00000f3d; 
    validation_data[ 3754] = 'h00001ebb; 
    validation_data[ 3755] = 'h00001b14; 
    validation_data[ 3756] = 'h00002dd0; 
    validation_data[ 3757] = 'h00002c1b; 
    validation_data[ 3758] = 'h00003054; 
    validation_data[ 3759] = 'h00001b85; 
    validation_data[ 3760] = 'h000020df; 
    validation_data[ 3761] = 'h00002b10; 
    validation_data[ 3762] = 'h000016d3; 
    validation_data[ 3763] = 'h00002035; 
    validation_data[ 3764] = 'h00002196; 
    validation_data[ 3765] = 'h00000963; 
    validation_data[ 3766] = 'h000016aa; 
    validation_data[ 3767] = 'h00000640; 
    validation_data[ 3768] = 'h00003425; 
    validation_data[ 3769] = 'h00001c38; 
    validation_data[ 3770] = 'h00002b8e; 
    validation_data[ 3771] = 'h00001452; 
    validation_data[ 3772] = 'h00001686; 
    validation_data[ 3773] = 'h00000a71; 
    validation_data[ 3774] = 'h00003dec; 
    validation_data[ 3775] = 'h00003870; 
    validation_data[ 3776] = 'h00000029; 
    validation_data[ 3777] = 'h000000c1; 
    validation_data[ 3778] = 'h00002675; 
    validation_data[ 3779] = 'h00000666; 
    validation_data[ 3780] = 'h00001eba; 
    validation_data[ 3781] = 'h0000127c; 
    validation_data[ 3782] = 'h00001f23; 
    validation_data[ 3783] = 'h00000af1; 
    validation_data[ 3784] = 'h000001b0; 
    validation_data[ 3785] = 'h0000040a; 
    validation_data[ 3786] = 'h00002fce; 
    validation_data[ 3787] = 'h00003ee3; 
    validation_data[ 3788] = 'h00000dcb; 
    validation_data[ 3789] = 'h00000079; 
    validation_data[ 3790] = 'h00000cd0; 
    validation_data[ 3791] = 'h00002a18; 
    validation_data[ 3792] = 'h00001ca5; 
    validation_data[ 3793] = 'h00001875; 
    validation_data[ 3794] = 'h000005fc; 
    validation_data[ 3795] = 'h000007a6; 
    validation_data[ 3796] = 'h00002ae5; 
    validation_data[ 3797] = 'h0000232a; 
    validation_data[ 3798] = 'h00001e12; 
    validation_data[ 3799] = 'h0000166f; 
    validation_data[ 3800] = 'h000023f5; 
    validation_data[ 3801] = 'h00000928; 
    validation_data[ 3802] = 'h0000165d; 
    validation_data[ 3803] = 'h00003302; 
    validation_data[ 3804] = 'h00000a58; 
    validation_data[ 3805] = 'h00001368; 
    validation_data[ 3806] = 'h000012ff; 
    validation_data[ 3807] = 'h00003213; 
    validation_data[ 3808] = 'h000023f4; 
    validation_data[ 3809] = 'h00002556; 
    validation_data[ 3810] = 'h00001582; 
    validation_data[ 3811] = 'h00003eb2; 
    validation_data[ 3812] = 'h00002a33; 
    validation_data[ 3813] = 'h00003c86; 
    validation_data[ 3814] = 'h00000d55; 
    validation_data[ 3815] = 'h00003489; 
    validation_data[ 3816] = 'h00002af2; 
    validation_data[ 3817] = 'h0000065a; 
    validation_data[ 3818] = 'h00001935; 
    validation_data[ 3819] = 'h00003536; 
    validation_data[ 3820] = 'h00003512; 
    validation_data[ 3821] = 'h00001f35; 
    validation_data[ 3822] = 'h000030b1; 
    validation_data[ 3823] = 'h00001e82; 
    validation_data[ 3824] = 'h000022c6; 
    validation_data[ 3825] = 'h00002218; 
    validation_data[ 3826] = 'h00000f3b; 
    validation_data[ 3827] = 'h00003b5f; 
    validation_data[ 3828] = 'h00002107; 
    validation_data[ 3829] = 'h00003fb6; 
    validation_data[ 3830] = 'h000031f2; 
    validation_data[ 3831] = 'h00000c49; 
    validation_data[ 3832] = 'h00000737; 
    validation_data[ 3833] = 'h00002ffc; 
    validation_data[ 3834] = 'h00001d65; 
    validation_data[ 3835] = 'h00003fd9; 
    validation_data[ 3836] = 'h00003ca1; 
    validation_data[ 3837] = 'h00002918; 
    validation_data[ 3838] = 'h00001be8; 
    validation_data[ 3839] = 'h00000bd2; 
    validation_data[ 3840] = 'h00000c75; 
    validation_data[ 3841] = 'h00002967; 
    validation_data[ 3842] = 'h00001c3a; 
    validation_data[ 3843] = 'h0000090a; 
    validation_data[ 3844] = 'h00000684; 
    validation_data[ 3845] = 'h000034a1; 
    validation_data[ 3846] = 'h0000012a; 
    validation_data[ 3847] = 'h00003ddf; 
    validation_data[ 3848] = 'h000000fa; 
    validation_data[ 3849] = 'h00001b6e; 
    validation_data[ 3850] = 'h000022bf; 
    validation_data[ 3851] = 'h00002912; 
    validation_data[ 3852] = 'h000023aa; 
    validation_data[ 3853] = 'h00000061; 
    validation_data[ 3854] = 'h00002a28; 
    validation_data[ 3855] = 'h000014c0; 
    validation_data[ 3856] = 'h00001177; 
    validation_data[ 3857] = 'h00002580; 
    validation_data[ 3858] = 'h00002d9b; 
    validation_data[ 3859] = 'h00003f13; 
    validation_data[ 3860] = 'h00002108; 
    validation_data[ 3861] = 'h00000a19; 
    validation_data[ 3862] = 'h0000094f; 
    validation_data[ 3863] = 'h00000ec7; 
    validation_data[ 3864] = 'h00001404; 
    validation_data[ 3865] = 'h00001914; 
    validation_data[ 3866] = 'h00001389; 
    validation_data[ 3867] = 'h000003aa; 
    validation_data[ 3868] = 'h00000117; 
    validation_data[ 3869] = 'h0000113d; 
    validation_data[ 3870] = 'h000016ba; 
    validation_data[ 3871] = 'h00000893; 
    validation_data[ 3872] = 'h000038c0; 
    validation_data[ 3873] = 'h0000050c; 
    validation_data[ 3874] = 'h000037ad; 
    validation_data[ 3875] = 'h0000061c; 
    validation_data[ 3876] = 'h0000076a; 
    validation_data[ 3877] = 'h000009e7; 
    validation_data[ 3878] = 'h00003491; 
    validation_data[ 3879] = 'h00000fda; 
    validation_data[ 3880] = 'h00003316; 
    validation_data[ 3881] = 'h00002426; 
    validation_data[ 3882] = 'h00003e01; 
    validation_data[ 3883] = 'h0000176f; 
    validation_data[ 3884] = 'h00003b6d; 
    validation_data[ 3885] = 'h00003a09; 
    validation_data[ 3886] = 'h00003908; 
    validation_data[ 3887] = 'h00000a25; 
    validation_data[ 3888] = 'h000006b9; 
    validation_data[ 3889] = 'h00002d7f; 
    validation_data[ 3890] = 'h0000351c; 
    validation_data[ 3891] = 'h00000d70; 
    validation_data[ 3892] = 'h00000625; 
    validation_data[ 3893] = 'h00003f3b; 
    validation_data[ 3894] = 'h000002dd; 
    validation_data[ 3895] = 'h000020e1; 
    validation_data[ 3896] = 'h00000694; 
    validation_data[ 3897] = 'h000000cc; 
    validation_data[ 3898] = 'h00000ed9; 
    validation_data[ 3899] = 'h0000322d; 
    validation_data[ 3900] = 'h0000123c; 
    validation_data[ 3901] = 'h00000e06; 
    validation_data[ 3902] = 'h000033dc; 
    validation_data[ 3903] = 'h000039a2; 
    validation_data[ 3904] = 'h00002ae9; 
    validation_data[ 3905] = 'h00000fb6; 
    validation_data[ 3906] = 'h00000a34; 
    validation_data[ 3907] = 'h00000ba7; 
    validation_data[ 3908] = 'h00002805; 
    validation_data[ 3909] = 'h00002623; 
    validation_data[ 3910] = 'h000020fd; 
    validation_data[ 3911] = 'h000028cd; 
    validation_data[ 3912] = 'h000014d9; 
    validation_data[ 3913] = 'h000007d1; 
    validation_data[ 3914] = 'h000025e5; 
    validation_data[ 3915] = 'h00002b97; 
    validation_data[ 3916] = 'h000038dd; 
    validation_data[ 3917] = 'h00001999; 
    validation_data[ 3918] = 'h00000273; 
    validation_data[ 3919] = 'h000031c2; 
    validation_data[ 3920] = 'h000027ad; 
    validation_data[ 3921] = 'h000010cf; 
    validation_data[ 3922] = 'h00000323; 
    validation_data[ 3923] = 'h00001d52; 
    validation_data[ 3924] = 'h00002947; 
    validation_data[ 3925] = 'h000033fc; 
    validation_data[ 3926] = 'h00002f12; 
    validation_data[ 3927] = 'h000011b4; 
    validation_data[ 3928] = 'h000027de; 
    validation_data[ 3929] = 'h00002b5f; 
    validation_data[ 3930] = 'h00003550; 
    validation_data[ 3931] = 'h00002126; 
    validation_data[ 3932] = 'h00002024; 
    validation_data[ 3933] = 'h00000263; 
    validation_data[ 3934] = 'h000025be; 
    validation_data[ 3935] = 'h00003995; 
    validation_data[ 3936] = 'h00000f7e; 
    validation_data[ 3937] = 'h00000d3c; 
    validation_data[ 3938] = 'h0000244e; 
    validation_data[ 3939] = 'h000010ba; 
    validation_data[ 3940] = 'h000030c2; 
    validation_data[ 3941] = 'h00002928; 
    validation_data[ 3942] = 'h000036c1; 
    validation_data[ 3943] = 'h0000388a; 
    validation_data[ 3944] = 'h00000bbc; 
    validation_data[ 3945] = 'h0000138e; 
    validation_data[ 3946] = 'h00000136; 
    validation_data[ 3947] = 'h0000228a; 
    validation_data[ 3948] = 'h000008f4; 
    validation_data[ 3949] = 'h00001ae6; 
    validation_data[ 3950] = 'h0000354c; 
    validation_data[ 3951] = 'h00003bf1; 
    validation_data[ 3952] = 'h0000147c; 
    validation_data[ 3953] = 'h000025fc; 
    validation_data[ 3954] = 'h00001bd3; 
    validation_data[ 3955] = 'h00003c1c; 
    validation_data[ 3956] = 'h00001f7b; 
    validation_data[ 3957] = 'h00003ac2; 
    validation_data[ 3958] = 'h00003e83; 
    validation_data[ 3959] = 'h00000d1c; 
    validation_data[ 3960] = 'h00003b99; 
    validation_data[ 3961] = 'h00000318; 
    validation_data[ 3962] = 'h000024c7; 
    validation_data[ 3963] = 'h0000268d; 
    validation_data[ 3964] = 'h0000059e; 
    validation_data[ 3965] = 'h00000a5c; 
    validation_data[ 3966] = 'h00000a9c; 
    validation_data[ 3967] = 'h00001790; 
    validation_data[ 3968] = 'h0000021b; 
    validation_data[ 3969] = 'h0000263d; 
    validation_data[ 3970] = 'h00001ae1; 
    validation_data[ 3971] = 'h000015ff; 
    validation_data[ 3972] = 'h0000272f; 
    validation_data[ 3973] = 'h0000375e; 
    validation_data[ 3974] = 'h00000e77; 
    validation_data[ 3975] = 'h0000347d; 
    validation_data[ 3976] = 'h00002784; 
    validation_data[ 3977] = 'h000015a5; 
    validation_data[ 3978] = 'h00003731; 
    validation_data[ 3979] = 'h00000fb9; 
    validation_data[ 3980] = 'h00002008; 
    validation_data[ 3981] = 'h000003c5; 
    validation_data[ 3982] = 'h00003f29; 
    validation_data[ 3983] = 'h00001dfc; 
    validation_data[ 3984] = 'h000011c4; 
    validation_data[ 3985] = 'h00003717; 
    validation_data[ 3986] = 'h00001e1b; 
    validation_data[ 3987] = 'h0000248e; 
    validation_data[ 3988] = 'h00000e46; 
    validation_data[ 3989] = 'h000029e4; 
    validation_data[ 3990] = 'h000037b1; 
    validation_data[ 3991] = 'h0000340d; 
    validation_data[ 3992] = 'h00002f27; 
    validation_data[ 3993] = 'h0000155c; 
    validation_data[ 3994] = 'h000039f2; 
    validation_data[ 3995] = 'h00000bcc; 
    validation_data[ 3996] = 'h0000318d; 
    validation_data[ 3997] = 'h00003c88; 
    validation_data[ 3998] = 'h0000376b; 
    validation_data[ 3999] = 'h00000cb5; 
    validation_data[ 4000] = 'h00003eba; 
    validation_data[ 4001] = 'h00000238; 
    validation_data[ 4002] = 'h00002353; 
    validation_data[ 4003] = 'h00003fb5; 
    validation_data[ 4004] = 'h00001030; 
    validation_data[ 4005] = 'h00001798; 
    validation_data[ 4006] = 'h00001d39; 
    validation_data[ 4007] = 'h00001d12; 
    validation_data[ 4008] = 'h00001b27; 
    validation_data[ 4009] = 'h00001b38; 
    validation_data[ 4010] = 'h000023de; 
    validation_data[ 4011] = 'h000020e2; 
    validation_data[ 4012] = 'h00002c60; 
    validation_data[ 4013] = 'h000034d6; 
    validation_data[ 4014] = 'h000015a2; 
    validation_data[ 4015] = 'h00000596; 
    validation_data[ 4016] = 'h000037ab; 
    validation_data[ 4017] = 'h000011ef; 
    validation_data[ 4018] = 'h00002f24; 
    validation_data[ 4019] = 'h00003e87; 
    validation_data[ 4020] = 'h00001eb0; 
    validation_data[ 4021] = 'h00002651; 
    validation_data[ 4022] = 'h00000f1e; 
    validation_data[ 4023] = 'h00003008; 
    validation_data[ 4024] = 'h00000166; 
    validation_data[ 4025] = 'h00002344; 
    validation_data[ 4026] = 'h00003af6; 
    validation_data[ 4027] = 'h000037e0; 
    validation_data[ 4028] = 'h00001b71; 
    validation_data[ 4029] = 'h00002e6e; 
    validation_data[ 4030] = 'h00000863; 
    validation_data[ 4031] = 'h00003022; 
    validation_data[ 4032] = 'h00002e31; 
    validation_data[ 4033] = 'h00003cf7; 
    validation_data[ 4034] = 'h00001762; 
    validation_data[ 4035] = 'h0000220a; 
    validation_data[ 4036] = 'h00003ef7; 
    validation_data[ 4037] = 'h000015a4; 
    validation_data[ 4038] = 'h0000070e; 
    validation_data[ 4039] = 'h0000292a; 
    validation_data[ 4040] = 'h00003d4b; 
    validation_data[ 4041] = 'h00002eba; 
    validation_data[ 4042] = 'h0000127e; 
    validation_data[ 4043] = 'h00000f03; 
    validation_data[ 4044] = 'h00002c7b; 
    validation_data[ 4045] = 'h000014c8; 
    validation_data[ 4046] = 'h00000cb0; 
    validation_data[ 4047] = 'h0000321e; 
    validation_data[ 4048] = 'h0000075c; 
    validation_data[ 4049] = 'h00000f16; 
    validation_data[ 4050] = 'h000027fe; 
    validation_data[ 4051] = 'h00003dd5; 
    validation_data[ 4052] = 'h000031b4; 
    validation_data[ 4053] = 'h0000140d; 
    validation_data[ 4054] = 'h00000932; 
    validation_data[ 4055] = 'h000038b5; 
    validation_data[ 4056] = 'h00003cfb; 
    validation_data[ 4057] = 'h00000a82; 
    validation_data[ 4058] = 'h0000146d; 
    validation_data[ 4059] = 'h00003965; 
    validation_data[ 4060] = 'h000016cf; 
    validation_data[ 4061] = 'h000000fc; 
    validation_data[ 4062] = 'h00000211; 
    validation_data[ 4063] = 'h00002583; 
    validation_data[ 4064] = 'h00003dee; 
    validation_data[ 4065] = 'h00001192; 
    validation_data[ 4066] = 'h0000162b; 
    validation_data[ 4067] = 'h00002696; 
    validation_data[ 4068] = 'h00002e4d; 
    validation_data[ 4069] = 'h00000685; 
    validation_data[ 4070] = 'h00002cbd; 
    validation_data[ 4071] = 'h00001065; 
    validation_data[ 4072] = 'h00002f3f; 
    validation_data[ 4073] = 'h00003798; 
    validation_data[ 4074] = 'h000034d5; 
    validation_data[ 4075] = 'h00001350; 
    validation_data[ 4076] = 'h00002461; 
    validation_data[ 4077] = 'h00002593; 
    validation_data[ 4078] = 'h00003ac3; 
    validation_data[ 4079] = 'h00001362; 
    validation_data[ 4080] = 'h000036c3; 
    validation_data[ 4081] = 'h00001e4f; 
    validation_data[ 4082] = 'h000034d3; 
    validation_data[ 4083] = 'h00001cc8; 
    validation_data[ 4084] = 'h00001884; 
    validation_data[ 4085] = 'h00000d20; 
    validation_data[ 4086] = 'h0000105d; 
    validation_data[ 4087] = 'h00000ee7; 
    validation_data[ 4088] = 'h0000070b; 
    validation_data[ 4089] = 'h000035a5; 
    validation_data[ 4090] = 'h000009ce; 
    validation_data[ 4091] = 'h00003e0e; 
    validation_data[ 4092] = 'h00001f7f; 
    validation_data[ 4093] = 'h00000d7b; 
    validation_data[ 4094] = 'h00001a1f; 
    validation_data[ 4095] = 'h000033ed; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule


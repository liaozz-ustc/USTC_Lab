
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h85efb51f;
    ram_cell[       1] = 32'h0;  // 32'hb0d237fc;
    ram_cell[       2] = 32'h0;  // 32'h45b9b456;
    ram_cell[       3] = 32'h0;  // 32'h6460b4f1;
    ram_cell[       4] = 32'h0;  // 32'h6f593d55;
    ram_cell[       5] = 32'h0;  // 32'hd96e0092;
    ram_cell[       6] = 32'h0;  // 32'hca6382f4;
    ram_cell[       7] = 32'h0;  // 32'h5729e353;
    ram_cell[       8] = 32'h0;  // 32'he896098f;
    ram_cell[       9] = 32'h0;  // 32'hd5c60a42;
    ram_cell[      10] = 32'h0;  // 32'h918d52cd;
    ram_cell[      11] = 32'h0;  // 32'h59307caf;
    ram_cell[      12] = 32'h0;  // 32'hcd9ecb6a;
    ram_cell[      13] = 32'h0;  // 32'h649194a4;
    ram_cell[      14] = 32'h0;  // 32'hb28e9213;
    ram_cell[      15] = 32'h0;  // 32'h9a2469b4;
    ram_cell[      16] = 32'h0;  // 32'hb8f81c4e;
    ram_cell[      17] = 32'h0;  // 32'h67ac76b4;
    ram_cell[      18] = 32'h0;  // 32'h906387e8;
    ram_cell[      19] = 32'h0;  // 32'hcc4ab185;
    ram_cell[      20] = 32'h0;  // 32'h2bf5b618;
    ram_cell[      21] = 32'h0;  // 32'hfd2610fc;
    ram_cell[      22] = 32'h0;  // 32'hce128811;
    ram_cell[      23] = 32'h0;  // 32'h4dee0a65;
    ram_cell[      24] = 32'h0;  // 32'hfe953dc0;
    ram_cell[      25] = 32'h0;  // 32'he2108e68;
    ram_cell[      26] = 32'h0;  // 32'h9f8ec77d;
    ram_cell[      27] = 32'h0;  // 32'h9e8e6809;
    ram_cell[      28] = 32'h0;  // 32'hcacd03f4;
    ram_cell[      29] = 32'h0;  // 32'h09de8c54;
    ram_cell[      30] = 32'h0;  // 32'h6354078f;
    ram_cell[      31] = 32'h0;  // 32'h4a6ae60b;
    ram_cell[      32] = 32'h0;  // 32'h82401255;
    ram_cell[      33] = 32'h0;  // 32'hd097f6e3;
    ram_cell[      34] = 32'h0;  // 32'h4ff166fe;
    ram_cell[      35] = 32'h0;  // 32'he1a1b122;
    ram_cell[      36] = 32'h0;  // 32'hd80e32f2;
    ram_cell[      37] = 32'h0;  // 32'hf73e1be3;
    ram_cell[      38] = 32'h0;  // 32'hf008a5d2;
    ram_cell[      39] = 32'h0;  // 32'hc4686370;
    ram_cell[      40] = 32'h0;  // 32'h4a95434c;
    ram_cell[      41] = 32'h0;  // 32'h07876318;
    ram_cell[      42] = 32'h0;  // 32'h532aaa8b;
    ram_cell[      43] = 32'h0;  // 32'h58257457;
    ram_cell[      44] = 32'h0;  // 32'h22f20888;
    ram_cell[      45] = 32'h0;  // 32'h1bed4edd;
    ram_cell[      46] = 32'h0;  // 32'he92aa070;
    ram_cell[      47] = 32'h0;  // 32'h84d641d6;
    ram_cell[      48] = 32'h0;  // 32'h9ad3b21a;
    ram_cell[      49] = 32'h0;  // 32'h34bb62c5;
    ram_cell[      50] = 32'h0;  // 32'h78bb0d2c;
    ram_cell[      51] = 32'h0;  // 32'h3ad8a8b3;
    ram_cell[      52] = 32'h0;  // 32'hbc74f080;
    ram_cell[      53] = 32'h0;  // 32'hb2e953b8;
    ram_cell[      54] = 32'h0;  // 32'hade79d2f;
    ram_cell[      55] = 32'h0;  // 32'h6c1aa1b3;
    ram_cell[      56] = 32'h0;  // 32'h96466344;
    ram_cell[      57] = 32'h0;  // 32'h61094b62;
    ram_cell[      58] = 32'h0;  // 32'h7ae378e0;
    ram_cell[      59] = 32'h0;  // 32'hb7390d2d;
    ram_cell[      60] = 32'h0;  // 32'h0ba5fe3a;
    ram_cell[      61] = 32'h0;  // 32'h15be617d;
    ram_cell[      62] = 32'h0;  // 32'hcb8afcfe;
    ram_cell[      63] = 32'h0;  // 32'h8ef47f0c;
    ram_cell[      64] = 32'h0;  // 32'h577cc574;
    ram_cell[      65] = 32'h0;  // 32'hc8d81bd2;
    ram_cell[      66] = 32'h0;  // 32'h5fc293af;
    ram_cell[      67] = 32'h0;  // 32'h87d0210d;
    ram_cell[      68] = 32'h0;  // 32'h616fbf6d;
    ram_cell[      69] = 32'h0;  // 32'hbd9fd4c9;
    ram_cell[      70] = 32'h0;  // 32'hbc10fcb1;
    ram_cell[      71] = 32'h0;  // 32'h5bf8819a;
    ram_cell[      72] = 32'h0;  // 32'h9325cb09;
    ram_cell[      73] = 32'h0;  // 32'h7e9fd9cc;
    ram_cell[      74] = 32'h0;  // 32'h5eba5d0f;
    ram_cell[      75] = 32'h0;  // 32'h49270ca3;
    ram_cell[      76] = 32'h0;  // 32'hd87b632f;
    ram_cell[      77] = 32'h0;  // 32'hd36b75d4;
    ram_cell[      78] = 32'h0;  // 32'hcfa324a1;
    ram_cell[      79] = 32'h0;  // 32'h80c27018;
    ram_cell[      80] = 32'h0;  // 32'hb5e5b9f5;
    ram_cell[      81] = 32'h0;  // 32'h2f184f29;
    ram_cell[      82] = 32'h0;  // 32'h9b8d1fc4;
    ram_cell[      83] = 32'h0;  // 32'h64cdb801;
    ram_cell[      84] = 32'h0;  // 32'h700950c3;
    ram_cell[      85] = 32'h0;  // 32'hf20751b1;
    ram_cell[      86] = 32'h0;  // 32'h231cb4ad;
    ram_cell[      87] = 32'h0;  // 32'h24581a44;
    ram_cell[      88] = 32'h0;  // 32'hc78e55a0;
    ram_cell[      89] = 32'h0;  // 32'hebad9bd7;
    ram_cell[      90] = 32'h0;  // 32'h9f74e02b;
    ram_cell[      91] = 32'h0;  // 32'h24063339;
    ram_cell[      92] = 32'h0;  // 32'h9a984248;
    ram_cell[      93] = 32'h0;  // 32'hc005297b;
    ram_cell[      94] = 32'h0;  // 32'hb69e4959;
    ram_cell[      95] = 32'h0;  // 32'hb02a9a88;
    ram_cell[      96] = 32'h0;  // 32'h28492746;
    ram_cell[      97] = 32'h0;  // 32'h2e9a5e4a;
    ram_cell[      98] = 32'h0;  // 32'h5b2bb9d7;
    ram_cell[      99] = 32'h0;  // 32'haed2e42d;
    ram_cell[     100] = 32'h0;  // 32'h6d1d7abf;
    ram_cell[     101] = 32'h0;  // 32'h5d77c813;
    ram_cell[     102] = 32'h0;  // 32'h44db699e;
    ram_cell[     103] = 32'h0;  // 32'hf30fb986;
    ram_cell[     104] = 32'h0;  // 32'he19149d5;
    ram_cell[     105] = 32'h0;  // 32'h946e30a6;
    ram_cell[     106] = 32'h0;  // 32'h3f368fcf;
    ram_cell[     107] = 32'h0;  // 32'hed78fa75;
    ram_cell[     108] = 32'h0;  // 32'ha37e48b5;
    ram_cell[     109] = 32'h0;  // 32'ha950d7d3;
    ram_cell[     110] = 32'h0;  // 32'h45d64741;
    ram_cell[     111] = 32'h0;  // 32'hc688bcaf;
    ram_cell[     112] = 32'h0;  // 32'haa95c183;
    ram_cell[     113] = 32'h0;  // 32'h47e0629f;
    ram_cell[     114] = 32'h0;  // 32'ha71d87ce;
    ram_cell[     115] = 32'h0;  // 32'haf263c51;
    ram_cell[     116] = 32'h0;  // 32'hf525cb93;
    ram_cell[     117] = 32'h0;  // 32'h8cce3dda;
    ram_cell[     118] = 32'h0;  // 32'hc6b1724c;
    ram_cell[     119] = 32'h0;  // 32'h47fdc2a6;
    ram_cell[     120] = 32'h0;  // 32'he62eb815;
    ram_cell[     121] = 32'h0;  // 32'h7d175383;
    ram_cell[     122] = 32'h0;  // 32'h66d61aa4;
    ram_cell[     123] = 32'h0;  // 32'h087dada5;
    ram_cell[     124] = 32'h0;  // 32'h7523156b;
    ram_cell[     125] = 32'h0;  // 32'h8bba573f;
    ram_cell[     126] = 32'h0;  // 32'h6c7df225;
    ram_cell[     127] = 32'h0;  // 32'h8ee432e7;
    ram_cell[     128] = 32'h0;  // 32'h93b0bf4d;
    ram_cell[     129] = 32'h0;  // 32'hedcb7013;
    ram_cell[     130] = 32'h0;  // 32'h12276712;
    ram_cell[     131] = 32'h0;  // 32'he494ebb8;
    ram_cell[     132] = 32'h0;  // 32'hc0530f91;
    ram_cell[     133] = 32'h0;  // 32'h056ad6d2;
    ram_cell[     134] = 32'h0;  // 32'h37e100d6;
    ram_cell[     135] = 32'h0;  // 32'ha87e934b;
    ram_cell[     136] = 32'h0;  // 32'h9045b3ae;
    ram_cell[     137] = 32'h0;  // 32'h12a423ea;
    ram_cell[     138] = 32'h0;  // 32'hcc3163d2;
    ram_cell[     139] = 32'h0;  // 32'h6587d462;
    ram_cell[     140] = 32'h0;  // 32'h8598d32b;
    ram_cell[     141] = 32'h0;  // 32'h8c3111a9;
    ram_cell[     142] = 32'h0;  // 32'h9d364634;
    ram_cell[     143] = 32'h0;  // 32'h301e8718;
    ram_cell[     144] = 32'h0;  // 32'hbac4e1a0;
    ram_cell[     145] = 32'h0;  // 32'h6af1ca6d;
    ram_cell[     146] = 32'h0;  // 32'h468d49ba;
    ram_cell[     147] = 32'h0;  // 32'hf7ae0c27;
    ram_cell[     148] = 32'h0;  // 32'hfd79fc3f;
    ram_cell[     149] = 32'h0;  // 32'h64036e3f;
    ram_cell[     150] = 32'h0;  // 32'h8cd33cdd;
    ram_cell[     151] = 32'h0;  // 32'h3feb4467;
    ram_cell[     152] = 32'h0;  // 32'hb539cb05;
    ram_cell[     153] = 32'h0;  // 32'ha5d96991;
    ram_cell[     154] = 32'h0;  // 32'h565581f8;
    ram_cell[     155] = 32'h0;  // 32'h9db96d29;
    ram_cell[     156] = 32'h0;  // 32'hc50a8dee;
    ram_cell[     157] = 32'h0;  // 32'h14ca5693;
    ram_cell[     158] = 32'h0;  // 32'h01b28faa;
    ram_cell[     159] = 32'h0;  // 32'h5ef5d637;
    ram_cell[     160] = 32'h0;  // 32'h34287bb6;
    ram_cell[     161] = 32'h0;  // 32'h279a27e0;
    ram_cell[     162] = 32'h0;  // 32'h85bc0ce9;
    ram_cell[     163] = 32'h0;  // 32'h3d66c174;
    ram_cell[     164] = 32'h0;  // 32'h668d864f;
    ram_cell[     165] = 32'h0;  // 32'hb86f34c2;
    ram_cell[     166] = 32'h0;  // 32'h3b2fe7a8;
    ram_cell[     167] = 32'h0;  // 32'hec0564be;
    ram_cell[     168] = 32'h0;  // 32'h25ae5f75;
    ram_cell[     169] = 32'h0;  // 32'ha85f4dd3;
    ram_cell[     170] = 32'h0;  // 32'h59e9e581;
    ram_cell[     171] = 32'h0;  // 32'h0f159830;
    ram_cell[     172] = 32'h0;  // 32'h1441abc3;
    ram_cell[     173] = 32'h0;  // 32'hdb7ab1be;
    ram_cell[     174] = 32'h0;  // 32'h54d55ddf;
    ram_cell[     175] = 32'h0;  // 32'h00cae3b9;
    ram_cell[     176] = 32'h0;  // 32'h38b7171f;
    ram_cell[     177] = 32'h0;  // 32'h3241d122;
    ram_cell[     178] = 32'h0;  // 32'h55a255f2;
    ram_cell[     179] = 32'h0;  // 32'h01782717;
    ram_cell[     180] = 32'h0;  // 32'h8e1de2ab;
    ram_cell[     181] = 32'h0;  // 32'hdb7021d7;
    ram_cell[     182] = 32'h0;  // 32'hc921d2b1;
    ram_cell[     183] = 32'h0;  // 32'h205ad2f5;
    ram_cell[     184] = 32'h0;  // 32'h04da7d93;
    ram_cell[     185] = 32'h0;  // 32'hb66f1ca1;
    ram_cell[     186] = 32'h0;  // 32'hae11bbdb;
    ram_cell[     187] = 32'h0;  // 32'h33730d23;
    ram_cell[     188] = 32'h0;  // 32'hde0716b5;
    ram_cell[     189] = 32'h0;  // 32'ha760a89c;
    ram_cell[     190] = 32'h0;  // 32'h0fac91bd;
    ram_cell[     191] = 32'h0;  // 32'h1a0531a1;
    ram_cell[     192] = 32'h0;  // 32'hcc94d59b;
    ram_cell[     193] = 32'h0;  // 32'h0e194f41;
    ram_cell[     194] = 32'h0;  // 32'h4cc976ef;
    ram_cell[     195] = 32'h0;  // 32'h9f9dc6ef;
    ram_cell[     196] = 32'h0;  // 32'hd328952a;
    ram_cell[     197] = 32'h0;  // 32'hc7b66eaf;
    ram_cell[     198] = 32'h0;  // 32'hd2c75a4d;
    ram_cell[     199] = 32'h0;  // 32'h0b412f9a;
    ram_cell[     200] = 32'h0;  // 32'h59924413;
    ram_cell[     201] = 32'h0;  // 32'h89c7a0d8;
    ram_cell[     202] = 32'h0;  // 32'h7460a5f4;
    ram_cell[     203] = 32'h0;  // 32'h07e54724;
    ram_cell[     204] = 32'h0;  // 32'h6ee0f1ec;
    ram_cell[     205] = 32'h0;  // 32'h250ad9eb;
    ram_cell[     206] = 32'h0;  // 32'h1db43ec4;
    ram_cell[     207] = 32'h0;  // 32'hb6dfd959;
    ram_cell[     208] = 32'h0;  // 32'h81aec487;
    ram_cell[     209] = 32'h0;  // 32'h6608db36;
    ram_cell[     210] = 32'h0;  // 32'h0dfa61f8;
    ram_cell[     211] = 32'h0;  // 32'h32091bb2;
    ram_cell[     212] = 32'h0;  // 32'ha3b156b3;
    ram_cell[     213] = 32'h0;  // 32'h8509c51c;
    ram_cell[     214] = 32'h0;  // 32'h46317a2a;
    ram_cell[     215] = 32'h0;  // 32'hdcd6c075;
    ram_cell[     216] = 32'h0;  // 32'hd1dc20ee;
    ram_cell[     217] = 32'h0;  // 32'h2f27c64f;
    ram_cell[     218] = 32'h0;  // 32'h4caa470a;
    ram_cell[     219] = 32'h0;  // 32'hf3a71d59;
    ram_cell[     220] = 32'h0;  // 32'h4c73f14d;
    ram_cell[     221] = 32'h0;  // 32'h3c6110b5;
    ram_cell[     222] = 32'h0;  // 32'ha3208d29;
    ram_cell[     223] = 32'h0;  // 32'h240a6638;
    ram_cell[     224] = 32'h0;  // 32'hb3dd631f;
    ram_cell[     225] = 32'h0;  // 32'h3fd13c1d;
    ram_cell[     226] = 32'h0;  // 32'hac21897b;
    ram_cell[     227] = 32'h0;  // 32'h225e8b02;
    ram_cell[     228] = 32'h0;  // 32'h46d8b073;
    ram_cell[     229] = 32'h0;  // 32'h191048c1;
    ram_cell[     230] = 32'h0;  // 32'he7138f12;
    ram_cell[     231] = 32'h0;  // 32'ha3aca775;
    ram_cell[     232] = 32'h0;  // 32'hab6297e6;
    ram_cell[     233] = 32'h0;  // 32'h7d0db7c2;
    ram_cell[     234] = 32'h0;  // 32'hacaa6e49;
    ram_cell[     235] = 32'h0;  // 32'h0d6fb2a2;
    ram_cell[     236] = 32'h0;  // 32'h40b901a2;
    ram_cell[     237] = 32'h0;  // 32'hf508cf7c;
    ram_cell[     238] = 32'h0;  // 32'hbc784761;
    ram_cell[     239] = 32'h0;  // 32'h8ffc740a;
    ram_cell[     240] = 32'h0;  // 32'hef17933e;
    ram_cell[     241] = 32'h0;  // 32'h25d2992a;
    ram_cell[     242] = 32'h0;  // 32'hba54c5b1;
    ram_cell[     243] = 32'h0;  // 32'he6f12db3;
    ram_cell[     244] = 32'h0;  // 32'h4933ebdd;
    ram_cell[     245] = 32'h0;  // 32'hb27acc58;
    ram_cell[     246] = 32'h0;  // 32'h65ac319a;
    ram_cell[     247] = 32'h0;  // 32'h5bafa292;
    ram_cell[     248] = 32'h0;  // 32'h0825dbfb;
    ram_cell[     249] = 32'h0;  // 32'h62d050ba;
    ram_cell[     250] = 32'h0;  // 32'he68a6297;
    ram_cell[     251] = 32'h0;  // 32'h27017d1b;
    ram_cell[     252] = 32'h0;  // 32'hbea85240;
    ram_cell[     253] = 32'h0;  // 32'h6348791f;
    ram_cell[     254] = 32'h0;  // 32'h55ab108e;
    ram_cell[     255] = 32'h0;  // 32'h342f4a2a;
    // src matrix A
    ram_cell[     256] = 32'h21d518de;
    ram_cell[     257] = 32'ha219256c;
    ram_cell[     258] = 32'hac7d5853;
    ram_cell[     259] = 32'h62820fba;
    ram_cell[     260] = 32'h74fa9c72;
    ram_cell[     261] = 32'hbe4056c2;
    ram_cell[     262] = 32'h9d48bb24;
    ram_cell[     263] = 32'h2d8d05c9;
    ram_cell[     264] = 32'h35b51ae7;
    ram_cell[     265] = 32'h087dd386;
    ram_cell[     266] = 32'hc5695d12;
    ram_cell[     267] = 32'hac0546ca;
    ram_cell[     268] = 32'hf5f652fe;
    ram_cell[     269] = 32'h27211684;
    ram_cell[     270] = 32'hb449067f;
    ram_cell[     271] = 32'ha24d9e5c;
    ram_cell[     272] = 32'hb4558db3;
    ram_cell[     273] = 32'h9aef5734;
    ram_cell[     274] = 32'h36cc25c0;
    ram_cell[     275] = 32'h650fbd4d;
    ram_cell[     276] = 32'h612addcd;
    ram_cell[     277] = 32'h16bdf3a4;
    ram_cell[     278] = 32'h7d525d95;
    ram_cell[     279] = 32'hba1ab7e2;
    ram_cell[     280] = 32'h9c3e2cc4;
    ram_cell[     281] = 32'hdddcdd4d;
    ram_cell[     282] = 32'hc793de84;
    ram_cell[     283] = 32'h7f5081dc;
    ram_cell[     284] = 32'hdd04dcb5;
    ram_cell[     285] = 32'h9e9bcc1d;
    ram_cell[     286] = 32'hf0d85b5d;
    ram_cell[     287] = 32'h484b6a73;
    ram_cell[     288] = 32'h59b64c43;
    ram_cell[     289] = 32'hf1c115f4;
    ram_cell[     290] = 32'h01840035;
    ram_cell[     291] = 32'haaa4d133;
    ram_cell[     292] = 32'h91879b3f;
    ram_cell[     293] = 32'h56487af9;
    ram_cell[     294] = 32'h1ae493fb;
    ram_cell[     295] = 32'h666531a2;
    ram_cell[     296] = 32'hb09600cb;
    ram_cell[     297] = 32'h24297d6f;
    ram_cell[     298] = 32'h4bb1f0fb;
    ram_cell[     299] = 32'hd3add05e;
    ram_cell[     300] = 32'h76de8f35;
    ram_cell[     301] = 32'h93bd9e61;
    ram_cell[     302] = 32'hc2ec4a97;
    ram_cell[     303] = 32'h60fb2f5a;
    ram_cell[     304] = 32'hc5cc26b2;
    ram_cell[     305] = 32'h3c1321b7;
    ram_cell[     306] = 32'h5d184e90;
    ram_cell[     307] = 32'hffe3cc67;
    ram_cell[     308] = 32'h202f578d;
    ram_cell[     309] = 32'ha5774283;
    ram_cell[     310] = 32'h33367d27;
    ram_cell[     311] = 32'h5efd68fe;
    ram_cell[     312] = 32'he4704784;
    ram_cell[     313] = 32'h4bf83c6e;
    ram_cell[     314] = 32'hb8a0d240;
    ram_cell[     315] = 32'h8dc4387c;
    ram_cell[     316] = 32'ha6611393;
    ram_cell[     317] = 32'h147786ea;
    ram_cell[     318] = 32'h3c2a98c5;
    ram_cell[     319] = 32'hac7b963b;
    ram_cell[     320] = 32'h33dbd8df;
    ram_cell[     321] = 32'hf178addc;
    ram_cell[     322] = 32'h50c2a633;
    ram_cell[     323] = 32'had36702c;
    ram_cell[     324] = 32'h5921f3ba;
    ram_cell[     325] = 32'h85e640f9;
    ram_cell[     326] = 32'h67c588bc;
    ram_cell[     327] = 32'hcb253c77;
    ram_cell[     328] = 32'h5be155a8;
    ram_cell[     329] = 32'h53a4f2ed;
    ram_cell[     330] = 32'h379d3ffd;
    ram_cell[     331] = 32'hbea36159;
    ram_cell[     332] = 32'ha1a7cc0b;
    ram_cell[     333] = 32'ha1b4dc27;
    ram_cell[     334] = 32'hc67dfdfe;
    ram_cell[     335] = 32'hf96686cf;
    ram_cell[     336] = 32'hf01c16b0;
    ram_cell[     337] = 32'he0e37583;
    ram_cell[     338] = 32'h19a4f6f0;
    ram_cell[     339] = 32'h44e542f0;
    ram_cell[     340] = 32'h84dbfe0c;
    ram_cell[     341] = 32'hc1f503a3;
    ram_cell[     342] = 32'h921a4b34;
    ram_cell[     343] = 32'h2af241d6;
    ram_cell[     344] = 32'h26b34545;
    ram_cell[     345] = 32'hdf74bd8d;
    ram_cell[     346] = 32'h8c65db5c;
    ram_cell[     347] = 32'h716cb571;
    ram_cell[     348] = 32'h3b366e61;
    ram_cell[     349] = 32'h08272f79;
    ram_cell[     350] = 32'hadea6066;
    ram_cell[     351] = 32'ha9bb00e5;
    ram_cell[     352] = 32'h0f4ada5f;
    ram_cell[     353] = 32'h749a8c7e;
    ram_cell[     354] = 32'h55ba312d;
    ram_cell[     355] = 32'h69cbc587;
    ram_cell[     356] = 32'h1555da82;
    ram_cell[     357] = 32'hefe80e3c;
    ram_cell[     358] = 32'he52ba588;
    ram_cell[     359] = 32'h4c54bbc9;
    ram_cell[     360] = 32'hcf6118ec;
    ram_cell[     361] = 32'h8edcf8b2;
    ram_cell[     362] = 32'hdea8e1b5;
    ram_cell[     363] = 32'hcb88cdba;
    ram_cell[     364] = 32'h4f5ca9b0;
    ram_cell[     365] = 32'he05a774d;
    ram_cell[     366] = 32'h1c8c3fb3;
    ram_cell[     367] = 32'hab85a415;
    ram_cell[     368] = 32'he5d05c71;
    ram_cell[     369] = 32'ha0686fe3;
    ram_cell[     370] = 32'h2d3eec32;
    ram_cell[     371] = 32'ha705666a;
    ram_cell[     372] = 32'h0154c69c;
    ram_cell[     373] = 32'hede20c3d;
    ram_cell[     374] = 32'h60522f42;
    ram_cell[     375] = 32'hfee8b26e;
    ram_cell[     376] = 32'hcac1e571;
    ram_cell[     377] = 32'h2321bc97;
    ram_cell[     378] = 32'hf792d35d;
    ram_cell[     379] = 32'h6332800f;
    ram_cell[     380] = 32'h342932c5;
    ram_cell[     381] = 32'h253bee5b;
    ram_cell[     382] = 32'hfd60f998;
    ram_cell[     383] = 32'hd25265a9;
    ram_cell[     384] = 32'hbe051a81;
    ram_cell[     385] = 32'h3432b2bb;
    ram_cell[     386] = 32'ha64e5df8;
    ram_cell[     387] = 32'h8b788042;
    ram_cell[     388] = 32'hedce8ce0;
    ram_cell[     389] = 32'hf2e75259;
    ram_cell[     390] = 32'h299d4cde;
    ram_cell[     391] = 32'hbc059848;
    ram_cell[     392] = 32'h8d42f4fc;
    ram_cell[     393] = 32'h0469ebc7;
    ram_cell[     394] = 32'hbe46b1d2;
    ram_cell[     395] = 32'h71bb93b3;
    ram_cell[     396] = 32'h003b0e5a;
    ram_cell[     397] = 32'hd06fe8bf;
    ram_cell[     398] = 32'he726cc44;
    ram_cell[     399] = 32'h072c97e2;
    ram_cell[     400] = 32'h8b8edc02;
    ram_cell[     401] = 32'hb96d8983;
    ram_cell[     402] = 32'hab9436a0;
    ram_cell[     403] = 32'hcd9530f2;
    ram_cell[     404] = 32'h595234e9;
    ram_cell[     405] = 32'hb4d33bb2;
    ram_cell[     406] = 32'h4de915b6;
    ram_cell[     407] = 32'h654a69a5;
    ram_cell[     408] = 32'hee5c7353;
    ram_cell[     409] = 32'h493e5940;
    ram_cell[     410] = 32'h3a3036f4;
    ram_cell[     411] = 32'h7ee72b6a;
    ram_cell[     412] = 32'hfcdcc529;
    ram_cell[     413] = 32'h02bd6dff;
    ram_cell[     414] = 32'h1ca382c9;
    ram_cell[     415] = 32'h36027a30;
    ram_cell[     416] = 32'h08ecb56f;
    ram_cell[     417] = 32'h15718f7f;
    ram_cell[     418] = 32'he9a99b4e;
    ram_cell[     419] = 32'h5c1a0fc3;
    ram_cell[     420] = 32'h7fd1ac88;
    ram_cell[     421] = 32'h2034abd9;
    ram_cell[     422] = 32'hc3cff123;
    ram_cell[     423] = 32'h354adedd;
    ram_cell[     424] = 32'hc68d5413;
    ram_cell[     425] = 32'hb3e4cc80;
    ram_cell[     426] = 32'h3c38aa03;
    ram_cell[     427] = 32'hd22fb005;
    ram_cell[     428] = 32'h99719b07;
    ram_cell[     429] = 32'h3633849d;
    ram_cell[     430] = 32'hadc30ad2;
    ram_cell[     431] = 32'h814896c8;
    ram_cell[     432] = 32'h0633fc52;
    ram_cell[     433] = 32'ha43aeef6;
    ram_cell[     434] = 32'hb00ca7f2;
    ram_cell[     435] = 32'h0f60e36c;
    ram_cell[     436] = 32'hc487f0e0;
    ram_cell[     437] = 32'hbd1a9422;
    ram_cell[     438] = 32'hebd9927e;
    ram_cell[     439] = 32'hd1e8483b;
    ram_cell[     440] = 32'ha5e6d8ab;
    ram_cell[     441] = 32'hbbcafeef;
    ram_cell[     442] = 32'h3985c706;
    ram_cell[     443] = 32'h4002ac8c;
    ram_cell[     444] = 32'h5fcd451c;
    ram_cell[     445] = 32'h3c19465f;
    ram_cell[     446] = 32'hb04e9a1e;
    ram_cell[     447] = 32'hdc63d015;
    ram_cell[     448] = 32'hc62e1203;
    ram_cell[     449] = 32'h96830346;
    ram_cell[     450] = 32'hf7dec83c;
    ram_cell[     451] = 32'hfbdb3c52;
    ram_cell[     452] = 32'h6b163d3f;
    ram_cell[     453] = 32'hc2ef45f6;
    ram_cell[     454] = 32'h6cbfdcbd;
    ram_cell[     455] = 32'h20c90ba2;
    ram_cell[     456] = 32'h0da68d15;
    ram_cell[     457] = 32'h4ac46ffe;
    ram_cell[     458] = 32'hd9a9c915;
    ram_cell[     459] = 32'hc1743b3e;
    ram_cell[     460] = 32'h272957cb;
    ram_cell[     461] = 32'h52cfcab0;
    ram_cell[     462] = 32'hd8dc5c09;
    ram_cell[     463] = 32'h5f9fb090;
    ram_cell[     464] = 32'hec35ad8e;
    ram_cell[     465] = 32'hcbdfe1db;
    ram_cell[     466] = 32'hc28aa6a3;
    ram_cell[     467] = 32'h8414e3d6;
    ram_cell[     468] = 32'he6212e10;
    ram_cell[     469] = 32'h8d92ae21;
    ram_cell[     470] = 32'h8032b6bf;
    ram_cell[     471] = 32'h2054d368;
    ram_cell[     472] = 32'hf5b5496c;
    ram_cell[     473] = 32'h51b011c4;
    ram_cell[     474] = 32'h4d881689;
    ram_cell[     475] = 32'he0215ff1;
    ram_cell[     476] = 32'h6c1c6dcb;
    ram_cell[     477] = 32'h14662bd2;
    ram_cell[     478] = 32'hf6e99e57;
    ram_cell[     479] = 32'hc56687a4;
    ram_cell[     480] = 32'h3b046772;
    ram_cell[     481] = 32'heb2c2021;
    ram_cell[     482] = 32'h68dbd890;
    ram_cell[     483] = 32'h3a0ef87b;
    ram_cell[     484] = 32'h482a7bde;
    ram_cell[     485] = 32'h90a091e9;
    ram_cell[     486] = 32'hfffe1e3c;
    ram_cell[     487] = 32'h929f4c78;
    ram_cell[     488] = 32'hdb4a2508;
    ram_cell[     489] = 32'h1fff539f;
    ram_cell[     490] = 32'h6be3a4a7;
    ram_cell[     491] = 32'hb485356e;
    ram_cell[     492] = 32'h4977f948;
    ram_cell[     493] = 32'h48c0a423;
    ram_cell[     494] = 32'h9f5a4798;
    ram_cell[     495] = 32'hbbd9dc11;
    ram_cell[     496] = 32'hdce61063;
    ram_cell[     497] = 32'ha10f7b1f;
    ram_cell[     498] = 32'h540eaeb0;
    ram_cell[     499] = 32'hba59af3f;
    ram_cell[     500] = 32'heb0cb6ef;
    ram_cell[     501] = 32'hbeac57e3;
    ram_cell[     502] = 32'h899a91aa;
    ram_cell[     503] = 32'hc13fe6f2;
    ram_cell[     504] = 32'h80ddb1c2;
    ram_cell[     505] = 32'h20d55390;
    ram_cell[     506] = 32'hf29fab62;
    ram_cell[     507] = 32'h0b760d0c;
    ram_cell[     508] = 32'h34118e2e;
    ram_cell[     509] = 32'hf1614402;
    ram_cell[     510] = 32'hab9f07e4;
    ram_cell[     511] = 32'h7eea91dc;
    // src matrix B
    ram_cell[     512] = 32'h5fbbf01c;
    ram_cell[     513] = 32'h0bab78c4;
    ram_cell[     514] = 32'h3811f14e;
    ram_cell[     515] = 32'h7e609430;
    ram_cell[     516] = 32'hb0309547;
    ram_cell[     517] = 32'h6159daaf;
    ram_cell[     518] = 32'h4d031cec;
    ram_cell[     519] = 32'hfe4471b6;
    ram_cell[     520] = 32'h83bdf8ec;
    ram_cell[     521] = 32'hb9beb45e;
    ram_cell[     522] = 32'h101851dc;
    ram_cell[     523] = 32'hdf57189a;
    ram_cell[     524] = 32'h2ed4cb35;
    ram_cell[     525] = 32'hd9e84a85;
    ram_cell[     526] = 32'h6916b1ee;
    ram_cell[     527] = 32'he0ef9e9b;
    ram_cell[     528] = 32'h99faf9fa;
    ram_cell[     529] = 32'h8789b819;
    ram_cell[     530] = 32'h764ee63c;
    ram_cell[     531] = 32'haf4a4a4f;
    ram_cell[     532] = 32'hebf47243;
    ram_cell[     533] = 32'h928813a8;
    ram_cell[     534] = 32'h5d5a5dc0;
    ram_cell[     535] = 32'hf45dc622;
    ram_cell[     536] = 32'hbdb52fd9;
    ram_cell[     537] = 32'h3faecea5;
    ram_cell[     538] = 32'h636e04ec;
    ram_cell[     539] = 32'h7be02bec;
    ram_cell[     540] = 32'h038971c5;
    ram_cell[     541] = 32'hd5aea748;
    ram_cell[     542] = 32'h16cd1e4a;
    ram_cell[     543] = 32'he943d544;
    ram_cell[     544] = 32'h5fe21b53;
    ram_cell[     545] = 32'h2e728a8f;
    ram_cell[     546] = 32'h6006e8c1;
    ram_cell[     547] = 32'h169b9ebd;
    ram_cell[     548] = 32'h41dbfd70;
    ram_cell[     549] = 32'h53e37778;
    ram_cell[     550] = 32'h1c21e157;
    ram_cell[     551] = 32'he8eae7ec;
    ram_cell[     552] = 32'h9904c714;
    ram_cell[     553] = 32'h6d57bd9f;
    ram_cell[     554] = 32'h3e162688;
    ram_cell[     555] = 32'h4b7e04e2;
    ram_cell[     556] = 32'h276fd51a;
    ram_cell[     557] = 32'hfcae19cf;
    ram_cell[     558] = 32'h6789e0e3;
    ram_cell[     559] = 32'hf7af69fa;
    ram_cell[     560] = 32'h88dbd6cb;
    ram_cell[     561] = 32'h08be7185;
    ram_cell[     562] = 32'haff1d780;
    ram_cell[     563] = 32'hd2c85637;
    ram_cell[     564] = 32'h65487dd2;
    ram_cell[     565] = 32'hbea6f851;
    ram_cell[     566] = 32'ha58bd1d6;
    ram_cell[     567] = 32'ha978fd94;
    ram_cell[     568] = 32'hd02a9680;
    ram_cell[     569] = 32'h6c03fb36;
    ram_cell[     570] = 32'h950f8e84;
    ram_cell[     571] = 32'h47d3e307;
    ram_cell[     572] = 32'hb4eb49b6;
    ram_cell[     573] = 32'h321419a9;
    ram_cell[     574] = 32'hec89ddce;
    ram_cell[     575] = 32'h982415f5;
    ram_cell[     576] = 32'hcca6ce8a;
    ram_cell[     577] = 32'he0ce81c2;
    ram_cell[     578] = 32'h62336ac8;
    ram_cell[     579] = 32'h0052989c;
    ram_cell[     580] = 32'h767b239e;
    ram_cell[     581] = 32'hc072d580;
    ram_cell[     582] = 32'h9202fc2c;
    ram_cell[     583] = 32'h37936786;
    ram_cell[     584] = 32'he8f00980;
    ram_cell[     585] = 32'hef5650ee;
    ram_cell[     586] = 32'h66cbdd0d;
    ram_cell[     587] = 32'h3de3e89e;
    ram_cell[     588] = 32'h911a6e15;
    ram_cell[     589] = 32'h8d0781a7;
    ram_cell[     590] = 32'hea41edd5;
    ram_cell[     591] = 32'h6e9cb0f1;
    ram_cell[     592] = 32'h1c7eac2f;
    ram_cell[     593] = 32'hf744f6e0;
    ram_cell[     594] = 32'h3ac1a89f;
    ram_cell[     595] = 32'h00cd253f;
    ram_cell[     596] = 32'h79d9db97;
    ram_cell[     597] = 32'h87d8b560;
    ram_cell[     598] = 32'h3ef2da54;
    ram_cell[     599] = 32'h09ed98fe;
    ram_cell[     600] = 32'h988ad956;
    ram_cell[     601] = 32'hc59c6417;
    ram_cell[     602] = 32'h96d76b0c;
    ram_cell[     603] = 32'h315d815e;
    ram_cell[     604] = 32'hec35d479;
    ram_cell[     605] = 32'h056683ca;
    ram_cell[     606] = 32'hb9cf032f;
    ram_cell[     607] = 32'h8908eced;
    ram_cell[     608] = 32'h85777c45;
    ram_cell[     609] = 32'h458e1b4c;
    ram_cell[     610] = 32'h008f6819;
    ram_cell[     611] = 32'hc3de8bc3;
    ram_cell[     612] = 32'h6585f278;
    ram_cell[     613] = 32'h9249afde;
    ram_cell[     614] = 32'hf4e8e571;
    ram_cell[     615] = 32'h19837ea3;
    ram_cell[     616] = 32'h4324e657;
    ram_cell[     617] = 32'heb19bbe7;
    ram_cell[     618] = 32'hacc8d950;
    ram_cell[     619] = 32'hcbe208f5;
    ram_cell[     620] = 32'h28065f54;
    ram_cell[     621] = 32'hf569407c;
    ram_cell[     622] = 32'he5004aed;
    ram_cell[     623] = 32'heb2a5fe8;
    ram_cell[     624] = 32'h52615f09;
    ram_cell[     625] = 32'h6cde6ecc;
    ram_cell[     626] = 32'h4e589db7;
    ram_cell[     627] = 32'he12613a6;
    ram_cell[     628] = 32'h363549ee;
    ram_cell[     629] = 32'h73bba4df;
    ram_cell[     630] = 32'heeca5b14;
    ram_cell[     631] = 32'h9c95492e;
    ram_cell[     632] = 32'h124135ab;
    ram_cell[     633] = 32'h66089e7d;
    ram_cell[     634] = 32'h76ab35a7;
    ram_cell[     635] = 32'hbe321d93;
    ram_cell[     636] = 32'hd73207b9;
    ram_cell[     637] = 32'h7814c789;
    ram_cell[     638] = 32'h62d7f37a;
    ram_cell[     639] = 32'hdf7907b6;
    ram_cell[     640] = 32'hcbea9dcd;
    ram_cell[     641] = 32'hb2589aa7;
    ram_cell[     642] = 32'h9857eee3;
    ram_cell[     643] = 32'h9ee4e5e0;
    ram_cell[     644] = 32'h03a3c2e9;
    ram_cell[     645] = 32'h90730bb0;
    ram_cell[     646] = 32'h70f491b6;
    ram_cell[     647] = 32'hc741c2a0;
    ram_cell[     648] = 32'h923a6b1e;
    ram_cell[     649] = 32'hc2e9a05a;
    ram_cell[     650] = 32'hbcb50982;
    ram_cell[     651] = 32'h53e52313;
    ram_cell[     652] = 32'h8f47bdcc;
    ram_cell[     653] = 32'hf2319bc9;
    ram_cell[     654] = 32'hf3e8b507;
    ram_cell[     655] = 32'he5f92317;
    ram_cell[     656] = 32'h9490e1fe;
    ram_cell[     657] = 32'h8ffbaa35;
    ram_cell[     658] = 32'hf18f0c1c;
    ram_cell[     659] = 32'h7b705674;
    ram_cell[     660] = 32'had218c51;
    ram_cell[     661] = 32'hb707c897;
    ram_cell[     662] = 32'h75effd2a;
    ram_cell[     663] = 32'h4126c460;
    ram_cell[     664] = 32'h7a9d8931;
    ram_cell[     665] = 32'h43dc916a;
    ram_cell[     666] = 32'hc86f5fef;
    ram_cell[     667] = 32'h00c6230f;
    ram_cell[     668] = 32'h5bcb0c1e;
    ram_cell[     669] = 32'h9cc57f15;
    ram_cell[     670] = 32'h4d8f4b91;
    ram_cell[     671] = 32'h5cde4856;
    ram_cell[     672] = 32'h9e51f254;
    ram_cell[     673] = 32'h9275e12a;
    ram_cell[     674] = 32'hda051e3e;
    ram_cell[     675] = 32'h53a6196e;
    ram_cell[     676] = 32'h767f5085;
    ram_cell[     677] = 32'h60ceebd2;
    ram_cell[     678] = 32'h0bbd69ed;
    ram_cell[     679] = 32'hffc5b3e2;
    ram_cell[     680] = 32'h58d83b43;
    ram_cell[     681] = 32'hd756a4ac;
    ram_cell[     682] = 32'h76742581;
    ram_cell[     683] = 32'he0c205f2;
    ram_cell[     684] = 32'h984822a4;
    ram_cell[     685] = 32'hb9d446f3;
    ram_cell[     686] = 32'h9c12bd3a;
    ram_cell[     687] = 32'h9095fb20;
    ram_cell[     688] = 32'h7da98613;
    ram_cell[     689] = 32'hc22acd5c;
    ram_cell[     690] = 32'hc38355bc;
    ram_cell[     691] = 32'h31ac69a6;
    ram_cell[     692] = 32'h656cc137;
    ram_cell[     693] = 32'h7753e76e;
    ram_cell[     694] = 32'h960278b2;
    ram_cell[     695] = 32'h76770183;
    ram_cell[     696] = 32'ha0358c12;
    ram_cell[     697] = 32'hd95679ea;
    ram_cell[     698] = 32'h9db9aa25;
    ram_cell[     699] = 32'ha24c1470;
    ram_cell[     700] = 32'h11805e33;
    ram_cell[     701] = 32'h2da6d3d8;
    ram_cell[     702] = 32'h997575b7;
    ram_cell[     703] = 32'h023bc217;
    ram_cell[     704] = 32'h5d2d6ea9;
    ram_cell[     705] = 32'hd7c1de6e;
    ram_cell[     706] = 32'h53510b0e;
    ram_cell[     707] = 32'h9619846c;
    ram_cell[     708] = 32'hdaaf0335;
    ram_cell[     709] = 32'hf7e1dea9;
    ram_cell[     710] = 32'h11b792e0;
    ram_cell[     711] = 32'had304a28;
    ram_cell[     712] = 32'hfed1f147;
    ram_cell[     713] = 32'h5fe7524f;
    ram_cell[     714] = 32'hb595ebda;
    ram_cell[     715] = 32'h21073295;
    ram_cell[     716] = 32'hccd1fa4b;
    ram_cell[     717] = 32'h2c01ef82;
    ram_cell[     718] = 32'hc10c6b30;
    ram_cell[     719] = 32'h5810ab21;
    ram_cell[     720] = 32'hcc7230ad;
    ram_cell[     721] = 32'h5d5d8019;
    ram_cell[     722] = 32'h7d2cea59;
    ram_cell[     723] = 32'h0e819cc4;
    ram_cell[     724] = 32'h029dedba;
    ram_cell[     725] = 32'ha01e2cb6;
    ram_cell[     726] = 32'hf3d76e36;
    ram_cell[     727] = 32'h2c7419f0;
    ram_cell[     728] = 32'hd516601e;
    ram_cell[     729] = 32'h7ed56b66;
    ram_cell[     730] = 32'h2875ae08;
    ram_cell[     731] = 32'h47c3cd21;
    ram_cell[     732] = 32'h7692cc65;
    ram_cell[     733] = 32'h9b412ab9;
    ram_cell[     734] = 32'h4a7db16f;
    ram_cell[     735] = 32'h143f11a1;
    ram_cell[     736] = 32'h8c9e8920;
    ram_cell[     737] = 32'h05ad4ee8;
    ram_cell[     738] = 32'hb7b6b189;
    ram_cell[     739] = 32'h8aebd5a4;
    ram_cell[     740] = 32'h3106a87e;
    ram_cell[     741] = 32'h50403d79;
    ram_cell[     742] = 32'h296cc2a5;
    ram_cell[     743] = 32'h1fbc8511;
    ram_cell[     744] = 32'hd05abb7c;
    ram_cell[     745] = 32'h455553be;
    ram_cell[     746] = 32'hd75123da;
    ram_cell[     747] = 32'h7567eaa1;
    ram_cell[     748] = 32'h0fbafb57;
    ram_cell[     749] = 32'h635bd27b;
    ram_cell[     750] = 32'h6e09288b;
    ram_cell[     751] = 32'h7977ce89;
    ram_cell[     752] = 32'h97337486;
    ram_cell[     753] = 32'hbc238415;
    ram_cell[     754] = 32'ha0378a61;
    ram_cell[     755] = 32'h6d9f98c5;
    ram_cell[     756] = 32'h5678a6dd;
    ram_cell[     757] = 32'h082ec0eb;
    ram_cell[     758] = 32'h93db2cf3;
    ram_cell[     759] = 32'hfd7b0687;
    ram_cell[     760] = 32'h4f54cb4f;
    ram_cell[     761] = 32'ha205f38c;
    ram_cell[     762] = 32'h7d8b0549;
    ram_cell[     763] = 32'h1f07837f;
    ram_cell[     764] = 32'h757970a3;
    ram_cell[     765] = 32'h2209c0e2;
    ram_cell[     766] = 32'h38b38e3a;
    ram_cell[     767] = 32'hcd37726d;
end

endmodule



module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hbd904917;
    ram_cell[       1] = 32'h0;  // 32'h19aecacd;
    ram_cell[       2] = 32'h0;  // 32'h7d008984;
    ram_cell[       3] = 32'h0;  // 32'hdc0440b1;
    ram_cell[       4] = 32'h0;  // 32'hd36ea304;
    ram_cell[       5] = 32'h0;  // 32'hdd41afdc;
    ram_cell[       6] = 32'h0;  // 32'hdb546741;
    ram_cell[       7] = 32'h0;  // 32'h8c70a6bc;
    ram_cell[       8] = 32'h0;  // 32'hc2f4c773;
    ram_cell[       9] = 32'h0;  // 32'hbbef7037;
    ram_cell[      10] = 32'h0;  // 32'h171d35c1;
    ram_cell[      11] = 32'h0;  // 32'hd5a8a5b0;
    ram_cell[      12] = 32'h0;  // 32'hf929d4b2;
    ram_cell[      13] = 32'h0;  // 32'h8747aaaf;
    ram_cell[      14] = 32'h0;  // 32'h11bdfb4e;
    ram_cell[      15] = 32'h0;  // 32'h9fed4d78;
    ram_cell[      16] = 32'h0;  // 32'h09be9639;
    ram_cell[      17] = 32'h0;  // 32'ha96fcfe4;
    ram_cell[      18] = 32'h0;  // 32'hb9411eca;
    ram_cell[      19] = 32'h0;  // 32'h710fc696;
    ram_cell[      20] = 32'h0;  // 32'hcc883696;
    ram_cell[      21] = 32'h0;  // 32'hb7a6eac8;
    ram_cell[      22] = 32'h0;  // 32'h4fdd2ccc;
    ram_cell[      23] = 32'h0;  // 32'hc48e47b1;
    ram_cell[      24] = 32'h0;  // 32'h5f8c6129;
    ram_cell[      25] = 32'h0;  // 32'h2eb333fc;
    ram_cell[      26] = 32'h0;  // 32'hfc1a38ff;
    ram_cell[      27] = 32'h0;  // 32'h709d7437;
    ram_cell[      28] = 32'h0;  // 32'h9b7b9537;
    ram_cell[      29] = 32'h0;  // 32'h51749dc7;
    ram_cell[      30] = 32'h0;  // 32'h7ec08709;
    ram_cell[      31] = 32'h0;  // 32'hb366895a;
    ram_cell[      32] = 32'h0;  // 32'h3bf2f015;
    ram_cell[      33] = 32'h0;  // 32'h45a9ec9d;
    ram_cell[      34] = 32'h0;  // 32'h72078a54;
    ram_cell[      35] = 32'h0;  // 32'h7071132d;
    ram_cell[      36] = 32'h0;  // 32'h4d02a478;
    ram_cell[      37] = 32'h0;  // 32'h4596ee01;
    ram_cell[      38] = 32'h0;  // 32'h3112c359;
    ram_cell[      39] = 32'h0;  // 32'he4d3c57a;
    ram_cell[      40] = 32'h0;  // 32'hf312905c;
    ram_cell[      41] = 32'h0;  // 32'h310fd820;
    ram_cell[      42] = 32'h0;  // 32'hafdcb01a;
    ram_cell[      43] = 32'h0;  // 32'hd3e71cdc;
    ram_cell[      44] = 32'h0;  // 32'h8c716485;
    ram_cell[      45] = 32'h0;  // 32'h26655846;
    ram_cell[      46] = 32'h0;  // 32'hfc250d43;
    ram_cell[      47] = 32'h0;  // 32'heca900b5;
    ram_cell[      48] = 32'h0;  // 32'h6c80410c;
    ram_cell[      49] = 32'h0;  // 32'h24fd10ef;
    ram_cell[      50] = 32'h0;  // 32'h9cf7b2df;
    ram_cell[      51] = 32'h0;  // 32'he0ebf6fa;
    ram_cell[      52] = 32'h0;  // 32'hd61534c5;
    ram_cell[      53] = 32'h0;  // 32'hfc92a19c;
    ram_cell[      54] = 32'h0;  // 32'hdca076cc;
    ram_cell[      55] = 32'h0;  // 32'h40253348;
    ram_cell[      56] = 32'h0;  // 32'hb91063f1;
    ram_cell[      57] = 32'h0;  // 32'ha426eb49;
    ram_cell[      58] = 32'h0;  // 32'h068881f0;
    ram_cell[      59] = 32'h0;  // 32'h9832cd64;
    ram_cell[      60] = 32'h0;  // 32'h90af2f72;
    ram_cell[      61] = 32'h0;  // 32'h75e9dc11;
    ram_cell[      62] = 32'h0;  // 32'h206323ea;
    ram_cell[      63] = 32'h0;  // 32'hff9dfaf3;
    ram_cell[      64] = 32'h0;  // 32'h5c975d00;
    ram_cell[      65] = 32'h0;  // 32'h96252782;
    ram_cell[      66] = 32'h0;  // 32'h754b01ae;
    ram_cell[      67] = 32'h0;  // 32'hf3681a9f;
    ram_cell[      68] = 32'h0;  // 32'h59dddb87;
    ram_cell[      69] = 32'h0;  // 32'hd6549ce9;
    ram_cell[      70] = 32'h0;  // 32'h6b1eb949;
    ram_cell[      71] = 32'h0;  // 32'ha5c62f8f;
    ram_cell[      72] = 32'h0;  // 32'h9adf970c;
    ram_cell[      73] = 32'h0;  // 32'h87e56ae6;
    ram_cell[      74] = 32'h0;  // 32'h03454804;
    ram_cell[      75] = 32'h0;  // 32'hd53561a6;
    ram_cell[      76] = 32'h0;  // 32'h6175fc19;
    ram_cell[      77] = 32'h0;  // 32'h46be90ce;
    ram_cell[      78] = 32'h0;  // 32'h07926dff;
    ram_cell[      79] = 32'h0;  // 32'h67c8821c;
    ram_cell[      80] = 32'h0;  // 32'hbc37df5b;
    ram_cell[      81] = 32'h0;  // 32'h2b5479f7;
    ram_cell[      82] = 32'h0;  // 32'h33e3d64e;
    ram_cell[      83] = 32'h0;  // 32'h74e3ef02;
    ram_cell[      84] = 32'h0;  // 32'h646147dd;
    ram_cell[      85] = 32'h0;  // 32'h6a43ead3;
    ram_cell[      86] = 32'h0;  // 32'h5244a722;
    ram_cell[      87] = 32'h0;  // 32'h2f58be6f;
    ram_cell[      88] = 32'h0;  // 32'h3715a15e;
    ram_cell[      89] = 32'h0;  // 32'h3813c025;
    ram_cell[      90] = 32'h0;  // 32'h7868cab5;
    ram_cell[      91] = 32'h0;  // 32'h040b4597;
    ram_cell[      92] = 32'h0;  // 32'hba89b1f6;
    ram_cell[      93] = 32'h0;  // 32'hb2fb070e;
    ram_cell[      94] = 32'h0;  // 32'h7696d7a1;
    ram_cell[      95] = 32'h0;  // 32'h5070f145;
    ram_cell[      96] = 32'h0;  // 32'h9d9e1ce3;
    ram_cell[      97] = 32'h0;  // 32'h9d4a0205;
    ram_cell[      98] = 32'h0;  // 32'h81a8cdc3;
    ram_cell[      99] = 32'h0;  // 32'h02fbbb2f;
    ram_cell[     100] = 32'h0;  // 32'h031b754d;
    ram_cell[     101] = 32'h0;  // 32'haf26e8ea;
    ram_cell[     102] = 32'h0;  // 32'hbf853ae7;
    ram_cell[     103] = 32'h0;  // 32'hdd6ff083;
    ram_cell[     104] = 32'h0;  // 32'h9c65bbf3;
    ram_cell[     105] = 32'h0;  // 32'h4708508e;
    ram_cell[     106] = 32'h0;  // 32'h841d86ea;
    ram_cell[     107] = 32'h0;  // 32'hc33e25a8;
    ram_cell[     108] = 32'h0;  // 32'hc756aa6e;
    ram_cell[     109] = 32'h0;  // 32'he42de840;
    ram_cell[     110] = 32'h0;  // 32'hfe56ff3f;
    ram_cell[     111] = 32'h0;  // 32'h14aeee4b;
    ram_cell[     112] = 32'h0;  // 32'ha1be27f1;
    ram_cell[     113] = 32'h0;  // 32'hc73e6516;
    ram_cell[     114] = 32'h0;  // 32'h9f443d9a;
    ram_cell[     115] = 32'h0;  // 32'hfbf5c5cd;
    ram_cell[     116] = 32'h0;  // 32'ha4d710cd;
    ram_cell[     117] = 32'h0;  // 32'h516beabc;
    ram_cell[     118] = 32'h0;  // 32'h664fece4;
    ram_cell[     119] = 32'h0;  // 32'hfde73a57;
    ram_cell[     120] = 32'h0;  // 32'h1f818e9a;
    ram_cell[     121] = 32'h0;  // 32'he0af8a62;
    ram_cell[     122] = 32'h0;  // 32'hb9971541;
    ram_cell[     123] = 32'h0;  // 32'hb97c420e;
    ram_cell[     124] = 32'h0;  // 32'h077ecacc;
    ram_cell[     125] = 32'h0;  // 32'ha434d8a6;
    ram_cell[     126] = 32'h0;  // 32'h7ae4427e;
    ram_cell[     127] = 32'h0;  // 32'h66d69f5d;
    ram_cell[     128] = 32'h0;  // 32'hcd3bd3a9;
    ram_cell[     129] = 32'h0;  // 32'h35d74cfe;
    ram_cell[     130] = 32'h0;  // 32'h189a81a5;
    ram_cell[     131] = 32'h0;  // 32'h80cbb290;
    ram_cell[     132] = 32'h0;  // 32'h09d12b35;
    ram_cell[     133] = 32'h0;  // 32'h6c43d78d;
    ram_cell[     134] = 32'h0;  // 32'h28935df3;
    ram_cell[     135] = 32'h0;  // 32'he6641117;
    ram_cell[     136] = 32'h0;  // 32'hefea855e;
    ram_cell[     137] = 32'h0;  // 32'h01b23062;
    ram_cell[     138] = 32'h0;  // 32'h9206fa2d;
    ram_cell[     139] = 32'h0;  // 32'hed70eb3f;
    ram_cell[     140] = 32'h0;  // 32'h5f00f67a;
    ram_cell[     141] = 32'h0;  // 32'h93c8b189;
    ram_cell[     142] = 32'h0;  // 32'h9842af5c;
    ram_cell[     143] = 32'h0;  // 32'hf45e5f8b;
    ram_cell[     144] = 32'h0;  // 32'h9c612ac7;
    ram_cell[     145] = 32'h0;  // 32'h595f800d;
    ram_cell[     146] = 32'h0;  // 32'hbe44ae02;
    ram_cell[     147] = 32'h0;  // 32'h37cf5cd8;
    ram_cell[     148] = 32'h0;  // 32'heda0b80a;
    ram_cell[     149] = 32'h0;  // 32'ha1d1384c;
    ram_cell[     150] = 32'h0;  // 32'hcc04294a;
    ram_cell[     151] = 32'h0;  // 32'h0202b6a1;
    ram_cell[     152] = 32'h0;  // 32'h28cefc60;
    ram_cell[     153] = 32'h0;  // 32'hedb8463e;
    ram_cell[     154] = 32'h0;  // 32'hc1cce7cc;
    ram_cell[     155] = 32'h0;  // 32'hd276e95e;
    ram_cell[     156] = 32'h0;  // 32'h87bd964c;
    ram_cell[     157] = 32'h0;  // 32'h5363987c;
    ram_cell[     158] = 32'h0;  // 32'h42544160;
    ram_cell[     159] = 32'h0;  // 32'hdd1db0d8;
    ram_cell[     160] = 32'h0;  // 32'h4a4dc84d;
    ram_cell[     161] = 32'h0;  // 32'h06d20044;
    ram_cell[     162] = 32'h0;  // 32'h7e8c19b9;
    ram_cell[     163] = 32'h0;  // 32'h556119d4;
    ram_cell[     164] = 32'h0;  // 32'h67843780;
    ram_cell[     165] = 32'h0;  // 32'h1fb6ec12;
    ram_cell[     166] = 32'h0;  // 32'ha78d4201;
    ram_cell[     167] = 32'h0;  // 32'h2b5f826a;
    ram_cell[     168] = 32'h0;  // 32'h5af9c2f8;
    ram_cell[     169] = 32'h0;  // 32'h557ef739;
    ram_cell[     170] = 32'h0;  // 32'h332115fd;
    ram_cell[     171] = 32'h0;  // 32'h0d96e67e;
    ram_cell[     172] = 32'h0;  // 32'h1c908565;
    ram_cell[     173] = 32'h0;  // 32'h16651975;
    ram_cell[     174] = 32'h0;  // 32'hd5603837;
    ram_cell[     175] = 32'h0;  // 32'h7c5ff0b0;
    ram_cell[     176] = 32'h0;  // 32'h341eaabf;
    ram_cell[     177] = 32'h0;  // 32'h43455512;
    ram_cell[     178] = 32'h0;  // 32'h6b3fafbd;
    ram_cell[     179] = 32'h0;  // 32'h48162d5a;
    ram_cell[     180] = 32'h0;  // 32'h53c5cce1;
    ram_cell[     181] = 32'h0;  // 32'h932084d4;
    ram_cell[     182] = 32'h0;  // 32'he18ea043;
    ram_cell[     183] = 32'h0;  // 32'he0c06f02;
    ram_cell[     184] = 32'h0;  // 32'hf54dbe85;
    ram_cell[     185] = 32'h0;  // 32'he7ef9b5e;
    ram_cell[     186] = 32'h0;  // 32'hae6eaea8;
    ram_cell[     187] = 32'h0;  // 32'hfa4ceb2b;
    ram_cell[     188] = 32'h0;  // 32'h11bc5040;
    ram_cell[     189] = 32'h0;  // 32'h77cd53f3;
    ram_cell[     190] = 32'h0;  // 32'h6e1f543f;
    ram_cell[     191] = 32'h0;  // 32'hda033465;
    ram_cell[     192] = 32'h0;  // 32'hbdc34140;
    ram_cell[     193] = 32'h0;  // 32'hd4c6d9cb;
    ram_cell[     194] = 32'h0;  // 32'h4acbfdcf;
    ram_cell[     195] = 32'h0;  // 32'h551fab9d;
    ram_cell[     196] = 32'h0;  // 32'h057c15a5;
    ram_cell[     197] = 32'h0;  // 32'h75af4c01;
    ram_cell[     198] = 32'h0;  // 32'h11f0fd60;
    ram_cell[     199] = 32'h0;  // 32'h4878750c;
    ram_cell[     200] = 32'h0;  // 32'hda4ef6a9;
    ram_cell[     201] = 32'h0;  // 32'h85941eaa;
    ram_cell[     202] = 32'h0;  // 32'h99c4ecf5;
    ram_cell[     203] = 32'h0;  // 32'ha9545264;
    ram_cell[     204] = 32'h0;  // 32'h371a825e;
    ram_cell[     205] = 32'h0;  // 32'h4564f97b;
    ram_cell[     206] = 32'h0;  // 32'h6f37644c;
    ram_cell[     207] = 32'h0;  // 32'h3b28cf34;
    ram_cell[     208] = 32'h0;  // 32'hcb8da98d;
    ram_cell[     209] = 32'h0;  // 32'h8f45d597;
    ram_cell[     210] = 32'h0;  // 32'h1d5184c2;
    ram_cell[     211] = 32'h0;  // 32'h2bc80f82;
    ram_cell[     212] = 32'h0;  // 32'h58fe0751;
    ram_cell[     213] = 32'h0;  // 32'h8b531a12;
    ram_cell[     214] = 32'h0;  // 32'h79ec1b3e;
    ram_cell[     215] = 32'h0;  // 32'h8f6e81d9;
    ram_cell[     216] = 32'h0;  // 32'h406a1258;
    ram_cell[     217] = 32'h0;  // 32'hc34a25fd;
    ram_cell[     218] = 32'h0;  // 32'hccf51ca9;
    ram_cell[     219] = 32'h0;  // 32'hf2054454;
    ram_cell[     220] = 32'h0;  // 32'h413af00c;
    ram_cell[     221] = 32'h0;  // 32'he1cc52c9;
    ram_cell[     222] = 32'h0;  // 32'h01e29388;
    ram_cell[     223] = 32'h0;  // 32'hc196cc2e;
    ram_cell[     224] = 32'h0;  // 32'h1f8abc91;
    ram_cell[     225] = 32'h0;  // 32'hc12cdd5e;
    ram_cell[     226] = 32'h0;  // 32'h0739e4fd;
    ram_cell[     227] = 32'h0;  // 32'h766d11e1;
    ram_cell[     228] = 32'h0;  // 32'he99b809a;
    ram_cell[     229] = 32'h0;  // 32'ha1821e3d;
    ram_cell[     230] = 32'h0;  // 32'hc9e76c52;
    ram_cell[     231] = 32'h0;  // 32'h39ba8f70;
    ram_cell[     232] = 32'h0;  // 32'hfe43efc6;
    ram_cell[     233] = 32'h0;  // 32'h85da41b7;
    ram_cell[     234] = 32'h0;  // 32'h81249707;
    ram_cell[     235] = 32'h0;  // 32'hbcc1b685;
    ram_cell[     236] = 32'h0;  // 32'hb602e9c9;
    ram_cell[     237] = 32'h0;  // 32'hf330d932;
    ram_cell[     238] = 32'h0;  // 32'hfd154019;
    ram_cell[     239] = 32'h0;  // 32'h4de964cb;
    ram_cell[     240] = 32'h0;  // 32'h9befe9b5;
    ram_cell[     241] = 32'h0;  // 32'h0cf43dc8;
    ram_cell[     242] = 32'h0;  // 32'hccdcbc57;
    ram_cell[     243] = 32'h0;  // 32'h84524fef;
    ram_cell[     244] = 32'h0;  // 32'h8356a485;
    ram_cell[     245] = 32'h0;  // 32'h815b5903;
    ram_cell[     246] = 32'h0;  // 32'h84bc9458;
    ram_cell[     247] = 32'h0;  // 32'hf4e46303;
    ram_cell[     248] = 32'h0;  // 32'hb3070f04;
    ram_cell[     249] = 32'h0;  // 32'hfeff4acd;
    ram_cell[     250] = 32'h0;  // 32'hf3542f7a;
    ram_cell[     251] = 32'h0;  // 32'h2b5af4be;
    ram_cell[     252] = 32'h0;  // 32'h37834c28;
    ram_cell[     253] = 32'h0;  // 32'h988b0986;
    ram_cell[     254] = 32'h0;  // 32'h751e4aa7;
    ram_cell[     255] = 32'h0;  // 32'hfb785470;
    // src matrix A
    ram_cell[     256] = 32'h56ed3902;
    ram_cell[     257] = 32'h09bd026b;
    ram_cell[     258] = 32'h8d94526d;
    ram_cell[     259] = 32'h7eee3348;
    ram_cell[     260] = 32'h36dbb5f2;
    ram_cell[     261] = 32'hc912e842;
    ram_cell[     262] = 32'h0b258f13;
    ram_cell[     263] = 32'h31b566e0;
    ram_cell[     264] = 32'hdd734b93;
    ram_cell[     265] = 32'h637ea145;
    ram_cell[     266] = 32'h044ca337;
    ram_cell[     267] = 32'h9fd0582e;
    ram_cell[     268] = 32'hd54da416;
    ram_cell[     269] = 32'h133edc14;
    ram_cell[     270] = 32'h27b4ae58;
    ram_cell[     271] = 32'haee18127;
    ram_cell[     272] = 32'h6e894de4;
    ram_cell[     273] = 32'he568e5aa;
    ram_cell[     274] = 32'h5e9e1e28;
    ram_cell[     275] = 32'h12debf6a;
    ram_cell[     276] = 32'h2d6dee68;
    ram_cell[     277] = 32'hb8fa1a38;
    ram_cell[     278] = 32'h2fb3126c;
    ram_cell[     279] = 32'hcb0aaa25;
    ram_cell[     280] = 32'hcec63764;
    ram_cell[     281] = 32'h89f1b206;
    ram_cell[     282] = 32'hbed26096;
    ram_cell[     283] = 32'hb98bcc7c;
    ram_cell[     284] = 32'hca6f0ade;
    ram_cell[     285] = 32'h997be185;
    ram_cell[     286] = 32'h33ff427f;
    ram_cell[     287] = 32'ha335445b;
    ram_cell[     288] = 32'h041d3702;
    ram_cell[     289] = 32'h9cbc422c;
    ram_cell[     290] = 32'h8630fa4d;
    ram_cell[     291] = 32'h4c45cd54;
    ram_cell[     292] = 32'hfc83063c;
    ram_cell[     293] = 32'hfbb8577d;
    ram_cell[     294] = 32'h49eb62d8;
    ram_cell[     295] = 32'h88a2009b;
    ram_cell[     296] = 32'h79f057ee;
    ram_cell[     297] = 32'h8867f464;
    ram_cell[     298] = 32'h39b75879;
    ram_cell[     299] = 32'h072fd1ed;
    ram_cell[     300] = 32'he4c0acf4;
    ram_cell[     301] = 32'h0190af05;
    ram_cell[     302] = 32'hc5551d02;
    ram_cell[     303] = 32'hd9023f37;
    ram_cell[     304] = 32'h74e17fb6;
    ram_cell[     305] = 32'h21ed31b3;
    ram_cell[     306] = 32'h823d6931;
    ram_cell[     307] = 32'he38c153c;
    ram_cell[     308] = 32'h354b7d69;
    ram_cell[     309] = 32'hb1718b15;
    ram_cell[     310] = 32'h3b069471;
    ram_cell[     311] = 32'hc086414a;
    ram_cell[     312] = 32'he6d57efb;
    ram_cell[     313] = 32'h2ec9ce06;
    ram_cell[     314] = 32'h083130f4;
    ram_cell[     315] = 32'h86432488;
    ram_cell[     316] = 32'hf788d848;
    ram_cell[     317] = 32'hbe76b299;
    ram_cell[     318] = 32'h6a018afa;
    ram_cell[     319] = 32'h27b2c28a;
    ram_cell[     320] = 32'h920f43b9;
    ram_cell[     321] = 32'h11e69126;
    ram_cell[     322] = 32'h48a1cd18;
    ram_cell[     323] = 32'h3dd9fc97;
    ram_cell[     324] = 32'hc0803384;
    ram_cell[     325] = 32'h12fff820;
    ram_cell[     326] = 32'h22a39c2d;
    ram_cell[     327] = 32'hc5d25377;
    ram_cell[     328] = 32'h111c6993;
    ram_cell[     329] = 32'h8a9e37c3;
    ram_cell[     330] = 32'h4d304847;
    ram_cell[     331] = 32'hd834176e;
    ram_cell[     332] = 32'h2322a5cb;
    ram_cell[     333] = 32'h5792f7ef;
    ram_cell[     334] = 32'h27c8de38;
    ram_cell[     335] = 32'hc2154d9c;
    ram_cell[     336] = 32'h2f716952;
    ram_cell[     337] = 32'hbb63818f;
    ram_cell[     338] = 32'hbb73add8;
    ram_cell[     339] = 32'h89effcf3;
    ram_cell[     340] = 32'h413a16d8;
    ram_cell[     341] = 32'h46435433;
    ram_cell[     342] = 32'hd76eff69;
    ram_cell[     343] = 32'hd3075515;
    ram_cell[     344] = 32'h1d124fed;
    ram_cell[     345] = 32'ha46e16ed;
    ram_cell[     346] = 32'hc7953cec;
    ram_cell[     347] = 32'hfa47334f;
    ram_cell[     348] = 32'h78e4a488;
    ram_cell[     349] = 32'h0145daac;
    ram_cell[     350] = 32'h4a74cb6c;
    ram_cell[     351] = 32'h566ce82f;
    ram_cell[     352] = 32'h1dd0486c;
    ram_cell[     353] = 32'h4f635d51;
    ram_cell[     354] = 32'h33e767cb;
    ram_cell[     355] = 32'hd8bac320;
    ram_cell[     356] = 32'hb5483794;
    ram_cell[     357] = 32'h7818567b;
    ram_cell[     358] = 32'h5812ecec;
    ram_cell[     359] = 32'hf811c76c;
    ram_cell[     360] = 32'h4dfd371d;
    ram_cell[     361] = 32'hfe4430e5;
    ram_cell[     362] = 32'hd0f15a6d;
    ram_cell[     363] = 32'h3b7a5a4e;
    ram_cell[     364] = 32'h0468663d;
    ram_cell[     365] = 32'h9a280d0d;
    ram_cell[     366] = 32'he627c9a7;
    ram_cell[     367] = 32'h8ac5f9bc;
    ram_cell[     368] = 32'h5d11395a;
    ram_cell[     369] = 32'ha1e5e3d0;
    ram_cell[     370] = 32'hf988102c;
    ram_cell[     371] = 32'hd9fbf322;
    ram_cell[     372] = 32'h8f45aa34;
    ram_cell[     373] = 32'hce66d0a1;
    ram_cell[     374] = 32'h703197c9;
    ram_cell[     375] = 32'hd51fb5b7;
    ram_cell[     376] = 32'ha5a73bfb;
    ram_cell[     377] = 32'h1f39deda;
    ram_cell[     378] = 32'h009f7d61;
    ram_cell[     379] = 32'hd80c47ef;
    ram_cell[     380] = 32'h6cfaa0cb;
    ram_cell[     381] = 32'h8d23d263;
    ram_cell[     382] = 32'h2d33ac27;
    ram_cell[     383] = 32'h44ade53d;
    ram_cell[     384] = 32'h70a52fa8;
    ram_cell[     385] = 32'hfcbf5923;
    ram_cell[     386] = 32'ha9744236;
    ram_cell[     387] = 32'h85d9dfd7;
    ram_cell[     388] = 32'h48a5295b;
    ram_cell[     389] = 32'h1217fe09;
    ram_cell[     390] = 32'h7b50e7ea;
    ram_cell[     391] = 32'hb55210a5;
    ram_cell[     392] = 32'hfd931c4b;
    ram_cell[     393] = 32'h14022303;
    ram_cell[     394] = 32'h4081a762;
    ram_cell[     395] = 32'h882e78dd;
    ram_cell[     396] = 32'h53aec270;
    ram_cell[     397] = 32'h5a517361;
    ram_cell[     398] = 32'h6dcfc27f;
    ram_cell[     399] = 32'hee7847f4;
    ram_cell[     400] = 32'h6523d120;
    ram_cell[     401] = 32'h25d80693;
    ram_cell[     402] = 32'hdfaa0e21;
    ram_cell[     403] = 32'hf1d1e596;
    ram_cell[     404] = 32'h85717e74;
    ram_cell[     405] = 32'h8e346b0d;
    ram_cell[     406] = 32'h80aa9917;
    ram_cell[     407] = 32'heeb0066c;
    ram_cell[     408] = 32'hf39654ae;
    ram_cell[     409] = 32'h99ebaa63;
    ram_cell[     410] = 32'h685b6033;
    ram_cell[     411] = 32'hcd874149;
    ram_cell[     412] = 32'h2d2abdc3;
    ram_cell[     413] = 32'ha7d211b4;
    ram_cell[     414] = 32'h1ca1ea74;
    ram_cell[     415] = 32'hbe9d76a3;
    ram_cell[     416] = 32'hf41cdf02;
    ram_cell[     417] = 32'h1abed6ad;
    ram_cell[     418] = 32'hc74b0331;
    ram_cell[     419] = 32'hbf6d7038;
    ram_cell[     420] = 32'hdb2b3f60;
    ram_cell[     421] = 32'h9b92f237;
    ram_cell[     422] = 32'h1211df19;
    ram_cell[     423] = 32'hf31a1a86;
    ram_cell[     424] = 32'hf94367d8;
    ram_cell[     425] = 32'h893a34fa;
    ram_cell[     426] = 32'h43dc53e1;
    ram_cell[     427] = 32'h491a5f27;
    ram_cell[     428] = 32'h568d106b;
    ram_cell[     429] = 32'hd72269e4;
    ram_cell[     430] = 32'h7de2ac85;
    ram_cell[     431] = 32'hca8fa7c3;
    ram_cell[     432] = 32'h37a94bb1;
    ram_cell[     433] = 32'hc6f6a2b3;
    ram_cell[     434] = 32'ha9e7d47b;
    ram_cell[     435] = 32'h471f2307;
    ram_cell[     436] = 32'h8fb45631;
    ram_cell[     437] = 32'h5ab0b11c;
    ram_cell[     438] = 32'hb7648e82;
    ram_cell[     439] = 32'h63c25ff8;
    ram_cell[     440] = 32'h52515f99;
    ram_cell[     441] = 32'h40f44fe8;
    ram_cell[     442] = 32'h5442a3fb;
    ram_cell[     443] = 32'hdc120c45;
    ram_cell[     444] = 32'h8320d2b9;
    ram_cell[     445] = 32'h79eac29c;
    ram_cell[     446] = 32'h9e2d618b;
    ram_cell[     447] = 32'hc4265ba0;
    ram_cell[     448] = 32'h6b7e2c15;
    ram_cell[     449] = 32'h28d566f7;
    ram_cell[     450] = 32'h9b05f172;
    ram_cell[     451] = 32'hd5ba8b1b;
    ram_cell[     452] = 32'h53d70893;
    ram_cell[     453] = 32'h4267fff3;
    ram_cell[     454] = 32'hdfc47f91;
    ram_cell[     455] = 32'h7b4c565d;
    ram_cell[     456] = 32'h9d0b6a29;
    ram_cell[     457] = 32'h1d94b7ed;
    ram_cell[     458] = 32'h17efdc29;
    ram_cell[     459] = 32'h2fa80708;
    ram_cell[     460] = 32'h34448739;
    ram_cell[     461] = 32'h26d7f2ae;
    ram_cell[     462] = 32'hf34bdd1a;
    ram_cell[     463] = 32'h107b0aba;
    ram_cell[     464] = 32'hf6477f9f;
    ram_cell[     465] = 32'h82c65f6d;
    ram_cell[     466] = 32'hea9dba55;
    ram_cell[     467] = 32'h47c3d77b;
    ram_cell[     468] = 32'hb652efdc;
    ram_cell[     469] = 32'h476cceca;
    ram_cell[     470] = 32'h8986c412;
    ram_cell[     471] = 32'h6c6df2fb;
    ram_cell[     472] = 32'h68209b72;
    ram_cell[     473] = 32'hb1e4fbdf;
    ram_cell[     474] = 32'he0069f8c;
    ram_cell[     475] = 32'hfe97625e;
    ram_cell[     476] = 32'h8204197a;
    ram_cell[     477] = 32'h6a9ef2d2;
    ram_cell[     478] = 32'h54bced03;
    ram_cell[     479] = 32'h9f09a2d7;
    ram_cell[     480] = 32'h27261062;
    ram_cell[     481] = 32'h183e2ebe;
    ram_cell[     482] = 32'h5d10e821;
    ram_cell[     483] = 32'ha4fca673;
    ram_cell[     484] = 32'he78c0669;
    ram_cell[     485] = 32'h7d827e83;
    ram_cell[     486] = 32'hcb0f65b7;
    ram_cell[     487] = 32'hd938247f;
    ram_cell[     488] = 32'h3c44a482;
    ram_cell[     489] = 32'h3c4e09be;
    ram_cell[     490] = 32'h5c7f0ab1;
    ram_cell[     491] = 32'h95dfd1d6;
    ram_cell[     492] = 32'hec05920a;
    ram_cell[     493] = 32'hc14484c6;
    ram_cell[     494] = 32'h17ff358f;
    ram_cell[     495] = 32'he776d6b5;
    ram_cell[     496] = 32'h41f3df14;
    ram_cell[     497] = 32'h4bc83455;
    ram_cell[     498] = 32'h5bb40275;
    ram_cell[     499] = 32'h330cf37c;
    ram_cell[     500] = 32'h71044e15;
    ram_cell[     501] = 32'ha225805e;
    ram_cell[     502] = 32'h29dcde3f;
    ram_cell[     503] = 32'hbe05065c;
    ram_cell[     504] = 32'h34e1ec04;
    ram_cell[     505] = 32'h6cbf942e;
    ram_cell[     506] = 32'h590e42aa;
    ram_cell[     507] = 32'ha2288732;
    ram_cell[     508] = 32'he6ffdf70;
    ram_cell[     509] = 32'h6e154476;
    ram_cell[     510] = 32'h25c2a366;
    ram_cell[     511] = 32'h663111f7;
    // src matrix B
    ram_cell[     512] = 32'hf71eecfc;
    ram_cell[     513] = 32'h8f0e2daf;
    ram_cell[     514] = 32'h896e02b4;
    ram_cell[     515] = 32'h9efad6f3;
    ram_cell[     516] = 32'hb7cd90be;
    ram_cell[     517] = 32'hfb3250e7;
    ram_cell[     518] = 32'h27bf334a;
    ram_cell[     519] = 32'hbddf275d;
    ram_cell[     520] = 32'h63a5417e;
    ram_cell[     521] = 32'h38100c5e;
    ram_cell[     522] = 32'h396b3f5a;
    ram_cell[     523] = 32'h10832964;
    ram_cell[     524] = 32'hafc13b9e;
    ram_cell[     525] = 32'h90619dbe;
    ram_cell[     526] = 32'h87fac01c;
    ram_cell[     527] = 32'h622c7073;
    ram_cell[     528] = 32'h54d196ca;
    ram_cell[     529] = 32'h8a710b0b;
    ram_cell[     530] = 32'h9731c242;
    ram_cell[     531] = 32'h7c7274a6;
    ram_cell[     532] = 32'h2d14c469;
    ram_cell[     533] = 32'h67c33f05;
    ram_cell[     534] = 32'ha4b3eb95;
    ram_cell[     535] = 32'h473bc563;
    ram_cell[     536] = 32'hd5a921a0;
    ram_cell[     537] = 32'he94afbaf;
    ram_cell[     538] = 32'h689a5189;
    ram_cell[     539] = 32'h93317d3a;
    ram_cell[     540] = 32'he1a82bdb;
    ram_cell[     541] = 32'haf110d32;
    ram_cell[     542] = 32'h07ebd549;
    ram_cell[     543] = 32'h6d4555f1;
    ram_cell[     544] = 32'he605ede9;
    ram_cell[     545] = 32'h01cda4b0;
    ram_cell[     546] = 32'h066b3c83;
    ram_cell[     547] = 32'hb82fd849;
    ram_cell[     548] = 32'hdae5afa4;
    ram_cell[     549] = 32'h34a775e0;
    ram_cell[     550] = 32'h81af1b8d;
    ram_cell[     551] = 32'hb8f6a461;
    ram_cell[     552] = 32'hc50f4101;
    ram_cell[     553] = 32'he748dbe1;
    ram_cell[     554] = 32'hdf1ed152;
    ram_cell[     555] = 32'h2df8a6e2;
    ram_cell[     556] = 32'h0ac701b7;
    ram_cell[     557] = 32'hd5388026;
    ram_cell[     558] = 32'h4870f597;
    ram_cell[     559] = 32'hbdeed43a;
    ram_cell[     560] = 32'hbd73f211;
    ram_cell[     561] = 32'hcdd18312;
    ram_cell[     562] = 32'h4cf0f2fb;
    ram_cell[     563] = 32'hcf69fac6;
    ram_cell[     564] = 32'hc2ea96bc;
    ram_cell[     565] = 32'h72c2fc7e;
    ram_cell[     566] = 32'h9fc0b37a;
    ram_cell[     567] = 32'h2a22d25b;
    ram_cell[     568] = 32'ha5a525b5;
    ram_cell[     569] = 32'h192bb680;
    ram_cell[     570] = 32'hcad639c1;
    ram_cell[     571] = 32'h20200fcb;
    ram_cell[     572] = 32'h256a5f18;
    ram_cell[     573] = 32'h3f000bde;
    ram_cell[     574] = 32'h59ef5e4e;
    ram_cell[     575] = 32'hd97302d9;
    ram_cell[     576] = 32'h2639c94f;
    ram_cell[     577] = 32'hd0b42a18;
    ram_cell[     578] = 32'h9ce585e3;
    ram_cell[     579] = 32'hd52f3d9c;
    ram_cell[     580] = 32'h6adaf88a;
    ram_cell[     581] = 32'haa68bd3b;
    ram_cell[     582] = 32'h9abd4f23;
    ram_cell[     583] = 32'h1fa605c4;
    ram_cell[     584] = 32'hd2518ac1;
    ram_cell[     585] = 32'hac6d6a74;
    ram_cell[     586] = 32'hd9719ef0;
    ram_cell[     587] = 32'h287a3a12;
    ram_cell[     588] = 32'ha8f5c571;
    ram_cell[     589] = 32'he1b6b330;
    ram_cell[     590] = 32'h8de1db4a;
    ram_cell[     591] = 32'h13da2fa7;
    ram_cell[     592] = 32'hadda34bb;
    ram_cell[     593] = 32'h1ad9f0de;
    ram_cell[     594] = 32'hfd4b341d;
    ram_cell[     595] = 32'hea0deaf5;
    ram_cell[     596] = 32'h37a54658;
    ram_cell[     597] = 32'h9cb668e0;
    ram_cell[     598] = 32'hd5703242;
    ram_cell[     599] = 32'h9a327bc0;
    ram_cell[     600] = 32'h0372e182;
    ram_cell[     601] = 32'h4d9ce7e5;
    ram_cell[     602] = 32'h32693ea7;
    ram_cell[     603] = 32'h5e7d8539;
    ram_cell[     604] = 32'h6438d82c;
    ram_cell[     605] = 32'h18754454;
    ram_cell[     606] = 32'h4d88071b;
    ram_cell[     607] = 32'hc7e7ea32;
    ram_cell[     608] = 32'hc5d4b6b3;
    ram_cell[     609] = 32'h861da966;
    ram_cell[     610] = 32'hd7681c51;
    ram_cell[     611] = 32'h37ed00f5;
    ram_cell[     612] = 32'h63b4037c;
    ram_cell[     613] = 32'h6b5563af;
    ram_cell[     614] = 32'hcdb3f114;
    ram_cell[     615] = 32'h9bfe8c65;
    ram_cell[     616] = 32'h664d3b32;
    ram_cell[     617] = 32'hf3c66bf5;
    ram_cell[     618] = 32'h41c1bf91;
    ram_cell[     619] = 32'hcc0cc2e9;
    ram_cell[     620] = 32'hf8cf9b2d;
    ram_cell[     621] = 32'h089b7594;
    ram_cell[     622] = 32'h4c818eda;
    ram_cell[     623] = 32'h322b0fd7;
    ram_cell[     624] = 32'ha133ca73;
    ram_cell[     625] = 32'h97d3dab1;
    ram_cell[     626] = 32'h524a2581;
    ram_cell[     627] = 32'hf1f33ecf;
    ram_cell[     628] = 32'hb0285480;
    ram_cell[     629] = 32'h0dcb897e;
    ram_cell[     630] = 32'hc811bdf8;
    ram_cell[     631] = 32'h2dbb8a8a;
    ram_cell[     632] = 32'h88fe88e4;
    ram_cell[     633] = 32'hff303ca8;
    ram_cell[     634] = 32'hc4c7cfc6;
    ram_cell[     635] = 32'habb9924e;
    ram_cell[     636] = 32'h62122ea3;
    ram_cell[     637] = 32'h3916dcca;
    ram_cell[     638] = 32'ha9a43fbc;
    ram_cell[     639] = 32'h1bfb9fee;
    ram_cell[     640] = 32'h837be522;
    ram_cell[     641] = 32'h14d33e2e;
    ram_cell[     642] = 32'h4622497e;
    ram_cell[     643] = 32'h29d91638;
    ram_cell[     644] = 32'h56411fdb;
    ram_cell[     645] = 32'h0267f79b;
    ram_cell[     646] = 32'hbb24f5c6;
    ram_cell[     647] = 32'h7dafb8c3;
    ram_cell[     648] = 32'h5164d033;
    ram_cell[     649] = 32'h79471a75;
    ram_cell[     650] = 32'h6f47d802;
    ram_cell[     651] = 32'hd28fe7b7;
    ram_cell[     652] = 32'h455ae0e3;
    ram_cell[     653] = 32'h5908e85a;
    ram_cell[     654] = 32'h0f091e68;
    ram_cell[     655] = 32'h3010d724;
    ram_cell[     656] = 32'hcf3f28a6;
    ram_cell[     657] = 32'hcddfa907;
    ram_cell[     658] = 32'h20b42e37;
    ram_cell[     659] = 32'h82da833b;
    ram_cell[     660] = 32'h3e01250d;
    ram_cell[     661] = 32'h22adb3a0;
    ram_cell[     662] = 32'h8f500461;
    ram_cell[     663] = 32'h1d12a8e2;
    ram_cell[     664] = 32'haa96f295;
    ram_cell[     665] = 32'h60484eb9;
    ram_cell[     666] = 32'hf394ecb1;
    ram_cell[     667] = 32'h37edb1ef;
    ram_cell[     668] = 32'hc3f8eb08;
    ram_cell[     669] = 32'h1f253d73;
    ram_cell[     670] = 32'hf459906c;
    ram_cell[     671] = 32'h15a801c9;
    ram_cell[     672] = 32'h8d1aaae5;
    ram_cell[     673] = 32'h4842f612;
    ram_cell[     674] = 32'hd45b8d95;
    ram_cell[     675] = 32'h0f83f52f;
    ram_cell[     676] = 32'h74d16961;
    ram_cell[     677] = 32'h10cd802b;
    ram_cell[     678] = 32'hbcc18bb5;
    ram_cell[     679] = 32'h97c596ac;
    ram_cell[     680] = 32'hb1546ffc;
    ram_cell[     681] = 32'h83a17808;
    ram_cell[     682] = 32'h040ee990;
    ram_cell[     683] = 32'hbfddae36;
    ram_cell[     684] = 32'he1ceb118;
    ram_cell[     685] = 32'h958af6f2;
    ram_cell[     686] = 32'hc912120b;
    ram_cell[     687] = 32'h5efee722;
    ram_cell[     688] = 32'h1dde31dd;
    ram_cell[     689] = 32'h7776ff1f;
    ram_cell[     690] = 32'hdd892573;
    ram_cell[     691] = 32'h51143d57;
    ram_cell[     692] = 32'hd6333016;
    ram_cell[     693] = 32'h9bcef1a6;
    ram_cell[     694] = 32'h2cf9a065;
    ram_cell[     695] = 32'h8d652175;
    ram_cell[     696] = 32'h9c06868d;
    ram_cell[     697] = 32'hbd85c11c;
    ram_cell[     698] = 32'hdd3bd66e;
    ram_cell[     699] = 32'h9f220323;
    ram_cell[     700] = 32'hf2576a7c;
    ram_cell[     701] = 32'hfcb69cf7;
    ram_cell[     702] = 32'h6eccc286;
    ram_cell[     703] = 32'h008c0822;
    ram_cell[     704] = 32'h68cc9934;
    ram_cell[     705] = 32'hca103edd;
    ram_cell[     706] = 32'h85d040e6;
    ram_cell[     707] = 32'hdd5544c5;
    ram_cell[     708] = 32'h4e5bac93;
    ram_cell[     709] = 32'h4a10c893;
    ram_cell[     710] = 32'h952e5b08;
    ram_cell[     711] = 32'h6f169f07;
    ram_cell[     712] = 32'ha1075847;
    ram_cell[     713] = 32'h8beffd17;
    ram_cell[     714] = 32'h187bb568;
    ram_cell[     715] = 32'h1783c699;
    ram_cell[     716] = 32'hca3e520b;
    ram_cell[     717] = 32'h063f6304;
    ram_cell[     718] = 32'h2cacfddd;
    ram_cell[     719] = 32'h7b1190ca;
    ram_cell[     720] = 32'h2f73abe0;
    ram_cell[     721] = 32'hd22e23de;
    ram_cell[     722] = 32'ha52ca1f5;
    ram_cell[     723] = 32'h3927a8f9;
    ram_cell[     724] = 32'hde31c0dd;
    ram_cell[     725] = 32'hf567c5a0;
    ram_cell[     726] = 32'hca8479ab;
    ram_cell[     727] = 32'h5feb3caa;
    ram_cell[     728] = 32'h8581d554;
    ram_cell[     729] = 32'h6cb43e1a;
    ram_cell[     730] = 32'h24eb410f;
    ram_cell[     731] = 32'h9da50bbf;
    ram_cell[     732] = 32'h9ca61cdd;
    ram_cell[     733] = 32'h0e3e8007;
    ram_cell[     734] = 32'hc3f07f6b;
    ram_cell[     735] = 32'hd47b31d8;
    ram_cell[     736] = 32'h7288e746;
    ram_cell[     737] = 32'hb36747de;
    ram_cell[     738] = 32'h295e14be;
    ram_cell[     739] = 32'h6257f197;
    ram_cell[     740] = 32'h595d4435;
    ram_cell[     741] = 32'hed3d8248;
    ram_cell[     742] = 32'h4da7c6f8;
    ram_cell[     743] = 32'h2e436a3b;
    ram_cell[     744] = 32'h794171a9;
    ram_cell[     745] = 32'h93a3c604;
    ram_cell[     746] = 32'hade87ba8;
    ram_cell[     747] = 32'h750d2e13;
    ram_cell[     748] = 32'h3163a0d7;
    ram_cell[     749] = 32'h758d4f8a;
    ram_cell[     750] = 32'he6f947c7;
    ram_cell[     751] = 32'h554ee657;
    ram_cell[     752] = 32'hc8b1f3a2;
    ram_cell[     753] = 32'h3e7305dd;
    ram_cell[     754] = 32'hdc12108e;
    ram_cell[     755] = 32'had6d1f51;
    ram_cell[     756] = 32'h28ead876;
    ram_cell[     757] = 32'h76969166;
    ram_cell[     758] = 32'h1da0a2b9;
    ram_cell[     759] = 32'h8b65a346;
    ram_cell[     760] = 32'h4d203dea;
    ram_cell[     761] = 32'hd90d7954;
    ram_cell[     762] = 32'h9ce61526;
    ram_cell[     763] = 32'h325065af;
    ram_cell[     764] = 32'h2f3e0e5a;
    ram_cell[     765] = 32'h619ccf2c;
    ram_cell[     766] = 32'h87ceec79;
    ram_cell[     767] = 32'h4be9f7ef;
end

endmodule

